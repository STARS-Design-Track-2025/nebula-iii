* NGSPICE file created from team_04.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

.subckt team_04 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XFILLER_0_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06883_ net999 net985 net979 _01808_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__and4_1
X_09671_ net337 _04423_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__nor2_1
X_08622_ net338 _03512_ _03506_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_38_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08553_ net522 net521 net406 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout162_A _05261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ net694 _02424_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__o31a_4
XANTENNA__07298__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ _03409_ _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__nor2_1
XANTENNA__07332__B _02255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07435_ datapath.rf.registers\[6\]\[19\] net814 net784 datapath.rf.registers\[5\]\[19\]
+ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a221o_1
XANTENNA__12665__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout427_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1169_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ datapath.rf.registers\[26\]\[21\] net941 net933 datapath.rf.registers\[23\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ net329 _03800_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nor2_1
XANTENNA__08262__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ datapath.rf.registers\[18\]\[22\] net791 net753 datapath.rf.registers\[22\]\[22\]
+ _02221_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ net363 _03885_ _03962_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a21o_1
XANTENNA__07470__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 datapath.rf.registers\[10\]\[14\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 datapath.rf.registers\[13\]\[14\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 datapath.rf.registers\[29\]\[14\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold373 datapath.rf.registers\[17\]\[12\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 datapath.rf.registers\[21\]\[30\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 datapath.rf.registers\[6\]\[7\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A _01806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net823 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_8
Xfanout831 net832 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_4
Xfanout842 net843 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07507__B _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _04855_ _04860_ _04863_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__or3_1
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout864 net867 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_4
Xfanout875 _01847_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_2
Xfanout886 _01841_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_4
X_09869_ _04725_ _04746_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__xnor2_1
Xfanout897 net899 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
Xhold1040 datapath.multiplication_module.multiplicand_i\[2\] vssd1 vssd1 vccd1 vccd1
+ net2406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 datapath.rf.registers\[0\]\[5\] vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 datapath.rf.registers\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net1473 _05885_ net156 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
Xhold1073 datapath.rf.registers\[31\]\[23\] vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ net245 net1854 net551 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XANTENNA__08619__A _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1084 datapath.rf.registers\[11\]\[27\] vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 datapath.rf.registers\[14\]\[29\] vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ _05499_ net176 _06230_ net179 vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14550_ net1361 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XANTENNA__07289__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ datapath.PC\[2\] _04664_ _05169_ _05238_ vssd1 vssd1 vccd1 vccd1 _06179_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13501_ clknet_leaf_78_clk _00451_ net1245 vssd1 vssd1 vccd1 vccd1 datapath.PC\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10832__A1 _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10713_ net842 _03637_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12575__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14481_ clknet_leaf_27_clk _01368_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11693_ screen.counter.currentCt\[17\] screen.counter.currentCt\[18\] _06132_ screen.counter.currentCt\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ clknet_leaf_87_clk _00388_ net1235 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ datapath.mulitply_result\[19\] net428 net662 vssd1 vssd1 vccd1 vccd1 _05501_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10575_ net1525 _03118_ net348 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ clknet_leaf_71_clk _00348_ net1229 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09450__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ net2024 net267 net476 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
X_13294_ clknet_leaf_109_clk _00284_ net1107 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12245_ net265 net2381 net484 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__mux2_1
XANTENNA__10823__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07213__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ columns.count\[1\] _06427_ net2380 vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__a21oi_1
X_11127_ _05265_ net1020 vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__nor2_4
XFILLER_0_155_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11058_ net1298 _05264_ net1297 vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__or3b_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08713__A0 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ datapath.PC\[25\] _03586_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07819__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10284__C1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12485__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ datapath.rf.registers\[0\]\[24\] net829 _02137_ _02146_ vssd1 vssd1 vccd1
+ vccd1 _02147_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07151_ net694 _02068_ _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08244__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07452__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07082_ datapath.rf.registers\[4\]\[27\] net810 net764 datapath.rf.registers\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07204__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout127 _06265_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout138 _05840_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout149 _06264_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_4
X_07984_ datapath.rf.registers\[25\]\[7\] net796 net759 datapath.rf.registers\[19\]\[7\]
+ _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a221o_1
X_09723_ _02522_ _02524_ _03873_ _04637_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_126_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06935_ _01800_ _01860_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__or2_1
XANTENNA__11303__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ net635 _04575_ _04577_ _03561_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__o2bb2a_1
X_06866_ datapath.rf.registers\[14\]\[31\] net800 net735 datapath.rf.registers\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ net656 _03529_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__nand2_1
X_06797_ datapath.MemWrite _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__nor2_1
X_09585_ net335 _04104_ net316 vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout544_A _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ net516 net515 net406 vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XANTENNA__10908__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ _03018_ net509 vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12395__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout809_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07418_ _02324_ _02344_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__or2_1
XANTENNA__07691__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08398_ _02702_ _02743_ _03322_ _02699_ _02657_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07349_ datapath.rf.registers\[6\]\[21\] net814 net810 datapath.rf.registers\[4\]\[21\]
+ _02268_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a221o_1
XANTENNA__08235__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10360_ screen.controlBus\[25\] screen.controlBus\[24\] screen.controlBus\[27\] screen.controlBus\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09019_ _03910_ _03911_ _03945_ net671 vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a22o_2
XANTENNA__10643__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ net337 _03935_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ net321 _06308_ _06309_ net325 net1890 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold170 datapath.multiplication_module.multiplicand_i\[28\] vssd1 vssd1 vccd1 vccd1
+ net1536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold181 datapath.multiplication_module.multiplicand_i\[13\] vssd1 vssd1 vccd1 vccd1
+ net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 datapath.multiplication_module.multiplicand_i\[5\] vssd1 vssd1 vccd1 vccd1
+ net1558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08340__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout650 net652 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_2
Xfanout672 _03558_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_2
Xfanout683 _03498_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_2
X_13981_ clknet_leaf_33_clk _00868_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ net289 net2319 net544 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ net163 net2554 net554 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ net205 _04816_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__nand2_1
X_12794_ net186 net2553 net563 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09120__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14533_ net1320 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11745_ screen.counter.ct\[17\] _06079_ _06098_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14464_ clknet_leaf_46_clk _01351_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11676_ screen.counter.currentCt\[13\] screen.counter.currentCt\[12\] _06122_ vssd1
+ vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__and3_1
X_14522__1348 vssd1 vssd1 vccd1 vccd1 net1348 _14522__1348/LO sky130_fd_sc_hd__conb_1
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ clknet_leaf_87_clk _00371_ net1221 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09959__C1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10627_ datapath.PC\[8\] _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14395_ clknet_leaf_19_clk _01282_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07434__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ clknet_leaf_99_clk _00331_ net1227 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10558_ _01444_ _05465_ _05466_ _05462_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[2\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11781__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ clknet_leaf_91_clk _00267_ net1204 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10489_ net121 net123 net124 net122 vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nor4b_1
XANTENNA__09187__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12228_ net194 net2248 net575 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12159_ net2368 net328 net324 _06417_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06960__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ mmio.memload_or_instruction\[24\] net1059 net1005 datapath.ru.latched_instruction\[24\]
+ net1038 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a32oi_2
XANTENNA__11297__B2 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06651_ _01452_ _01577_ _01579_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_88_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06582_ mmio.memload_or_instruction\[27\] net1062 vssd1 vssd1 vccd1 vccd1 _01512_
+ sky130_fd_sc_hd__and2_2
X_09370_ _02905_ net357 _04165_ net389 vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08321_ net646 _03244_ _03211_ _03205_ _03203_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11413__A _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ net505 net504 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07203_ datapath.rf.registers\[26\]\[24\] net822 net788 datapath.rf.registers\[23\]\[24\]
+ _02129_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ datapath.rf.registers\[16\]\[3\] net730 _03092_ _03103_ _03104_ vssd1 vssd1
+ vccd1 vccd1 _03110_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12943__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07134_ datapath.rf.registers\[11\]\[26\] net970 net901 datapath.rf.registers\[20\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07425__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11772__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07065_ _01972_ net533 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08441__B _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11524__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07967_ datapath.rf.registers\[6\]\[7\] net896 net860 datapath.rf.registers\[28\]\[7\]
+ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a221o_1
XANTENNA__06951__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09706_ _02172_ _04500_ _04631_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__and4_1
XFILLER_0_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06918_ datapath.rf.registers\[17\]\[31\] net881 net878 datapath.rf.registers\[29\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XANTENNA__11288__B2 mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ datapath.rf.registers\[31\]\[9\] net818 net723 datapath.rf.registers\[27\]\[9\]
+ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ _03347_ _04563_ net642 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a21o_1
X_06849_ _01639_ net998 net982 net977 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__and4_2
XANTENNA_fanout926_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _04478_ _04490_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08519_ net656 _03444_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__nand2_4
XANTENNA__10799__A0 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09499_ net380 _04154_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ screen.register.currentXbus\[13\] _05709_ _05772_ screen.register.currentYbus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__a22o_1
XANTENNA__07664__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08335__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12853__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08208__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11461_ screen.register.currentXbus\[25\] _05700_ _05772_ screen.register.currentYbus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09405__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13200_ clknet_leaf_4_clk _00192_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10412_ datapath.multiplication_module.mul_prev _01636_ vssd1 vssd1 vccd1 vccd1 _05332_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11392_ screen.register.currentYbus\[15\] net132 _05881_ net161 vssd1 vssd1 vccd1
+ vccd1 _00373_ sky130_fd_sc_hd__a22o_1
X_14180_ clknet_leaf_17_clk _01067_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13131_ clknet_leaf_18_clk _00123_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10343_ net1297 net1298 _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__or3_2
XFILLER_0_131_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13062_ clknet_leaf_106_clk _00054_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10274_ net337 _03898_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12013_ datapath.mulitply_result\[6\] datapath.multiplication_module.multiplicand_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__nand2_1
XANTENNA__10723__B1 _05567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09463__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout480 _06449_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06942__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout491 _03556_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11279__B2 mmio.memload_or_instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13964_ clknet_leaf_30_clk _00851_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09341__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ net1576 net235 net545 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
X_13895_ clknet_leaf_25_clk _00782_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ net249 net2074 net553 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ net263 net2311 net561 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11233__A datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14516_ clknet_leaf_115_clk _01403_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_140_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11728_ screen.counter.ct\[10\] _06076_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14447_ clknet_leaf_6_clk _01334_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12763__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11659_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07407__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11203__B2 _05048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14378_ clknet_leaf_9_clk _01265_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold906 datapath.rf.registers\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 datapath.multiplication_module.multiplicand_i\[17\] vssd1 vssd1 vccd1 vccd1
+ net2283 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ clknet_leaf_77_clk net1367 net1246 vssd1 vssd1 vccd1 vccd1 mmio.WEN2 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08080__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold928 datapath.rf.registers\[24\]\[21\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10962__A0 _05590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold939 datapath.rf.registers\[22\]\[31\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08870_ net420 _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07186__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ datapath.rf.registers\[2\]\[10\] net920 net848 datapath.rf.registers\[1\]\[10\]
+ _02745_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a221o_1
XANTENNA__06933__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__inv_2
XANTENNA__08135__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__A0 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06703_ datapath.ru.latched_instruction\[13\] net1041 _01630_ vssd1 vssd1 vccd1 vccd1
+ _01631_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12938__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ _02588_ net519 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__nand2_1
XANTENNA__06697__A1 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ net396 _04213_ _04348_ net400 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__a211o_1
X_06634_ mmio.memload_or_instruction\[14\] mmio.memload_or_instruction\[13\] mmio.memload_or_instruction\[12\]
+ mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__and4b_1
XANTENNA__07894__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ net507 _03061_ net684 vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__o21a_1
X_06565_ mmio.memload_or_instruction\[18\] net1058 vssd1 vssd1 vccd1 vccd1 _01495_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08438__A2 _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09096__C1 _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08304_ datapath.rf.registers\[17\]\[1\] _01735_ _01758_ vssd1 vssd1 vccd1 vccd1
+ _03231_ sky130_fd_sc_hd__and3_1
XANTENNA__07646__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06496_ datapath.PC\[13\] vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
X_09284_ _02905_ _02855_ net354 vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08235_ datapath.rf.registers\[18\]\[2\] net792 net733 datapath.rf.registers\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a22o_1
XANTENNA__12673__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1151_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout507_A _03039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09548__A _03785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ datapath.rf.registers\[7\]\[3\] net993 _01739_ vssd1 vssd1 vccd1 vccd1 _03093_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_151_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07117_ datapath.rf.registers\[18\]\[26\] net790 net731 datapath.rf.registers\[16\]\[26\]
+ _02041_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a221o_1
X_08097_ datapath.rf.registers\[26\]\[4\] net941 net889 datapath.rf.registers\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07048_ datapath.rf.registers\[19\]\[28\] net945 net917 datapath.rf.registers\[10\]\[28\]
+ _01974_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout876_A _01844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10921__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10181__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__A mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ net376 _03925_ _03917_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__o21a_1
XANTENNA__09433__D _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10961_ net297 net2386 net586 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__mux2_1
XANTENNA__12848__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net181 net2355 net569 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__mux2_1
X_13680_ clknet_leaf_110_clk _00615_ net1103 vssd1 vssd1 vccd1 vccd1 columns.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10892_ net289 net1578 net595 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ net1825 net170 net441 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08346__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12562_ net191 net2450 net450 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07101__A2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14301_ clknet_leaf_32_clk _01188_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11513_ screen.register.currentYbus\[20\] _05735_ _05737_ screen.register.currentYbus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a22o_1
XANTENNA__12583__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ net209 net1763 net458 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire155 _05263_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_1
X_14232_ clknet_leaf_40_clk _01119_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11444_ _05304_ _05784_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08062__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ clknet_leaf_59_clk _01050_ net1267 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11375_ _02926_ net669 vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13114_ clknet_leaf_23_clk _00106_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ mmio.wishbone.curr_state\[2\] mmio.wishbone.curr_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _05252_ sky130_fd_sc_hd__nor2_2
X_14094_ clknet_leaf_116_clk _00981_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13045_ clknet_leaf_28_clk _00037_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10257_ net835 _04935_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07168__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__A _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1231 net1254 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_4
Xfanout1242 net1254 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_2
X_10188_ _05114_ net834 _04418_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__or3b_1
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10172__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1264 net1266 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06915__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1275 datapath.PC\[18\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_2
XFILLER_0_89_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1286 screen.counter.ct\[16\] vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__buf_1
Xfanout1297 screen.counter.ct\[3\] vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__clkbuf_2
X_13947_ clknet_leaf_19_clk _00834_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12758__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06679__A1 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07876__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_26_clk _00765_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07340__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ net167 net2116 net558 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
XANTENNA__07628__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12493__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08020_ datapath.rf.registers\[15\]\[6\] net856 net852 datapath.rf.registers\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold703 datapath.rf.registers\[8\]\[13\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 datapath.rf.registers\[16\]\[30\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 datapath.rf.registers\[28\]\[21\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold736 datapath.rf.registers\[16\]\[28\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 datapath.rf.registers\[19\]\[25\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold758 datapath.rf.registers\[14\]\[30\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold769 datapath.rf.registers\[16\]\[24\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _04895_ _04897_ datapath.PC\[28\] net1272 vssd1 vssd1 vccd1 vccd1 _04898_
+ sky130_fd_sc_hd__o2bb2a_1
X_08922_ _03715_ _03716_ net375 vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a21o_1
XANTENNA__10741__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__C1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _03421_ _03748_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout192_A _05544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07804_ datapath.rf.registers\[29\]\[11\] net876 net856 datapath.rf.registers\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
X_08784_ _02079_ net359 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ _02660_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__or2_1
XANTENNA__12668__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout457_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ datapath.rf.registers\[16\]\[14\] net960 net936 datapath.rf.registers\[21\]\[14\]
+ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09405_ net639 _04321_ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__a21o_1
X_06617_ datapath.ru.latched_instruction\[9\] _01515_ _01544_ _01545_ _01546_ vssd1
+ vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09069__C1 _03995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07597_ _02501_ net521 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__and2_1
XANTENNA__07619__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ _04261_ _04262_ net399 vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__a21o_1
X_06548_ mmio.key_data\[2\] mmio.memload_or_instruction\[2\] net1060 vssd1 vssd1 vccd1
+ vccd1 _01478_ sky130_fd_sc_hd__mux2_2
XFILLER_0_145_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09267_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__inv_2
XANTENNA__10916__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06479_ datapath.ru.latched_instruction\[7\] vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
X_08218_ net696 _03135_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__or3_1
X_09198_ net510 _02973_ _03497_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08149_ datapath.rf.registers\[26\]\[3\] net940 net869 datapath.rf.registers\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07398__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _05748_ _05752_ _05805_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__or3_2
X_10111_ _01424_ net1243 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__nor2_1
X_11091_ _05739_ _05740_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nor2_1
X_10042_ net537 _04471_ _04968_ net1056 vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a211o_1
Xhold30 keypad.decode.d2 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 keypad.apps.button\[1\] vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 net61 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 screen.controlBus\[15\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold74 net116 vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 net70 vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_3_clk _00688_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold96 net53 vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12578__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11993_ _06277_ _06278_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__xnor2_1
X_13732_ clknet_leaf_101_clk _00619_ net1223 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_67_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10944_ net242 net1807 net592 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
XANTENNA__07322__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13663_ clknet_leaf_57_clk _00601_ net1257 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10875_ net244 net1970 net600 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12614_ net1872 net253 net440 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ clknet_leaf_81_clk net1386 net1238 vssd1 vssd1 vccd1 vccd1 screen.register.xFill2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12545_ net267 net2506 net448 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10826__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12476_ net278 net1814 net456 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XANTENNA__08092__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ clknet_leaf_15_clk _01102_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11427_ net1017 _05745_ _05746_ _05798_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__a311o_1
XANTENNA__08035__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07389__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output86_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ clknet_leaf_42_clk _01033_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11358_ keypad.apps.button\[4\] _05829_ _05861_ keypad.apps.button\[3\] vssd1 vssd1
+ vccd1 vccd1 _05864_ sky130_fd_sc_hd__or4b_1
XFILLER_0_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ datapath.PC\[0\] _05235_ net1245 vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14077_ clknet_leaf_24_clk _00964_ net1143 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ net9 net1044 net1033 net2593 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__o22a_1
X_13028_ clknet_leaf_102_clk _00020_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1050 _05397_ vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_2
Xfanout1061 net1062 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
Xfanout1072 net1076 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07155__B _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1083 net1084 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
Xfanout1094 net1096 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07561__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire425_A _01971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12488__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ datapath.rf.registers\[17\]\[17\] net765 net729 datapath.rf.registers\[2\]\[17\]
+ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a221o_1
XANTENNA__07849__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07313__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07451_ datapath.rf.registers\[22\]\[19\] net953 net858 datapath.rf.registers\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07382_ datapath.rf.registers\[7\]\[20\] net826 net801 datapath.rf.registers\[14\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09121_ _02743_ _02744_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11421__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_98_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08003_ net512 _02927_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08026__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12951__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 datapath.rf.registers\[11\]\[2\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 datapath.rf.registers\[22\]\[19\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 datapath.mulitply_result\[20\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold533 datapath.rf.registers\[31\]\[3\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 datapath.rf.registers\[27\]\[4\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 datapath.rf.registers\[16\]\[19\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 datapath.rf.registers\[16\]\[9\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold577 datapath.rf.registers\[5\]\[29\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 datapath.rf.registers\[29\]\[15\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net1057 _03591_ _04880_ net845 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__a31o_1
Xhold599 datapath.rf.registers\[15\]\[21\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _02390_ _02391_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__and2b_1
X_09885_ _04809_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__and2b_1
Xhold1200 datapath.rf.registers\[11\]\[6\] vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13927__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 datapath.rf.registers\[19\]\[31\] vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 datapath.rf.registers\[31\]\[29\] vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07065__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08836_ _03630_ _03762_ net401 vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__mux2_1
Xhold1233 datapath.rf.registers\[17\]\[26\] vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 datapath.rf.registers\[19\]\[27\] vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 screen.counter.currentCt\[1\] vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 datapath.rf.registers\[23\]\[28\] vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12398__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1277 datapath.rf.registers\[6\]\[1\] vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net338 _03693_ net315 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout741_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ datapath.rf.registers\[11\]\[13\] net968 net896 datapath.rf.registers\[6\]\[13\]
+ _02642_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _01682_ net622 vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07649_ datapath.rf.registers\[7\]\[14\] net824 net796 datapath.rf.registers\[25\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ datapath.PC\[21\] datapath.PC\[22\] _05503_ vssd1 vssd1 vccd1 vccd1 _05514_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09319_ net365 _03670_ _03671_ net373 vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_11_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08265__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_114_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10591_ net2406 net506 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[3\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12330_ net2418 net194 net478 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08343__C _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net195 net2401 net485 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__mux2_1
XANTENNA__12861__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__C1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ clknet_leaf_3_clk _00887_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11212_ net1599 net143 net137 _05103_ vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__a22o_1
XANTENNA__09736__A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ _06438_ _06439_ _06436_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__o21a_1
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
X_11143_ _05726_ net1014 _05747_ _05791_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__or4_1
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07791__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
X_11074_ net1022 _05715_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__nor2_1
XANTENNA__10127__A1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _04474_ _04949_ _04951_ _04921_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__o211a_1
XANTENNA__11875__A1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output124_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ net172 net2588 net581 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__mux2_1
X_13715_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[0\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ net287 net1611 net591 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13646_ clknet_leaf_68_clk _00584_ net1225 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ net288 net1556 net599 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08256__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_105_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13577_ clknet_leaf_88_clk _00527_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10789_ net1277 _05485_ datapath.PC\[10\] vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12528_ net1790 net192 net454 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08008__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12771__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ net213 net2236 net462 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
XANTENNA__08559__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14129_ clknet_leaf_8_clk _01016_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout309 _05860_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
XANTENNA__09508__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ datapath.rf.registers\[21\]\[30\] net746 net727 datapath.rf.registers\[2\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a22o_1
XANTENNA__06990__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _03449_ _04433_ _04591_ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o211a_1
X_06882_ net1001 net983 net979 _01808_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__and4_1
XANTENNA__07534__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ net333 net377 _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_38_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08552_ net523 _02431_ net406 vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07503_ datapath.rf.registers\[0\]\[18\] net692 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__or2_1
XANTENNA__12291__A1 _05519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _03405_ _03406_ _02701_ _03379_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o211a_1
XANTENNA__12946__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07434_ datapath.rf.registers\[15\]\[19\] net805 net735 datapath.rf.registers\[12\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07365_ datapath.rf.registers\[22\]\[21\] net953 net905 datapath.rf.registers\[24\]\[21\]
+ _02291_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout322_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08444__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _03808_ _04030_ net380 vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14126__RESET_B net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07296_ datapath.rf.registers\[20\]\[22\] net803 net732 datapath.rf.registers\[16\]\[22\]
+ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a221o_1
XANTENNA__08163__C _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09035_ net367 _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12681__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1231_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold330 datapath.rf.registers\[13\]\[3\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 datapath.rf.registers\[29\]\[4\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 datapath.rf.registers\[5\]\[6\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 datapath.rf.registers\[23\]\[12\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 datapath.rf.registers\[2\]\[25\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 datapath.rf.registers\[1\]\[25\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 datapath.rf.registers\[15\]\[30\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net812 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__buf_4
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_4
Xfanout832 _01736_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_8
X_09937_ _04855_ _04860_ _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__o21ai_1
Xfanout843 _01720_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout956_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_4
Xfanout865 net867 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_4
Xfanout876 _01844_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_4
X_09868_ _04792_ _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__nor2_1
Xfanout887 _01841_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
Xhold1030 datapath.rf.registers\[14\]\[17\] vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_4
XANTENNA__07525__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1041 datapath.rf.registers\[25\]\[20\] vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _03706_ _03741_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a21o_1
Xhold1052 datapath.rf.registers\[4\]\[26\] vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 datapath.rf.registers\[10\]\[15\] vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ datapath.PC\[5\] _02998_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__or2_1
Xhold1074 datapath.rf.registers\[7\]\[22\] vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 datapath.rf.registers\[26\]\[31\] vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net834 _04825_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__nand2_1
Xhold1096 datapath.rf.registers\[16\]\[4\] vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10230__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__C _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ _05384_ _06177_ _01578_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__a21o_1
XANTENNA__12856__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ clknet_leaf_79_clk _00450_ net1243 vssd1 vssd1 vccd1 vccd1 datapath.PC\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ net842 _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14480_ clknet_leaf_0_clk _01367_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10832__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11692_ net1517 _06134_ _06136_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13431_ clknet_leaf_79_clk _00387_ net1244 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08238__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10643_ _03872_ _05499_ net845 vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ clknet_leaf_95_clk _00347_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ datapath.multiplication_module.multiplier_i\[3\] _03176_ net348 vssd1 vssd1
+ vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[2\] sky130_fd_sc_hd__mux2_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__A2 _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12313_ net2434 net270 net478 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XANTENNA__12591__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ clknet_4_13_0_clk _00283_ net1266 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
X_12244_ net269 net2570 net485 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ columns.count\[1\] columns.count\[2\] _06427_ vssd1 vssd1 vccd1 vccd1 _06429_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11000__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _05699_ net1020 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__nor2_4
XANTENNA__06972__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ net1022 _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__nor2_4
XANTENNA__11848__A1 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07516__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ net536 net1051 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nand2_1
XANTENNA__09269__A2 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12766__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11959_ net259 net2158 net578 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13629_ clknet_leaf_54_clk _00567_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_17_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09426__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ _02070_ _02072_ _02074_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_95_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07081_ datapath.rf.registers\[1\]\[27\] net742 _02007_ _01736_ vssd1 vssd1 vccd1
+ vccd1 _02008_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09376__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__A _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07755__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_26_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07983_ datapath.rf.registers\[9\]\[7\] net778 net734 datapath.rf.registers\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a22o_1
Xfanout139 _05840_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
XANTENNA__06963__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _04644_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nor2_1
X_06934_ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__inv_2
XANTENNA__11839__B2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09653_ _03347_ _04563_ _03556_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06865_ _01781_ _01787_ _01789_ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout272_A _05622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08439__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ net654 net637 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ net639 _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__and2_1
X_06796_ _01602_ net835 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ _03460_ _03461_ net409 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
XANTENNA__12676__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_35_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ _03066_ _03391_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and2b_1
XANTENNA__07140__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07417_ net524 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08397_ _02702_ _02743_ _03322_ _02699_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout704_A _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07348_ _02272_ _02273_ _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10578__A1 _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07279_ _02201_ _02203_ _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07994__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ _03938_ _03940_ _03944_ _03915_ net429 vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a311o_1
X_10290_ net394 _05215_ _05216_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold160 datapath.rf.registers\[14\]\[0\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 datapath.rf.registers\[17\]\[3\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold182 datapath.rf.registers\[4\]\[7\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold193 net76 vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06954__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _03505_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 datapath.MemRead vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_4
X_13980_ clknet_leaf_55_clk _00867_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
Xfanout684 _03497_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout695 net697 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_4
X_12931_ net182 net1635 net544 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__mux2_1
X_12862_ net168 net2257 net555 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ datapath.PC\[14\] net303 _06217_ _05161_ vssd1 vssd1 vccd1 vccd1 _00458_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12586__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ net188 net2638 net563 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14532_ net1319 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
X_11744_ net1284 net664 vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__nand2_1
XANTENNA__10805__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14463_ clknet_leaf_37_clk _01350_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11675_ screen.counter.currentCt\[11\] screen.counter.currentCt\[12\] _06120_ screen.counter.currentCt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a31o_1
X_13414_ clknet_leaf_87_clk _00370_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ datapath.PC\[6\] datapath.PC\[7\] _05483_ vssd1 vssd1 vccd1 vccd1 _05484_
+ sky130_fd_sc_hd__and3_1
X_14394_ clknet_leaf_23_clk _01281_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ clknet_leaf_99_clk _00330_ net1227 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_77_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ net1050 _05426_ _05456_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__or3b_1
XANTENNA__11230__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07985__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ clknet_leaf_92_clk _00266_ net1204 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10488_ net121 net122 net124 net123 vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__or4b_2
XANTENNA__09187__A1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ net199 net1751 net576 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07737__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12158_ _06413_ _06416_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_9_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06945__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net1290 net1291 _05749_ _05758_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__or4_1
X_12089_ _06352_ _06354_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__nor2_1
XANTENNA__08147__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06650_ _01579_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__inv_2
XANTENNA__07370__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06581_ mmio.memload_or_instruction\[16\] net1058 vssd1 vssd1 vccd1 vccd1 _01511_
+ sky130_fd_sc_hd__and2_2
XANTENNA__12496__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14471__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ net649 _03244_ _03211_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08275__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11413__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ net650 _03148_ _03175_ _03177_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a31o_2
XFILLER_0_117_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07202_ datapath.rf.registers\[14\]\[24\] net801 net736 datapath.rf.registers\[12\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ _03097_ _03106_ _03107_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07133_ net652 _02059_ _01729_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_119_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07976__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ datapath.rf.registers\[0\]\[28\] net692 _01978_ _01990_ vssd1 vssd1 vccd1
+ vccd1 _01991_ sky130_fd_sc_hd__o22a_4
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1027_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07966_ datapath.rf.registers\[10\]\[7\] net916 net908 datapath.rf.registers\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a22o_1
X_09705_ _01864_ _01910_ _01996_ _03596_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__and4_1
X_06917_ net999 net983 net980 _01812_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__and4_4
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07897_ datapath.rf.registers\[13\]\[9\] net793 net720 datapath.rf.registers\[28\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a22o_1
XANTENNA__08169__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout654_A _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__A2 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09350__B2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _02040_ _03346_ _01996_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__o21ai_1
X_06848_ net996 _01731_ _01742_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ _04489_ _04491_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__a21o_1
XANTENNA__10919__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06779_ _01465_ _01469_ _01497_ _01504_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout821_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08518_ _01625_ _03443_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09498_ net376 _04147_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ _02547_ net520 vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ screen.register.currentXbus\[1\] _05704_ _05776_ screen.register.currentYbus\[9\]
+ _05773_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a221o_1
X_10411_ _05037_ _05331_ vssd1 vssd1 vccd1 vccd1 mmio.ack_center.key_en sky130_fd_sc_hd__nor2_1
XANTENNA__08613__A0 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ net423 net714 vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07967__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ clknet_leaf_12_clk _00122_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10342_ net1300 net1301 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13061_ clknet_leaf_95_clk _00053_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ net400 _05198_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_72_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12012_ net322 _06293_ _06294_ net326 net2581 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a32o_1
XANTENNA__10723__A1 _01492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11920__B1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_8
Xfanout481 _06449_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11279__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout492 _03555_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
X_13963_ clknet_leaf_56_clk _00850_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08144__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09341__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12914_ net1737 net240 net547 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
X_13894_ clknet_leaf_111_clk _00781_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12845_ net253 net2284 net553 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ net268 net1876 net561 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__mux2_1
XANTENNA__07104__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ net1292 net663 _06157_ net712 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a22o_1
X_14515_ clknet_leaf_59_clk _01402_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11658_ screen.counter.currentCt\[7\] screen.counter.currentCt\[6\] _06110_ vssd1
+ vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and3_1
X_14446_ clknet_leaf_118_clk _01333_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ net1452 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_142_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14377_ clknet_leaf_2_clk _01264_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11203__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11589_ _05705_ _05760_ _05805_ _05763_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold907 datapath.rf.registers\[22\]\[25\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold918 datapath.rf.registers\[20\]\[13\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ clknet_leaf_75_clk _00318_ net1250 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold929 datapath.rf.registers\[24\]\[15\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13259_ clknet_leaf_63_clk _00249_ net1271 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06918__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ datapath.rf.registers\[10\]\[10\] net916 net868 datapath.rf.registers\[27\]\[10\]
+ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09580__A1 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ net652 _02677_ net627 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
X_06702_ _01628_ _01629_ net1008 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__o21a_1
XANTENNA__08135__A2 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__A1 _03087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ net519 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__inv_2
XANTENNA__07343__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ _04058_ _04059_ net396 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a21oi_1
X_06633_ mmio.memload_or_instruction\[24\] mmio.memload_or_instruction\[26\] mmio.memload_or_instruction\[25\]
+ mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ _03068_ _03390_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__xnor2_1
X_06564_ net1306 net1302 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ _01494_ sky130_fd_sc_hd__or3b_2
XFILLER_0_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08303_ datapath.rf.registers\[1\]\[1\] net974 _01735_ vssd1 vssd1 vccd1 vccd1 _03230_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ net636 _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__and2_1
X_06495_ datapath.PC\[10\] vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
XANTENNA__12954__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout235_A _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ datapath.rf.registers\[10\]\[2\] _01772_ _03149_ _03150_ _03158_ vssd1 vssd1
+ vccd1 vccd1 _03161_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08165_ datapath.rf.registers\[9\]\[3\] net993 _01754_ vssd1 vssd1 vccd1 vccd1 _03092_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_151_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1144_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07116_ datapath.rf.registers\[6\]\[26\] net814 net727 datapath.rf.registers\[2\]\[26\]
+ _02042_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a221o_1
X_08096_ datapath.rf.registers\[21\]\[4\] net936 net909 datapath.rf.registers\[30\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a22o_1
XANTENNA__08171__C _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ datapath.rf.registers\[16\]\[28\] net962 net938 datapath.rf.registers\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XANTENNA__07068__B _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout771_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A _01848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__B _04209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net374 _03924_ _03918_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_149_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07582__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__B net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__inv_2
XANTENNA__10222__B _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08126__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10469__B1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ net289 net1969 net586 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ net689 _04543_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a21o_1
X_10891_ net183 net1501 net595 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__mux2_1
XANTENNA__08627__B _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ net1809 net171 net442 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08346__C _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ net195 net2557 net449 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11512_ screen.register.currentXbus\[4\] _05720_ _05736_ screen.register.currentYbus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__a22o_1
X_14300_ clknet_leaf_53_clk _01187_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12492_ net213 net2482 net458 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__mux2_1
X_14231_ clknet_leaf_46_clk _01118_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11443_ screen.register.currentYbus\[0\] _05772_ _05912_ _05914_ _05915_ vssd1 vssd1
+ vccd1 vccd1 _05916_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_124_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09458__B _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ clknet_leaf_36_clk _01049_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11374_ net2586 net132 _05872_ net161 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13113_ clknet_leaf_47_clk _00105_ net1197 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10325_ _05248_ _05251_ vssd1 vssd1 vccd1 vccd1 mmio.WEN sky130_fd_sc_hd__nand2_1
XFILLER_0_132_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14093_ clknet_leaf_0_clk _00980_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06612__A2 _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ clknet_leaf_116_clk _00036_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10256_ net844 _04661_ _05182_ net835 vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__o211a_1
Xfanout1210 net1212 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_2
Xfanout1221 net1222 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08365__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1235 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_4
X_10187_ _04081_ _04417_ _04047_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__o21a_1
Xfanout1243 net1244 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__B1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__buf_2
Xfanout1265 net1266 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__clkbuf_2
Xfanout1276 datapath.PC\[12\] vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_2
Xfanout1287 screen.counter.ct\[15\] vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
Xfanout1298 net1299 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08117__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_13946_ clknet_leaf_23_clk _00833_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07325__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13877_ clknet_leaf_29_clk _00764_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12828_ net172 net1881 net559 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11424__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12774__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ net192 net2599 net567 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14429_ clknet_leaf_24_clk _01316_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold704 datapath.rf.registers\[12\]\[0\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold715 datapath.rf.registers\[25\]\[22\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 datapath.rf.registers\[27\]\[13\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 datapath.rf.registers\[18\]\[29\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 datapath.rf.registers\[10\]\[10\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ net207 _04896_ net1313 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a21oi_1
Xhold759 datapath.rf.registers\[9\]\[27\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
X_08921_ net367 _03847_ _03846_ net371 vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a211o_1
XANTENNA__10148__C1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06801__A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11419__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10699__B1 _05546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _03336_ _03748_ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__o21a_1
X_07803_ datapath.rf.registers\[6\]\[11\] net896 net892 datapath.rf.registers\[14\]\[11\]
+ _02729_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a221o_1
X_08783_ net362 _03621_ _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a21o_1
XANTENNA__12949__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout185_A _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08108__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07734_ datapath.rf.registers\[18\]\[12\] net789 net730 datapath.rf.registers\[16\]\[12\]
+ _02659_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a221o_1
XANTENNA__09305__B2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ datapath.rf.registers\[8\]\[14\] net924 net864 datapath.rf.registers\[13\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ net335 _03763_ _04326_ net640 vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__o211a_1
X_06616_ datapath.ru.latched_instruction\[22\] _01486_ _01510_ datapath.ru.latched_instruction\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_9_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09069__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07596_ _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__inv_2
XANTENNA__08166__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07619__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ net387 _04259_ net394 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__o21a_1
X_06547_ mmio.key_data\[4\] net1060 _01475_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__o21a_2
XANTENNA__12684__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _03127_ _03388_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07095__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ datapath.ru.latched_instruction\[6\] vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08217_ _03137_ _03139_ _03141_ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__or4_1
X_09197_ net415 _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nand2_1
XANTENNA__12376__A0 _05607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ datapath.rf.registers\[30\]\[3\] net909 net884 datapath.rf.registers\[9\]\[3\]
+ _03074_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__a221o_1
XANTENNA__08044__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout986_A _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10932__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08079_ datapath.rf.registers\[18\]\[5\] net789 net770 datapath.rf.registers\[30\]\[5\]
+ _03005_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__a221o_1
X_10110_ _05035_ _05036_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__or2_2
XFILLER_0_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11090_ _05728_ net1021 vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__nor2_1
XANTENNA__08347__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ net1275 net540 vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__nor2_1
Xhold20 screen.register.xFill1 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__A1 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 datapath.i_ack vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08752__C1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 net48 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 net58 vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 datapath.multiplication_module.multiplier_i\[1\] vssd1 vssd1 vccd1 vccd1 net1430
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12859__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 net83 vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11763__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13800_ clknet_leaf_14_clk _00687_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold86 datapath.multiplication_module.multiplicand_i\[20\] vssd1 vssd1 vccd1 vccd1
+ net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net89 vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ datapath.mulitply_result\[1\] datapath.multiplication_module.multiplicand_i\[1\]
+ _06272_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10943_ net235 net2312 net590 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
X_13731_ clknet_leaf_104_clk _00618_ net1121 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10311__C1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10874_ net236 net2352 net598 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__mux2_1
X_13662_ clknet_leaf_57_clk _00600_ net1259 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12613_ net1782 net257 net440 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__mux2_1
X_13593_ clknet_leaf_80_clk screen.register.xFill net1233 vssd1 vssd1 vccd1 vccd1
+ screen.register.xFill1 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12594__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12544_ net271 net2154 net449 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12475_ net280 net2268 net456 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XANTENNA__11003__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14214_ clknet_leaf_114_clk _01101_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11426_ _05799_ _05817_ _05762_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a21oi_1
XANTENNA_6 _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ clknet_leaf_42_clk _01032_ net1162 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11357_ net2628 net2251 _05862_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XANTENNA__10842__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10308_ datapath.PC\[0\] _05234_ _05184_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__mux2_1
X_14076_ clknet_leaf_55_clk _00963_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ net8 net1044 net1033 mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1
+ vccd1 _00302_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_111_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ clknet_leaf_104_clk _00019_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10239_ _05092_ _05103_ _05113_ _05154_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__or4_1
XANTENNA__07546__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10145__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__A1 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__buf_4
Xfanout1051 net1054 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
Xfanout1062 _01455_ vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07010__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1073 net1075 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12769__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929_ clknet_leaf_2_clk _00816_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13604__D net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07450_ datapath.rf.registers\[23\]\[19\] net933 net901 datapath.rf.registers\[20\]\[19\]
+ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07381_ datapath.rf.registers\[6\]\[20\] net815 net794 datapath.rf.registers\[13\]\[20\]
+ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09120_ _04041_ _04045_ net675 _04008_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_33_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07077__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09051_ _02656_ _02657_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_142_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11421__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ net512 _02927_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__and2b_1
Xhold501 datapath.rf.registers\[17\]\[1\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 datapath.rf.registers\[21\]\[0\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 datapath.rf.registers\[22\]\[27\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 datapath.rf.registers\[19\]\[6\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 datapath.rf.registers\[10\]\[22\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 datapath.rf.registers\[4\]\[14\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07785__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 datapath.rf.registers\[13\]\[9\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold578 datapath.rf.registers\[29\]\[22\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06531__A mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold589 datapath.rf.registers\[31\]\[4\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ datapath.PC\[29\] _03590_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
X_08904_ net673 _03786_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__o21ai_2
XANTENNA__11333__A1 _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _04757_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07537__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__B2 datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1201 datapath.rf.registers\[16\]\[15\] vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 datapath.rf.registers\[28\]\[20\] vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 datapath.rf.registers\[31\]\[14\] vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ _03757_ _03761_ net394 vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__mux2_1
Xhold1234 datapath.rf.registers\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12679__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 datapath.rf.registers\[23\]\[29\] vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout567_A _06465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 datapath.rf.registers\[24\]\[10\] vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1215_A datapath.mulitply_result\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ net398 _03692_ _03516_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__o21a_1
Xhold1267 datapath.rf.registers\[19\]\[16\] vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 screen.counter.ct\[11\] vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
X_07717_ datapath.rf.registers\[4\]\[13\] net928 net884 datapath.rf.registers\[9\]\[13\]
+ _02643_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a221o_1
XANTENNA__10199__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ net333 net377 _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout734_A _01777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08177__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ datapath.rf.registers\[14\]\[14\] net799 net734 datapath.rf.registers\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10927__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ datapath.rf.registers\[31\]\[16\] net950 net894 datapath.rf.registers\[14\]\[16\]
+ _02505_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09318_ net376 _04243_ _04244_ net331 vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_62_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10590_ net2325 net505 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[2\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09462__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06706__A _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _03687_ _03689_ net388 vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12260_ net196 net1740 net486 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11211_ net1518 net144 net138 _05123_ vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__a22o_1
X_12191_ columns.count\[7\] _06434_ columns.count\[8\] vssd1 vssd1 vccd1 vccd1 _06439_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__09736__B _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _05747_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nor2_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__07240__A2 _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__09517__A1 _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11257__A1_N _02234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
X_11073_ net1023 _05705_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or2_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__11324__B2 _01456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ net1052 _04950_ _04948_ net704 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__a211o_1
XANTENNA__12589__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11875__A2 _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11975_ net187 net2498 net580 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
X_13714_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[31\]
+ net1262 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ net181 net2172 net591 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__mux2_1
XANTENNA__07700__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ net180 net2441 net599 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__mux2_1
X_13645_ clknet_leaf_69_clk _00583_ net1225 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07059__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13576_ clknet_leaf_88_clk _00526_ net1219 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09453__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10788_ net2225 net271 net604 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11260__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12527_ net1664 net196 net453 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12458_ net218 net2235 net462 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11409_ net530 net714 vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__nor2_1
X_12389_ net226 net1697 net469 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07767__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14128_ clknet_leaf_4_clk _01015_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ datapath.rf.registers\[10\]\[30\] net749 _01876_ net832 vssd1 vssd1 vccd1
+ vccd1 _01877_ sky130_fd_sc_hd__a211o_1
X_14059_ clknet_leaf_18_clk _00946_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07519__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ _01673_ _01675_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a211oi_4
XANTENNA__12499__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ net371 net362 _03546_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__or3_1
XANTENNA__08278__A datapath.rf.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ _03476_ _03477_ net409 vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07502_ datapath.rf.registers\[14\]\[18\] net893 _02412_ _02425_ _02428_ vssd1 vssd1
+ vccd1 vccd1 _02429_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_141_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08482_ _03378_ _03380_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__nor2_1
XANTENNA__07298__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07433_ datapath.rf.registers\[9\]\[19\] net779 net770 datapath.rf.registers\[30\]\[19\]
+ _02359_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ datapath.rf.registers\[4\]\[21\] net930 net870 datapath.rf.registers\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ net369 _03924_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a21o_1
XANTENNA__10054__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11251__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12962__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ datapath.rf.registers\[25\]\[22\] net798 net721 datapath.rf.registers\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1057_A _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ net497 net494 net520 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07470__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 datapath.rf.registers\[12\]\[26\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 datapath.rf.registers\[6\]\[19\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1224_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 datapath.rf.registers\[3\]\[29\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold353 datapath.rf.registers\[29\]\[28\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 datapath.rf.registers\[22\]\[29\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold375 datapath.rf.registers\[10\]\[5\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10762__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 datapath.rf.registers\[22\]\[5\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 _01753_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_4
Xhold397 datapath.rf.registers\[9\]\[24\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_4
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
X_09936_ _04861_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__xnor2_1
Xfanout833 net838 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_4
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_4
Xfanout855 _01855_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_4
Xfanout877 _01844_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_2
X_09867_ _04744_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__xnor2_1
Xfanout888 net891 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_4
Xhold1020 datapath.rf.registers\[29\]\[2\] vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 _01836_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout949_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1031 datapath.rf.registers\[26\]\[21\] vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 datapath.rf.registers\[7\]\[2\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12202__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1053 datapath.rf.registers\[4\]\[4\] vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _03739_ _03742_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__o21ai_1
X_09798_ _04723_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__and2b_1
Xhold1064 datapath.rf.registers\[18\]\[15\] vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 datapath.rf.registers\[26\]\[0\] vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1086 datapath.rf.registers\[6\]\[10\] vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 datapath.rf.registers\[30\]\[23\] vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ _03674_ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ net430 _06176_ _05852_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07289__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _05556_ _05557_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__nor2_1
X_11691_ screen.counter.currentCt\[18\] _06134_ net666 vssd1 vssd1 vccd1 vccd1 _06136_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08635__B _03560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13430_ clknet_leaf_79_clk _00386_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10642_ _05497_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11242__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_100_clk _00346_ net1227 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_10573_ net1416 _03244_ net348 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[1\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12872__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ net1643 net273 net477 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
X_13292_ clknet_leaf_60_clk _00282_ net1266 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09738__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ net273 net1766 net487 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__mux2_1
XANTENNA__11545__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ net2230 _06427_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__xor2_1
XANTENNA__07213__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11125_ _05710_ net1020 vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__nor2_4
X_11056_ net1298 _05702_ net1297 vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__or3b_2
X_10007_ net836 _04499_ _04518_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__nor3_1
XANTENNA__07921__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11958_ net263 net1887 net578 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__mux2_1
XANTENNA__10284__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10909_ net243 net2241 net596 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__mux2_1
X_11889_ net1483 _05874_ net156 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13628_ clknet_leaf_23_clk _00566_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12782__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13559_ clknet_leaf_79_clk _00509_ net1244 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14563__A screen.screenLogic.currentWrx vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07080_ datapath.rf.registers\[20\]\[27\] net803 net753 datapath.rf.registers\[22\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07452__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07204__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout129 _06265_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_2
X_07982_ datapath.rf.registers\[31\]\[7\] net817 net765 datapath.rf.registers\[17\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a22o_1
X_09721_ _02613_ _03377_ _04646_ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a211o_1
X_06933_ datapath.rf.registers\[0\]\[31\] net692 _01859_ _01822_ vssd1 vssd1 vccd1
+ vccd1 _01860_ sky130_fd_sc_hd__o22a_4
XANTENNA__11839__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09652_ net625 _04564_ _04566_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__a31o_1
X_06864_ datapath.rf.registers\[9\]\[31\] net779 net731 datapath.rf.registers\[16\]\[31\]
+ _01790_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a221o_1
XANTENNA__07912__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08603_ net706 _03504_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__or2_1
X_09583_ net333 _04093_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__nor2_1
X_06795_ _01595_ _01597_ _01718_ _01592_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__or4b_1
XANTENNA__12957__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ net518 net517 net406 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ net509 _03018_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout432_A _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ datapath.rf.registers\[0\]\[20\] net693 _02330_ _02342_ vssd1 vssd1 vccd1
+ vccd1 _02343_ sky130_fd_sc_hd__o22a_2
XFILLER_0_135_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ _02702_ _02743_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__or3_1
XANTENNA__07691__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__C _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1282_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ datapath.rf.registers\[18\]\[21\] net790 net763 datapath.rf.registers\[17\]\[21\]
+ _02264_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12692__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07278_ datapath.rf.registers\[10\]\[23\] net918 net858 datapath.rf.registers\[15\]\[23\]
+ _02202_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09017_ _03449_ _03942_ _03943_ _03941_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__o211a_1
XANTENNA__08928__C1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold150 datapath.rf.registers\[0\]\[4\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold161 net98 vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold172 datapath.rf.registers\[0\]\[14\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 datapath.rf.registers\[22\]\[12\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold194 net92 vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10940__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_2
Xfanout641 net642 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_4
Xfanout652 _01724_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_4
X_09919_ _04668_ _04839_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nor2_1
Xfanout663 net665 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_2
XANTENNA__08156__B1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 _03558_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_4
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout696 _01828_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_4
X_12930_ net630 _05669_ _06450_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_70_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ net172 net2435 net555 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__mux2_1
XANTENNA__12867__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11812_ _05647_ net175 _06216_ net178 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12792_ net192 net2175 net563 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07550__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ net1318 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11743_ net1286 net664 _06166_ net713 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14462_ clknet_leaf_52_clk _01349_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11674_ net1534 _06122_ _06124_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13413_ clknet_leaf_89_clk _00369_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11215__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10625_ datapath.PC\[5\] _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__and2_1
X_14530__1352 vssd1 vssd1 vccd1 vccd1 net1352 _14530__1352/LO sky130_fd_sc_hd__conb_1
X_14393_ clknet_leaf_48_clk _01280_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13344_ clknet_leaf_97_clk _00329_ net1220 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_10556_ net1050 _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07434__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ net121 net122 net124 net123 vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__nor4b_1
X_13275_ clknet_leaf_110_clk _00265_ net1107 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11011__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12226_ net211 net2350 net576 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10850__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _06414_ _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ net1285 net1281 net1282 net1284 vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__or4b_1
X_12088_ datapath.mulitply_result\[18\] datapath.multiplication_module.multiplicand_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11039_ _05265_ _05266_ _05271_ _05677_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__nor4_1
XANTENNA__12777__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06580_ net1305 net1303 mmio.memload_or_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ _01510_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_121_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ net646 _03147_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07201_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11206__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08181_ datapath.rf.registers\[25\]\[3\] net796 net762 datapath.rf.registers\[19\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07132_ datapath.rf.registers\[0\]\[26\] _02058_ net828 vssd1 vssd1 vccd1 vccd1 _02059_
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07425__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06804__A _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07063_ net694 _01980_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__or3_1
XANTENNA__06523__B datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07965_ datapath.rf.registers\[17\]\[7\] net880 net852 datapath.rf.registers\[5\]\[7\]
+ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a221o_1
X_09704_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__inv_2
X_06916_ net999 net983 net980 net976 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_52_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07896_ datapath.rf.registers\[14\]\[9\] net800 net779 datapath.rf.registers\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__a22o_1
XANTENNA__08169__C _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _04558_ _04560_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__nor2_1
XANTENNA__12687__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ net973 _01735_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout647_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06778_ _01491_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__nand2b_1
X_09566_ net615 _04485_ _04492_ net676 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ _01625_ _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout814_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ _04422_ _04423_ net337 vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07664__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ _02457_ _02477_ _02522_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_156_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08379_ net696 _03296_ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__nor3_1
XANTENNA__10935__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ _05080_ _05168_ _05244_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__or4_1
XANTENNA__09297__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ net2620 net132 _05880_ net161 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__a22o_1
XANTENNA__07416__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ keypad.decode.sticky\[4\] keypad.decode.sticky\[3\] net1032 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky_n\[3\] sky130_fd_sc_hd__mux2_1
XFILLER_0_61_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10236__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ clknet_leaf_102_clk _00052_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ net392 _04322_ _04323_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08377__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ _06291_ _06292_ _06290_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_72_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11920__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08129__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net463 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_8
Xfanout471 _06454_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
Xfanout482 _06449_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_6
X_13962_ clknet_leaf_11_clk _00849_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout493 _03555_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13063__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ net1636 net247 net546 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
XANTENNA__12597__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ clknet_leaf_92_clk _00780_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12844_ net259 net1869 net553 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12775_ net269 net2079 net563 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__mux2_1
XANTENNA__11006__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14514_ clknet_leaf_33_clk _01401_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11726_ _06076_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07655__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ clknet_leaf_119_clk _01332_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06863__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ screen.counter.currentCt\[5\] screen.counter.currentCt\[6\] _06108_ screen.counter.currentCt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a31o_1
XANTENNA__10845__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ net1512 net346 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[20\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07407__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14376_ clknet_leaf_14_clk _01263_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11588_ _05298_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold908 datapath.rf.registers\[17\]\[30\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ clknet_leaf_76_clk _00317_ net1248 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_10539_ _05402_ _05407_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__nor2_1
XANTENNA__08080__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold919 datapath.rf.registers\[27\]\[21\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13258_ clknet_leaf_65_clk _00248_ net1268 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ _05613_ net1693 net573 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13189_ clknet_leaf_94_clk _00181_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07040__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__A2 _04107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ datapath.rf.registers\[0\]\[12\] _02676_ net827 vssd1 vssd1 vccd1 vccd1 _02677_
+ sky130_fd_sc_hd__mux2_8
X_06701_ _01414_ net1030 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__nor2_1
X_07681_ datapath.rf.registers\[0\]\[14\] net690 _02607_ vssd1 vssd1 vccd1 vccd1 _02608_
+ sky130_fd_sc_hd__o21a_4
XANTENNA__08540__A0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06632_ _01555_ _01556_ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__nor3_1
X_09420_ net329 _04345_ _04346_ _04344_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__a31o_1
XANTENNA__12300__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06563_ datapath.ru.latched_instruction\[30\] _01492_ vssd1 vssd1 vccd1 vccd1 _01493_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _04269_ _04275_ _04276_ _04272_ net675 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_23_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08302_ datapath.rf.registers\[11\]\[1\] net996 _01763_ vssd1 vssd1 vccd1 vccd1 _03229_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09282_ net330 _03850_ _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_118_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06494_ datapath.PC\[7\] vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
XANTENNA__07646__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08233_ datapath.rf.registers\[15\]\[2\] net808 net737 datapath.rf.registers\[8\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06854__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout130_A _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A _05502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08164_ datapath.rf.registers\[30\]\[3\] net987 _01752_ vssd1 vssd1 vccd1 vccd1 _03091_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07115_ datapath.rf.registers\[7\]\[26\] net825 net775 datapath.rf.registers\[11\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a22o_1
XANTENNA__12970__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08095_ datapath.rf.registers\[31\]\[4\] net950 net898 datapath.rf.registers\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07046_ datapath.rf.registers\[3\]\[28\] net965 net862 datapath.rf.registers\[28\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a22o_1
XANTENNA__08359__B1 _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ net363 _03919_ _03920_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_149_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07948_ _02865_ _02872_ _02874_ net831 _01422_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a32o_2
XANTENNA_fanout931_A _01820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ datapath.rf.registers\[17\]\[9\] net881 net865 datapath.rf.registers\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a22o_1
X_09618_ net707 _04544_ net624 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a21o_1
XANTENNA__12210__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _05479_ net630 _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__or3_4
XANTENNA__08196__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09549_ _02260_ _03424_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09087__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ net196 net2010 net450 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _05978_ _05979_ net975 _05917_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__or4bb_1
X_12491_ net219 net2448 net458 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__mux2_1
X_14230_ clknet_leaf_26_clk _01117_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ screen.register.currentXbus\[24\] _05700_ _05707_ screen.register.currentXbus\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a22o_1
XANTENNA__12880__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11373_ _02971_ net669 vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__and2_1
X_14161_ clknet_leaf_27_clk _01048_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08062__A2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10324_ _05035_ _05036_ _05250_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__or3_2
X_13112_ clknet_leaf_39_clk _00104_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09755__A _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07270__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ clknet_leaf_31_clk _00979_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10255_ datapath.PC\[0\] _03286_ _04737_ _04738_ vssd1 vssd1 vccd1 vccd1 _05182_
+ sky130_fd_sc_hd__a22o_1
X_13043_ clknet_leaf_60_clk _00035_ net1267 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09011__A1 _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1200 _00004_ vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_4
Xfanout1222 net1255 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_2
X_10186_ datapath.PC\[10\] net1248 _05109_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_
+ sky130_fd_sc_hd__o22a_1
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10413__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1244 net1245 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1255 net1273 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_2
XANTENNA__08770__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1266 net1267 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__clkbuf_4
Xfanout1277 datapath.PC\[9\] vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_2
Xfanout1288 screen.counter.ct\[14\] vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__clkbuf_2
Xfanout290 _05583_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
Xfanout1299 screen.counter.ct\[2\] vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13945_ clknet_leaf_60_clk _00832_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13876_ clknet_leaf_115_clk _00763_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07876__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09078__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ net186 net2117 net558 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__mux2_1
XANTENNA__10486__D_N net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12758_ net198 net1691 net568 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__mux2_1
XANTENNA__07628__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11709_ net1298 net663 _06146_ net712 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ net1879 net217 net434 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14428_ clknet_leaf_54_clk _01315_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold705 datapath.rf.registers\[15\]\[28\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__A2 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12790__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14359_ clknet_leaf_44_clk _01246_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09250__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap424 _02104_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_2
Xhold716 datapath.rf.registers\[5\]\[28\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 datapath.rf.registers\[20\]\[5\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap435 _06463_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_2
Xhold738 datapath.rf.registers\[22\]\[26\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07261__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold749 datapath.rf.registers\[26\]\[13\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08920_ _02343_ net523 net359 vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06801__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10699__A1 _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11419__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _03336_ _03748_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_71_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07802_ datapath.rf.registers\[26\]\[11\] net940 net696 _02728_ vssd1 vssd1 vccd1
+ vccd1 _02729_ sky130_fd_sc_hd__a211o_1
X_08782_ net368 _03707_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__and3_1
X_07733_ datapath.rf.registers\[31\]\[12\] net817 net759 datapath.rf.registers\[19\]\[12\]
+ _02658_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout178_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ datapath.rf.registers\[18\]\[14\] net912 net896 datapath.rf.registers\[6\]\[14\]
+ _02590_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a221o_1
XANTENNA__07867__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06529__A mmio.memload_or_instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ net492 _04327_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__nand2_1
X_06615_ datapath.ru.latched_instruction\[25\] _01484_ _01486_ datapath.ru.latched_instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a22o_1
XANTENNA__12965__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ _02501_ net521 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout345_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06546_ mmio.key_data\[4\] net1060 _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__o21ai_1
X_09334_ net509 net358 _04260_ net389 vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__a211o_1
XANTENNA__07619__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08816__B2 _03560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06477_ datapath.ru.latched_instruction\[3\] vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
X_09265_ _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08292__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ datapath.rf.registers\[8\]\[2\] net925 net855 datapath.rf.registers\[5\]\[2\]
+ _03142_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09196_ _04119_ _04122_ net413 vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__mux2_1
X_08147_ datapath.rf.registers\[6\]\[3\] net896 _03073_ net696 vssd1 vssd1 vccd1 vccd1
+ _03074_ sky130_fd_sc_hd__a211o_1
XANTENNA__07252__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ datapath.rf.registers\[14\]\[5\] net799 net795 datapath.rf.registers\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout881_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07029_ datapath.rf.registers\[20\]\[28\] net802 net746 datapath.rf.registers\[21\]\[28\]
+ _01953_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a221o_1
XANTENNA__12205__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ _04965_ _04966_ _04472_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__a21oi_1
Xhold10 keypad.debounce.debounce\[4\] vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 keypad.debounce.debounce\[6\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 datapath.multiplication_module.multiplicand_i\[22\] vssd1 vssd1 vccd1 vccd1
+ net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 datapath.rf.registers\[0\]\[13\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 datapath.multiplication_module.multiplicand_i\[11\] vssd1 vssd1 vccd1 vccd1
+ net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 net45 vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 columns.count\[5\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 screen.controlBus\[18\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 screen.controlBus\[28\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _06275_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nor2_1
X_13730_ clknet_leaf_94_clk datapath.multiplication_module.multiplier_i_n\[15\] net1206
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[15\] sky130_fd_sc_hd__dfrtp_1
X_10942_ net241 datapath.rf.registers\[28\]\[16\] net593 vssd1 vssd1 vccd1 vccd1 _00131_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13661_ clknet_leaf_56_clk _00599_ net1257 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_119_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12875__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ net241 net2590 net601 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12612_ net2423 net261 net440 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13592_ clknet_leaf_86_clk _00542_ net1235 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10075__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06818__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ net273 net1777 net451 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11080__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07491__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ net284 net2153 net459 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14213_ clknet_leaf_109_clk _01100_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11425_ _05747_ _05779_ _05783_ _05784_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__and4bb_1
XANTENNA__08035__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ clknet_leaf_46_clk _01031_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11356_ _05863_ _05862_ keypad.apps.app_c\[0\] vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_128_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06902__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10307_ _01621_ _05223_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__o21ai_2
X_14075_ clknet_leaf_52_clk _00962_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11287_ net7 net1046 net1035 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1
+ vccd1 _00301_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ clknet_leaf_33_clk _00018_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ datapath.PC\[14\] net1250 _05163_ _05164_ vssd1 vssd1 vccd1 vccd1 _05165_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10143__B _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_2
XANTENNA__11954__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_4
X_10169_ _04418_ _05095_ _05094_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a21bo_1
Xfanout1052 net1054 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_2
Xfanout1063 _01455_ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_4
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
Xfanout1085 net1125 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 net1102 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ clknet_leaf_13_clk _00815_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_137_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07849__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13859_ clknet_leaf_107_clk _00746_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12785__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07380_ datapath.rf.registers\[11\]\[20\] net776 net761 datapath.rf.registers\[19\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ net672 _03970_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ net646 _02926_ _02907_ net512 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08026__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06639__A_N mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold502 datapath.rf.registers\[12\]\[2\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 datapath.rf.registers\[15\]\[22\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 datapath.mulitply_result\[8\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06812__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 datapath.rf.registers\[13\]\[18\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 datapath.rf.registers\[9\]\[19\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 datapath.rf.registers\[14\]\[8\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 datapath.rf.registers\[18\]\[16\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09127__A2_N net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold579 datapath.rf.registers\[17\]\[9\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net838 _04585_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08903_ _03787_ _03825_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _04702_ _04704_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nand2_1
XANTENNA__08734__A0 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 datapath.rf.registers\[11\]\[13\] vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ _03759_ _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_146_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 datapath.rf.registers\[29\]\[20\] vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1002_A _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 datapath.rf.registers\[26\]\[16\] vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 datapath.rf.registers\[27\]\[29\] vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 datapath.rf.registers\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 datapath.mulitply_result\[1\] vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ _03688_ _03691_ net395 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__mux2_1
Xhold1268 screen.register.currentXbus\[21\] vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout462_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06760__A2 _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1279 net86 vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
X_07716_ datapath.rf.registers\[21\]\[13\] net936 net900 datapath.rf.registers\[20\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
X_08696_ net363 _03621_ _03622_ net375 vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_49_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08177__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12695__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07647_ datapath.rf.registers\[20\]\[14\] net804 net751 datapath.rf.registers\[22\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout727_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07578_ datapath.rf.registers\[12\]\[16\] net890 net859 datapath.rf.registers\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09998__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ net370 _04137_ _04138_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and3_1
X_06529_ mmio.memload_or_instruction\[28\] net1059 vssd1 vssd1 vccd1 vccd1 _01459_
+ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_62_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08265__A2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07473__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ net393 _04174_ _03520_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10943__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ net416 _03879_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__or2_1
X_11210_ net1580 net143 net137 _05092_ vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__a22o_1
XANTENNA__07225__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12190_ _01445_ _06433_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__and2_1
X_11141_ _05678_ _05731_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nor2_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
X_11072_ net1023 _05705_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__nor2_1
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
X_10023_ _01431_ _03785_ net538 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__mux2_1
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11974_ net189 net2310 net580 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
XANTENNA__09150__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[30\]
+ net1259 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ net631 _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or2_4
X_13644_ clknet_leaf_69_clk _00582_ net1228 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ net630 _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13575_ clknet_leaf_87_clk _00525_ net1220 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08256__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ _01514_ net709 _05620_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__o22a_2
XANTENNA__11014__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12526_ net1794 net212 net453 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11949__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08008__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10853__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12457_ net225 net2262 net461 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11408_ screen.register.currentYbus\[23\] net132 _05889_ net161 vssd1 vssd1 vccd1
+ vccd1 _00381_ sky130_fd_sc_hd__a22o_1
XANTENNA__07728__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07216__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12388_ net244 net1783 net469 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
XANTENNA__11563__A2 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ clknet_leaf_5_clk _01014_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11339_ datapath.ru.latched_instruction\[18\] net311 net307 _01495_ vssd1 vssd1 vccd1
+ vccd1 _00341_ sky130_fd_sc_hd__a22o_1
XANTENNA__10154__A _05048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ clknet_leaf_11_clk _00945_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08716__A0 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net1873 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__clkbuf_1
X_06880_ datapath.rf.registers\[3\]\[31\] net965 net962 datapath.rf.registers\[16\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_145_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08278__B net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ net526 net524 net406 vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ _02413_ _02414_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_141_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ _02700_ _03407_ _02701_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07432_ datapath.rf.registers\[23\]\[19\] net786 net766 datapath.rf.registers\[3\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a22o_1
XANTENNA__06807__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07363_ datapath.rf.registers\[2\]\[21\] net921 net881 datapath.rf.registers\[17\]\[21\]
+ _02289_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13347__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ net373 _04027_ _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and3_1
XANTENNA__07455__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11251__B2 _02499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ datapath.rf.registers\[26\]\[22\] net822 net772 datapath.rf.registers\[30\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ net503 net619 net496 net521 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07207__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 datapath.rf.registers\[23\]\[9\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06542__A mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 datapath.rf.registers\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 datapath.rf.registers\[25\]\[23\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 datapath.rf.registers\[24\]\[14\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 datapath.rf.registers\[13\]\[21\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 datapath.rf.registers\[3\]\[26\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 datapath.rf.registers\[31\]\[15\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 datapath.rf.registers\[21\]\[14\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 screen.counter.ct\[19\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _01753_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_4
Xfanout812 _01749_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_4
X_09935_ datapath.PC\[31\] _01728_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__xnor2_1
Xfanout823 _01744_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
Xfanout856 _01853_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
Xfanout867 _01850_ vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_4
X_09866_ _04726_ _04728_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__nand2_1
Xfanout878 _01844_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_4
Xhold1010 datapath.rf.registers\[29\]\[30\] vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 screen.controlBus\[2\] vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07373__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__B1 _04304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 net891 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_4
Xhold1032 datapath.rf.registers\[7\]\[20\] vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net614 _03738_ _03743_ net674 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__o31a_1
Xhold1043 datapath.rf.registers\[4\]\[6\] vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ datapath.PC\[6\] _02972_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout844_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1054 datapath.rf.registers\[14\]\[23\] vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 datapath.rf.registers\[21\]\[31\] vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 datapath.rf.registers\[28\]\[30\] vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 datapath.rf.registers\[16\]\[18\] vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _03670_ _03671_ net365 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__a21o_1
Xhold1098 datapath.rf.registers\[29\]\[26\] vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10938__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ net412 _03604_ _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a21o_1
X_10710_ datapath.PC\[29\] _05549_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__nor2_1
XANTENNA__07694__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _06134_ _06135_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10641_ net1275 _05491_ datapath.PC\[19\] vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08238__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13360_ clknet_leaf_99_clk _00345_ net1224 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07446__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ net1430 _03285_ net348 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[0\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11242__B2 _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12311_ net1548 net277 net476 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13291_ clknet_leaf_60_clk _00281_ net1266 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09738__A2 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ net277 net2041 net484 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__mux2_1
X_12173_ _06427_ _06428_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11124_ _05707_ _05709_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__or3_1
XANTENNA__09763__A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06972__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11055_ net1300 net1301 net1297 net1299 vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__or4_4
XANTENNA__08379__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _04833_ _04835_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__nor2_1
XANTENNA__11009__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ net268 net1907 net578 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
XANTENNA__10848__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ net234 net2193 net594 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__mux2_1
XANTENNA__07730__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11888_ net158 _05873_ net150 screen.controlBus\[7\] vssd1 vssd1 vccd1 vccd1 _00486_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13627_ clknet_leaf_47_clk _00565_ net1197 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10839_ net1976 net234 net602 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07437__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ clknet_leaf_79_clk _00508_ net1244 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11784__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ net1571 net279 net452 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13489_ clknet_leaf_82_clk _00442_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10992__A0 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07981_ datapath.rf.registers\[13\]\[7\] net795 net737 datapath.rf.registers\[8\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a22o_1
XANTENNA__06963__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _02614_ _03409_ _03947_ _03376_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__a31o_1
X_06932_ net694 _01835_ _01846_ _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or4_1
XANTENNA__07905__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09651_ net654 _04577_ _04574_ _04576_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or4b_1
X_06863_ datapath.rf.registers\[5\]\[31\] net784 net756 datapath.rf.registers\[24\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a22o_1
X_08602_ net706 _03504_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__nor2_1
X_09582_ net319 _04506_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a21bo_1
X_06794_ _01597_ net840 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_2
X_08533_ net520 net519 net405 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout160_A _05261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07640__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08464_ _03064_ _03390_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07140__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07132__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07415_ net695 _02332_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__or3_1
XANTENNA__12973__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08395_ _02792_ _02834_ _03320_ _02788_ _02744_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11256__A1_N net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07428__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ datapath.rf.registers\[7\]\[21\] net825 net741 datapath.rf.registers\[1\]\[21\]
+ _02267_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07277_ datapath.rf.registers\[25\]\[23\] net873 net866 datapath.rf.registers\[13\]\[23\]
+ _02194_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09016_ _01632_ _02526_ net687 _02521_ _01634_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A _01757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 datapath.multiplication_module.multiplier_i\[9\] vssd1 vssd1 vccd1 vccd1
+ net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 screen.counter.currentCt\[18\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 datapath.multiplication_module.multiplicand_i\[14\] vssd1 vssd1 vccd1 vccd1
+ net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net41 vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 datapath.rf.registers\[4\]\[0\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07600__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 datapath.rf.registers\[31\]\[0\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A _01806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 _03508_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
XANTENNA__06954__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout631 _05480_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_2
Xfanout642 _03354_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
X_09918_ net1274 datapath.PC\[25\] datapath.PC\[26\] datapath.PC\[27\] net628 vssd1
+ vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__o41a_1
XANTENNA__12213__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 _01623_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_2
Xfanout664 net665 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_2
XANTENNA__09353__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout675 net677 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout686 net687 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09849_ _04668_ _04775_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2b_1
XANTENNA__10241__B _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ net187 net2511 net554 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__mux2_1
X_11811_ net833 _04813_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ net198 net1713 net564 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__mux2_1
X_14530_ net1352 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
X_11742_ net1286 _06072_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xor2_1
XANTENNA__07667__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07131__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11072__B _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14461_ clknet_leaf_24_clk _01348_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11673_ screen.counter.currentCt\[12\] _06122_ net667 vssd1 vssd1 vccd1 vccd1 _06124_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__12883__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13412_ clknet_leaf_89_clk _00368_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10624_ net1278 datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _05482_
+ sky130_fd_sc_hd__and3_1
X_14392_ clknet_leaf_40_clk _01279_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13343_ clknet_leaf_97_clk _00328_ net1220 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10555_ _05449_ _05455_ _05457_ _05434_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ clknet_leaf_110_clk _00264_ net1106 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net121 net122 net123 net124 vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__or4b_1
XFILLER_0_122_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ net214 net2046 net575 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07198__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ datapath.mulitply_result\[29\] datapath.multiplication_module.multiplicand_i\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06945__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__inv_2
X_12087_ datapath.mulitply_result\[18\] datapath.multiplication_module.multiplicand_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ _05679_ _05682_ _05684_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11962__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07370__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ net1504 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07122__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12793__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07200_ _02106_ net531 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_41_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08180_ datapath.rf.registers\[14\]\[3\] net799 net777 datapath.rf.registers\[11\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__a22o_1
XANTENNA__08572__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07131_ datapath.rf.registers\[26\]\[26\] net821 _02054_ _02056_ _02057_ vssd1 vssd1
+ vccd1 vccd1 _02058_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08083__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06804__B _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ _01982_ _01984_ _01986_ _01988_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__or4_1
XANTENNA__07830__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09032__C1 _03958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07189__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07964_ datapath.rf.registers\[19\]\[7\] net944 net904 datapath.rf.registers\[24\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ _02085_ _04542_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nand2_1
X_06915_ datapath.rf.registers\[10\]\[31\] net917 net886 datapath.rf.registers\[9\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12968__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07895_ datapath.rf.registers\[12\]\[9\] net735 net731 datapath.rf.registers\[16\]\[9\]
+ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a221o_1
X_09634_ _04558_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__or2_1
X_06846_ net991 _01733_ _01735_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__and3_4
XANTENNA__07897__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ _03560_ _04486_ _04488_ net610 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a2bb2o_1
X_06777_ datapath.ru.latched_instruction\[12\] _01510_ _01519_ datapath.ru.latched_instruction\[11\]
+ _01463_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout542_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ _01627_ _01631_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07649__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ net398 _04175_ _03516_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__o21a_1
X_08447_ _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout807_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _03298_ _03300_ _03302_ _03304_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__or4_1
XANTENNA__08074__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ _02235_ net527 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__nand2_1
XANTENNA__12208__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09271__C1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10340_ keypad.decode.sticky\[3\] keypad.decode.sticky\[2\] net1032 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky_n\[2\] sky130_fd_sc_hd__mux2_1
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07821__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10951__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ net384 _05197_ _05196_ net394 vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__o211a_1
XANTENNA__09023__C1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12010_ _06290_ _06291_ _06292_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_72_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06927__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_4
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_4
Xfanout472 net475 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_8
X_13961_ clknet_leaf_3_clk _00848_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12878__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout483 _06449_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_2
X_12912_ net1684 net249 net545 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
XANTENNA__07888__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ clknet_leaf_102_clk _00779_ net1121 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07352__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ net262 net2280 net553 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_100_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09629__B2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12774_ net273 net1780 net562 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07104__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14513_ clknet_leaf_8_clk _01400_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11725_ net1293 _06069_ screen.counter.ct\[9\] vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11811__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09488__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444_ clknet_leaf_35_clk _01331_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11656_ net1514 _06110_ _06112_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08065__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ net1495 net346 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[19\]
+ sky130_fd_sc_hd__and2_1
X_14375_ clknet_leaf_24_clk _01262_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11587_ _05763_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__nand2_1
XANTENNA__11022__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13326_ clknet_leaf_76_clk _00316_ net1248 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07812__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10538_ _05445_ _05447_ keypad.alpha vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a21oi_1
Xhold909 datapath.rf.registers\[30\]\[24\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11957__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10861__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ clknet_leaf_65_clk _00247_ net1268 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
X_10469_ _05372_ _05383_ _01636_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a21o_1
X_12208_ net281 net2486 net573 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
XANTENNA__06640__A _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10175__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ clknet_leaf_17_clk _00180_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06918__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _06393_ _06399_ _06398_ _06397_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12788__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ mmio.memload_or_instruction\[13\] net1061 net1027 vssd1 vssd1 vccd1 vccd1
+ _01628_ sky130_fd_sc_hd__and3_1
X_07680_ net696 _02596_ _02600_ _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__or4_1
XANTENNA__07879__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08567__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07343__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ _01557_ _01558_ _01559_ _01560_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09350_ _04269_ _04275_ _04276_ _04272_ net675 vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a32oi_4
X_06562_ net1305 net1303 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ _01492_ sky130_fd_sc_hd__or3b_4
XANTENNA__09096__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08301_ _03215_ _03219_ _03223_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_23_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ net378 _04068_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06493_ datapath.PC\[6\] vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ datapath.rf.registers\[23\]\[2\] net989 _01739_ vssd1 vssd1 vccd1 vccd1 _03159_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_142_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06815__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08163_ datapath.rf.registers\[27\]\[3\] net987 _01763_ vssd1 vssd1 vccd1 vccd1 _03090_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08056__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07114_ datapath.rf.registers\[5\]\[26\] net784 net741 datapath.rf.registers\[1\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a22o_1
XANTENNA__07803__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08094_ datapath.rf.registers\[29\]\[4\] net876 net860 datapath.rf.registers\[28\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07045_ net648 net425 net626 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08359__A1 _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09556__B1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ net367 _03921_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__and3_1
XANTENNA__09308__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _02862_ _02867_ _02873_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__nor3_1
XANTENNA__12698__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__A2 _05383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ datapath.rf.registers\[2\]\[9\] net921 net870 datapath.rf.registers\[27\]\[9\]
+ _02804_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a221o_1
XANTENNA__08531__A1 _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _03431_ _04542_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__xor2_2
X_06829_ _01639_ net998 net982 _01682_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__and4_4
XANTENNA_fanout924_A _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__B _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _03785_ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__nand2_1
XANTENNA__10946__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09479_ net369 _04131_ _04240_ net376 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _05294_ net1014 _05767_ _05297_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ net222 net2186 net457 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11441_ screen.register.currentYbus\[16\] _05775_ _05913_ vssd1 vssd1 vccd1 vccd1
+ _05914_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08598__A1 _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ clknet_leaf_0_clk _01047_ net1070 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11372_ net2536 net133 _05871_ net162 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__a22o_1
XANTENNA__08940__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ clknet_leaf_44_clk _00103_ net1185 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ _05081_ _05166_ _05167_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__or4_1
X_14091_ clknet_leaf_17_clk _00978_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13042_ clknet_leaf_34_clk _00034_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ datapath.PC\[1\] net1245 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__or2_1
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1222 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_2
X_10185_ net204 _05111_ net1309 vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a21o_1
Xfanout1223 net1226 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__A2 _02499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08770__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1245 net1253 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__buf_2
Xfanout1256 net1261 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__clkbuf_4
Xfanout1267 net1273 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_2
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout1278 datapath.PC\[2\] vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
Xfanout1289 screen.counter.ct\[14\] vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__buf_1
XANTENNA__09490__B _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12401__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ clknet_leaf_42_clk _00831_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07325__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13875_ clknet_leaf_59_clk _00762_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11017__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12826_ net189 net2610 net559 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12757_ net212 net1778 net568 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11708_ net1298 _05264_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__xnor2_1
X_12688_ net1965 net224 net433 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
XANTENNA__08038__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14427_ clknet_leaf_21_clk _01314_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _06100_ _06101_ net664 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__and3b_1
XFILLER_0_141_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10157__A _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14358_ clknet_leaf_25_clk _01245_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold706 datapath.rf.registers\[21\]\[27\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold717 datapath.rf.registers\[18\]\[24\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13309_ clknet_leaf_117_clk _00299_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold728 datapath.rf.registers\[18\]\[7\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 datapath.rf.registers\[17\]\[13\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ clknet_leaf_7_clk _01176_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09538__B1 _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10604__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ net706 _03776_ net491 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__o21a_1
XANTENNA__10699__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ datapath.rf.registers\[20\]\[11\] net900 net848 datapath.rf.registers\[1\]\[11\]
+ _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a221o_1
XANTENNA__10323__C _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ net497 net494 _02038_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__a21o_1
XANTENNA__06772__B1 _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ datapath.rf.registers\[26\]\[12\] net820 net770 datapath.rf.registers\[30\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__a22o_1
XANTENNA__12311__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10620__A _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ datapath.rf.registers\[28\]\[14\] net860 net852 datapath.rf.registers\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
X_09402_ net624 _04328_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06614_ datapath.ru.latched_instruction\[15\] _01462_ _01484_ datapath.ru.latched_instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__o22ai_1
XANTENNA__09069__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ _02500_ net521 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ net499 net621 net489 net508 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o211a_1
X_06545_ net1306 net1302 mmio.memload_or_instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ _01475_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout240_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ net675 _04186_ _04188_ _04190_ _04118_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__o41a_2
XFILLER_0_117_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06476_ datapath.ru.latched_instruction\[2\] vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
X_08215_ datapath.rf.registers\[24\]\[2\] net907 net848 datapath.rf.registers\[1\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a22o_1
XANTENNA__08029__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ net341 _03644_ _04120_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout505_A _03146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08146_ datapath.rf.registers\[19\]\[3\] net947 net855 datapath.rf.registers\[5\]\[3\]
+ _03071_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08077_ datapath.rf.registers\[17\]\[5\] net765 net759 datapath.rf.registers\[19\]\[5\]
+ _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__a221o_1
XANTENNA__09529__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07028_ datapath.rf.registers\[30\]\[28\] net771 net760 datapath.rf.registers\[19\]\[28\]
+ _01954_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08201__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 keypad.debounce.debounce\[2\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 datapath.multiplication_module.multiplier_i\[5\] vssd1 vssd1 vccd1 vccd1 net1388
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 datapath.multiplication_module.multiplier_i\[10\] vssd1 vssd1 vccd1 vccd1
+ net1410 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _03414_ _03873_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06763__B1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 net55 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 screen.controlBus\[23\] vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 screen.controlBus\[9\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12221__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 net90 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ datapath.mulitply_result\[2\] datapath.multiplication_module.multiplicand_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__nor2_1
Xhold99 net56 vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07307__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ net246 net1704 net592 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
XANTENNA__10311__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660_ clknet_leaf_57_clk _00598_ net1259 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ net246 net1683 net600 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__mux2_1
X_12611_ net2328 net267 net440 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13591_ clknet_leaf_87_clk _00541_ net1235 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_117_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11361__A _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ net278 net1882 net448 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ net294 net1831 net458 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XANTENNA__12891__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ clknet_leaf_16_clk _01099_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11424_ screen.register.currentYbus\[31\] net132 _05897_ net161 vssd1 vssd1 vccd1
+ vccd1 _00389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _02812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14143_ clknet_leaf_36_clk _01030_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11355_ keypad.apps.app_c\[1\] _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _04619_ _05232_ _05231_ _05229_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__o2bb2a_1
X_14074_ clknet_leaf_21_clk _00961_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11286_ net6 net1044 net1033 mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1
+ vccd1 _00300_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_111_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ clknet_leaf_42_clk _00017_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10237_ net205 _05156_ net1311 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a21o_1
XANTENNA__07546__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_8
Xfanout1031 _01574_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_2
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_4
X_10168_ net834 _04007_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nor2_1
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_1
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_2
Xfanout1086 net1089 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
Xfanout1097 net1098 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_10099_ net837 _05023_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__and3_1
X_13927_ clknet_leaf_20_clk _00814_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11970__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13858_ clknet_leaf_43_clk _00745_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12809_ net268 net1870 net557 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__mux2_1
XANTENNA__10586__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08259__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13789_ clknet_leaf_33_clk _00676_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10066__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09208__C1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08000_ net646 _02926_ _02907_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08580__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 datapath.rf.registers\[20\]\[12\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold514 datapath.rf.registers\[12\]\[18\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12306__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold525 datapath.rf.registers\[25\]\[29\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 datapath.rf.registers\[18\]\[5\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 net69 vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06812__B _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08982__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold558 datapath.rf.registers\[30\]\[7\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _04875_ _04877_ datapath.PC\[30\] net1272 vssd1 vssd1 vccd1 vccd1 _04878_
+ sky130_fd_sc_hd__o2bb2a_1
Xhold569 datapath.rf.registers\[3\]\[31\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06993__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ _03824_ _03826_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ _04786_ _04805_ _04807_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or3_1
XANTENNA__07537__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08833_ net529 net352 _03726_ net388 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a211o_1
Xhold1203 datapath.rf.registers\[6\]\[30\] vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 datapath.rf.registers\[16\]\[31\] vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 datapath.rf.registers\[17\]\[31\] vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1236 net96 vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 screen.register.currentYbus\[0\] vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _03689_ _03690_ net388 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__mux2_1
Xhold1258 datapath.multiplication_module.multiplicand_i\[25\] vssd1 vssd1 vccd1 vccd1
+ net2624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 datapath.rf.registers\[30\]\[30\] vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ datapath.rf.registers\[30\]\[13\] net908 net876 datapath.rf.registers\[29\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12976__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ net362 _03546_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1197_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07646_ datapath.rf.registers\[10\]\[14\] net748 net730 datapath.rf.registers\[16\]\[14\]
+ _02571_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07170__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ datapath.rf.registers\[3\]\[16\] net966 net874 datapath.rf.registers\[25\]\[16\]
+ _02503_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ net361 _04239_ _04242_ net373 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__o211a_1
X_06528_ mmio.key_data\[0\] mmio.memload_or_instruction\[0\] net1059 vssd1 vssd1 vccd1
+ vccd1 _01458_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ net384 _03686_ _03524_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ net336 _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout991_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08129_ datapath.rf.registers\[6\]\[4\] net814 net766 datapath.rf.registers\[3\]\[4\]
+ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__a221o_1
XANTENNA__12216__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ net1023 _05728_ net1021 _05725_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11309__A0 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XANTENNA__06984__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
X_11071_ net1300 net1301 net1299 net1297 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__or4b_4
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
X_10022_ net837 _03785_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__or2_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ net194 net2596 net580 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XANTENNA__09150__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ _05478_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__or2_1
X_13712_ clknet_leaf_57_clk datapath.multiplication_module.multiplicand_i_n\[29\]
+ net1259 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07161__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07700__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10855_ _05479_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__or2_1
X_13643_ clknet_leaf_69_clk _00581_ net1229 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ clknet_leaf_87_clk _00524_ net1219 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10599__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ datapath.mulitply_result\[9\] net428 net658 vssd1 vssd1 vccd1 vccd1 _05621_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09453__A2 _04367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12525_ net1747 net213 net453 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12456_ net231 net2015 net462 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11407_ _02191_ _05695_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12387_ net236 net1960 net468 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ clknet_leaf_116_clk _01013_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07767__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11338_ datapath.ru.latched_instruction\[17\] net311 net307 _01479_ vssd1 vssd1 vccd1
+ vccd1 _00340_ sky130_fd_sc_hd__a22o_1
XANTENNA__06975__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ clknet_leaf_2_clk _00944_ net1075 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11269_ mmio.wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__and2_1
XANTENNA__07519__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__A1 _03087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ net2411 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07463__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire423_A _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12796__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10287__A0 _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ datapath.rf.registers\[10\]\[18\] net917 net870 datapath.rf.registers\[27\]\[18\]
+ _02426_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_18_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08480_ _03405_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07431_ _02351_ _02353_ _02355_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08294__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06807__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07362_ datapath.rf.registers\[20\]\[21\] net901 net889 datapath.rf.registers\[12\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ _04023_ _04024_ net366 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07293_ datapath.rf.registers\[14\]\[22\] net801 net764 datapath.rf.registers\[17\]\[22\]
+ _02219_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09032_ _02568_ net683 _03948_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 datapath.rf.registers\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 datapath.rf.registers\[15\]\[25\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout203_A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold322 datapath.rf.registers\[19\]\[4\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 datapath.rf.registers\[30\]\[4\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 datapath.rf.registers\[7\]\[25\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 datapath.mulitply_result\[21\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 datapath.rf.registers\[21\]\[9\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10762__A1 datapath.mulitply_result\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 datapath.rf.registers\[22\]\[10\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 datapath.rf.registers\[12\]\[17\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net803 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
Xhold399 datapath.rf.registers\[7\]\[3\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09934_ _04858_ _04859_ _04856_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__o21ai_1
Xfanout813 net816 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_4
Xfanout824 _01740_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_8
Xfanout835 net838 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 _01719_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
Xfanout857 _01853_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _04790_ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__nand2_1
Xhold1000 datapath.rf.registers\[10\]\[6\] vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 _01848_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
XANTENNA_fanout572_A _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout879 _01844_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
Xhold1011 datapath.rf.registers\[17\]\[29\] vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 datapath.rf.registers\[20\]\[17\] vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1033 datapath.rf.registers\[11\]\[18\] vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net610 _03731_ _03720_ _03560_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__o2bb2a_1
X_09796_ datapath.PC\[6\] _02972_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__and2_1
Xhold1044 datapath.rf.registers\[0\]\[9\] vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1055 datapath.rf.registers\[28\]\[22\] vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1066 datapath.rf.registers\[31\]\[9\] vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 datapath.rf.registers\[30\]\[26\] vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _03672_ _03673_ net362 vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a21o_1
Xhold1088 datapath.rf.registers\[2\]\[5\] vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 datapath.rf.registers\[15\]\[23\] vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__A1 _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ net413 net341 _03471_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__and3_1
XANTENNA__07143__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__S net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ datapath.rf.registers\[23\]\[15\] net933 net878 datapath.rf.registers\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a22o_1
X_10640_ net1275 datapath.PC\[19\] _05491_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10954__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _05413_ _05432_ _05475_ _05477_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[4\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ net2409 net280 net476 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
X_13290_ clknet_leaf_112_clk _00280_ net1103 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12241_ net280 net2472 net484 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__mux2_1
XANTENNA__09199__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07749__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net2531 _06426_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11123_ _05705_ net1020 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ net1022 _05703_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__nor2_2
X_10005_ _04920_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07382__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__A2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output122_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11814__A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ net271 net2432 net580 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__mux2_1
XANTENNA__07134__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10907_ net238 net1641 net597 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__mux2_1
X_11887_ net157 _05872_ net150 net2256 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _05664_ _05663_ net711 _01479_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__o2bb2a_2
X_13626_ clknet_leaf_40_clk _00564_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13557_ clknet_leaf_79_clk _00507_ net1244 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10769_ _01457_ net709 _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__o21a_2
XANTENNA__10864__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ net2366 net280 net452 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__mux2_1
X_13488_ clknet_leaf_83_clk _00441_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12439_ net293 net1660 net460 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ clknet_leaf_23_clk _00996_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_07980_ net646 _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__nand2_1
X_06931_ _01849_ _01852_ _01854_ _01857_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__or4_1
X_09650_ net339 _04021_ net316 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_143_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06862_ datapath.rf.registers\[8\]\[31\] net738 net715 datapath.rf.registers\[29\]\[31\]
+ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a221o_1
X_08601_ net398 _03527_ _03516_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__o21a_1
XANTENNA__07912__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ _02126_ net685 net681 _02127_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__o221a_1
X_06793_ _01595_ _01718_ _01592_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__or3b_2
XANTENNA__09114__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _03288_ _03446_ _03457_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_46_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07125__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08463_ _03125_ _03388_ _03123_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout153_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06537__B _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ _02334_ _02336_ _02338_ _02340_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__or4_1
X_08394_ _02793_ _02835_ _03320_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__or3b_1
XFILLER_0_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ datapath.rf.registers\[19\]\[21\] net760 net735 datapath.rf.registers\[12\]\[21\]
+ _02266_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1062_A _01455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
X_07276_ datapath.rf.registers\[8\]\[23\] net926 net905 datapath.rf.registers\[24\]\[23\]
+ _02195_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a221o_1
XANTENNA__06553__A mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09015_ net419 _03648_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold130 keypad.decode.push vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 datapath.multiplication_module.multiplier_i\[14\] vssd1 vssd1 vccd1 vccd1
+ net1507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__A1 _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 net43 vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 datapath.rf.registers\[22\]\[0\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 datapath.rf.registers\[0\]\[6\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold185 datapath.multiplication_module.multiplicand_i\[15\] vssd1 vssd1 vccd1 vccd1
+ net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 datapath.multiplication_module.multiplicand_i\[3\] vssd1 vssd1 vccd1 vccd1
+ net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_2
Xfanout621 _03508_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_2
Xfanout632 _04677_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
X_09917_ _04842_ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nand2_1
Xfanout654 _01623_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout665 _06099_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08156__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net677 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_13_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ datapath.PC\[25\] net628 _04773_ _04774_ _04669_ vssd1 vssd1 vccd1 vccd1
+ _04775_ sky130_fd_sc_hd__a221o_1
Xfanout687 _03495_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07364__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout698 net699 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ net632 _04705_ net1276 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _06215_ datapath.PC\[13\] net306 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ net209 net2083 net564 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__mux2_1
XANTENNA__07116__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11741_ screen.counter.ct\[15\] net664 _06165_ net713 vssd1 vssd1 vccd1 vccd1 _00438_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10120__C1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11672_ _06122_ _06123_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__nor2_1
X_14460_ clknet_leaf_57_clk _01347_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13411_ clknet_leaf_89_clk _00367_ net1214 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10623_ _05478_ _05479_ net631 vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10684__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14391_ clknet_leaf_50_clk _01278_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13342_ clknet_leaf_97_clk _00327_ net1220 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_10554_ net1026 _05459_ _05402_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13273_ clknet_leaf_110_clk _00263_ net1106 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
X_10485_ keypad.apps.button\[0\] net1032 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09774__A _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ net219 net2243 net576 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12155_ datapath.mulitply_result\[29\] datapath.multiplication_module.multiplicand_i\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__and2_1
XANTENNA__12404__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11106_ net1292 net1293 screen.counter.ct\[11\] screen.counter.ct\[10\] vssd1 vssd1
+ vccd1 vccd1 _05756_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_9_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12086_ net321 _06355_ _06356_ net325 net1853 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_88_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08147__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ _05313_ _05322_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_108_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07107__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06638__A _01456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ net1936 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11939_ net152 _05891_ net127 screen.register.currentXbus\[25\] vssd1 vssd1 vccd1
+ vccd1 _00536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08607__A0 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ clknet_leaf_20_clk _00547_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_07130_ _02043_ _02044_ _02051_ _02053_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__or4_1
XANTENNA__10607__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08291__C _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07061_ datapath.rf.registers\[14\]\[28\] net893 net889 datapath.rf.registers\[12\]\[28\]
+ _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a221o_1
XANTENNA__06538__C_N mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11914__B1 _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06820__B _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ datapath.rf.registers\[31\]\[7\] net948 net856 datapath.rf.registers\[15\]\[7\]
+ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_79_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06914_ net1002 net983 net981 _01801_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__and4_4
X_09702_ _01800_ _01861_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__and2_1
X_07894_ datapath.rf.registers\[3\]\[9\] net767 net749 datapath.rf.registers\[10\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a22o_1
XANTENNA__07346__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06845_ net993 _01743_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__and2_4
X_09633_ _04546_ _04555_ _04559_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout368_A _03540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _01717_ _04476_ net625 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__o21ai_1
X_06776_ datapath.ru.latched_instruction\[26\] _01613_ _01702_ vssd1 vssd1 vccd1 vccd1
+ _01703_ sky130_fd_sc_hd__a21o_1
XANTENNA__09099__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _03352_ net688 _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _04162_ _04179_ net399 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ _02457_ _02477_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ datapath.rf.registers\[20\]\[0\] net903 net852 datapath.rf.registers\[5\]\[0\]
+ _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07328_ datapath.rf.registers\[0\]\[22\] net693 _02242_ _02254_ vssd1 vssd1 vccd1
+ vccd1 _02255_ sky130_fd_sc_hd__o22a_2
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07259_ datapath.rf.registers\[31\]\[23\] net818 net760 datapath.rf.registers\[19\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ _03207_ _03146_ net353 vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__mux2_1
XANTENNA__11905__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12224__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 net443 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08003__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _06459_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_8
X_13960_ clknet_leaf_12_clk _00847_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07337__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout484 net487 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_6
Xfanout495 _03544_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_2
X_12911_ net2224 net255 net545 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
X_13891_ clknet_leaf_105_clk _00778_ net1101 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12842_ net267 net2128 net553 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11436__A2 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12773_ net279 net2094 net562 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__mux2_1
XANTENNA__12894__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14512_ clknet_leaf_3_clk _01399_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ net1293 net663 _06155_ net712 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11655_ screen.counter.currentCt\[6\] _06110_ net667 vssd1 vssd1 vccd1 vccd1 _06112_
+ sky130_fd_sc_hd__o21ai_1
X_14443_ clknet_leaf_101_clk _01330_ net1223 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06863__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10606_ net2283 net346 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[18\]
+ sky130_fd_sc_hd__and2_1
X_11586_ _05750_ _06046_ _06047_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__or4_1
X_14374_ clknet_leaf_111_clk _01261_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10537_ _05399_ net1026 _05446_ _05442_ net1050 vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__o32a_1
X_13325_ clknet_leaf_117_clk _00315_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13256_ clknet_leaf_65_clk _00246_ net1269 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09014__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10468_ _05378_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ net284 net2304 net574 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
X_13187_ clknet_leaf_103_clk _00179_ net1121 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10399_ _05315_ _05316_ _05317_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__o211a_1
XANTENNA__06640__B _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ _06397_ _06398_ _06399_ _06393_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a211o_1
XANTENNA__07040__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11255__A1_N net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ datapath.mulitply_result\[15\] datapath.multiplication_module.multiplicand_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_06630_ datapath.ru.latched_instruction\[8\] datapath.ru.latched_instruction\[9\]
+ datapath.ru.latched_instruction\[10\] datapath.ru.latched_instruction\[11\] vssd1
+ vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08286__C _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ datapath.ru.latched_instruction\[4\] _01476_ _01490_ vssd1 vssd1 vccd1 vccd1
+ _01491_ sky130_fd_sc_hd__o21ai_1
X_08300_ datapath.rf.registers\[24\]\[1\] net758 _03224_ _03225_ _03226_ vssd1 vssd1
+ vccd1 vccd1 _03227_ sky130_fd_sc_hd__a2111o_1
X_09280_ net383 _04205_ _04206_ net332 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__a31o_1
X_06492_ datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
XANTENNA__07500__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ datapath.rf.registers\[11\]\[2\] net994 _01763_ vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_118_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06854__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__B _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08162_ datapath.rf.registers\[0\]\[3\] net830 vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07113_ _02018_ net532 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_151_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06606__A2 _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ net509 _03018_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07044_ datapath.rf.registers\[0\]\[28\] net828 _01970_ vssd1 vssd1 vccd1 vccd1 _01971_
+ sky130_fd_sc_hd__o21ai_2
XANTENNA__06831__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07567__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net497 net494 net521 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout485_A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ datapath.rf.registers\[6\]\[8\] net815 net794 datapath.rf.registers\[13\]\[8\]
+ _02858_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a221o_1
XANTENNA__07319__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07877_ datapath.rf.registers\[7\]\[9\] net957 net930 datapath.rf.registers\[4\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a22o_1
X_09616_ _03345_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__xnor2_1
X_06828_ net990 _01754_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__and2_2
X_06759_ _01415_ net1004 _01661_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__and3_1
X_09547_ _03831_ _03871_ _04472_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout917_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09478_ _04249_ _04250_ net382 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08429_ _01620_ _01633_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12219__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11440_ screen.register.currentXbus\[0\] _05704_ _05776_ screen.register.currentYbus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10962__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _03017_ _05695_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__and2_1
X_10322_ _05237_ _05242_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or2_1
X_13110_ clknet_leaf_26_clk _00102_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07837__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14090_ clknet_leaf_10_clk _00977_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07270__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ clknet_leaf_27_clk _00033_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__inv_2
XANTENNA__07558__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_2
X_10184_ _04805_ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__nand2_1
Xfanout1213 net1216 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12889__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1224 net1226 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
Xfanout1235 net1254 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__buf_2
Xfanout1246 net1253 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_4
Xfanout1257 net1261 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1268 net1269 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__clkbuf_4
Xfanout270 net272 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1279 screen.counter.ct\[21\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_2
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
Xfanout292 _05590_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
X_13943_ clknet_leaf_44_clk _00830_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11094__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13874_ clknet_leaf_34_clk _00761_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12825_ net194 net2233 net558 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07089__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ net216 net2488 net567 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__mux2_1
XANTENNA__08607__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ net1300 net663 _06145_ net712 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a22o_1
X_12687_ net1749 net232 net434 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14426_ clknet_leaf_51_clk _01313_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11638_ screen.counter.currentCt\[0\] _06087_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11968__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14357_ clknet_leaf_29_clk _01244_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10872__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11569_ _05307_ _06033_ _05734_ _05746_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07797__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 datapath.rf.registers\[25\]\[31\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_75_clk _00298_ net1250 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold718 datapath.rf.registers\[23\]\[7\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08994__C1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07261__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold729 datapath.rf.registers\[4\]\[25\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ clknet_leaf_4_clk _01175_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13239_ clknet_leaf_75_clk _00229_ net1251 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__A1 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ datapath.rf.registers\[11\]\[11\] net968 net924 datapath.rf.registers\[8\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
X_08780_ net502 net618 net496 net533 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08578__A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ datapath.rf.registers\[20\]\[12\] net804 net717 datapath.rf.registers\[29\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08297__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ datapath.rf.registers\[10\]\[14\] net916 net856 datapath.rf.registers\[15\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
XANTENNA__07721__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06613_ _01537_ _01538_ _01540_ _01542_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__or4_1
X_09401_ _04312_ _04327_ net688 vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07593_ datapath.rf.registers\[0\]\[16\] net693 _02507_ _02519_ vssd1 vssd1 vccd1
+ vccd1 _02520_ sky130_fd_sc_hd__o22a_1
X_06544_ datapath.ru.latched_instruction\[8\] _01472_ _01473_ datapath.ru.latched_instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__o22ai_2
X_09332_ net505 _03087_ net353 vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09263_ net624 _04183_ _04189_ _01622_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06475_ datapath.ru.latched_instruction\[1\] vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout233_A _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08214_ datapath.rf.registers\[22\]\[2\] net955 net919 datapath.rf.registers\[10\]\[2\]
+ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ net341 _03644_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__a21oi_1
X_08145_ datapath.rf.registers\[7\]\[3\] net959 net851 datapath.rf.registers\[1\]\[3\]
+ _03069_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1142_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08076_ datapath.rf.registers\[20\]\[5\] net804 net769 datapath.rf.registers\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_1
XANTENNA__07252__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07027_ datapath.rf.registers\[15\]\[28\] net806 net749 datapath.rf.registers\[10\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold1250_A mmio.memload_or_instruction\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11336__A1 _01461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold12 keypad.debounce.debounce\[14\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 keypad.debounce.debounce\[10\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08752__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 keypad.apps.button\[2\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net613 _03882_ _03904_ net674 vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__o31a_1
Xhold45 datapath.multiplication_module.multiplicand_i\[4\] vssd1 vssd1 vccd1 vccd1
+ net1411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 screen.counter.ct\[5\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 net47 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 datapath.multiplication_module.multiplier_i\[12\] vssd1 vssd1 vccd1 vccd1
+ net1444 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ datapath.rf.registers\[17\]\[8\] net764 net757 datapath.rf.registers\[24\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a22o_1
Xhold89 net88 vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ net251 net2112 net590 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__mux2_1
XANTENNA__07712__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10311__A2 _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ net251 net2180 net598 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__mux2_1
XANTENNA__10957__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ net1933 net269 net441 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__mux2_1
X_13590_ clknet_leaf_79_clk _00540_ net1243 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ net280 net2566 net448 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__mux2_1
XANTENNA__06818__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12472_ net292 net2490 net459 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XANTENNA__07491__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14211_ clknet_leaf_104_clk _01098_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11423_ _01799_ net669 vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07779__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ keypad.apps.app_c\[0\] keypad.apps.app_c\[1\] _05835_ _05861_ keypad.apps.button\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_105_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14142_ clknet_leaf_51_clk _01029_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10305_ net625 net680 net492 net676 vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07286__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ net5 net1044 net1033 mmio.memload_or_instruction\[12\] vssd1 vssd1 vccd1
+ vccd1 _00299_ sky130_fd_sc_hd__o22a_1
X_14073_ clknet_leaf_48_clk _00960_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09782__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ net202 _05160_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__and3_1
X_13024_ clknet_leaf_50_clk _00016_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1010 _01581_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 _05732_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
Xfanout1032 _01450_ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__buf_2
X_10167_ net701 _04420_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nand2_1
XANTENNA__12412__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1043 _01454_ vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
Xfanout1054 _03568_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_2
Xfanout1065 net1076 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_4
Xfanout1076 net1125 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_2
Xfanout1087 net1089 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_2
X_10098_ _03586_ _05024_ net1052 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__a21o_1
Xfanout1098 net1102 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09153__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10838__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ clknet_leaf_108_clk _00813_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13434__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13857_ clknet_leaf_41_clk _00744_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10867__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12808_ net271 net1787 net558 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__mux2_1
X_13788_ clknet_leaf_58_clk _00675_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11263__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12739_ net281 net2425 net565 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ clknet_leaf_2_clk _01296_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold504 datapath.rf.registers\[19\]\[10\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold515 datapath.rf.registers\[19\]\[29\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold526 datapath.rf.registers\[6\]\[16\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06812__C _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold537 datapath.rf.registers\[9\]\[8\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 datapath.rf.registers\[28\]\[9\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold559 datapath.rf.registers\[5\]\[23\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net207 _04876_ net1312 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a21oi_1
X_08901_ net615 _03799_ _03827_ net676 vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ _04805_ _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08832_ net527 net354 _03758_ net386 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a211o_1
XANTENNA__12322__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1204 datapath.rf.registers\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 datapath.mulitply_result\[5\] vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 datapath.rf.registers\[31\]\[22\] vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 screen.counter.currentCt\[3\] vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 screen.register.currentXbus\[3\] vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ net529 net531 net353 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__mux2_1
Xhold1259 datapath.rf.registers\[23\]\[20\] vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout183_A _05579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07714_ datapath.rf.registers\[18\]\[13\] net912 net864 datapath.rf.registers\[13\]\[13\]
+ _02638_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a221o_1
X_08694_ _01904_ net534 net359 vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10777__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ datapath.rf.registers\[8\]\[14\] net738 net717 datapath.rf.registers\[29\]\[14\]
+ _02570_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout350_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ datapath.rf.registers\[16\]\[16\] net963 net915 datapath.rf.registers\[18\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a22o_1
XANTENNA__09447__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11181__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06527_ mmio.key_data\[6\] mmio.memload_or_instruction\[6\] net1060 vssd1 vssd1 vccd1
+ vccd1 _01457_ sky130_fd_sc_hd__mux2_2
XANTENNA__11254__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09998__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ _04237_ _04238_ net365 vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_62_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09246_ net399 _04172_ _04163_ net336 vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07473__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09177_ net398 _03891_ _03516_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__o21ai_1
X_08128_ datapath.rf.registers\[26\]\[4\] net820 net738 datapath.rf.registers\[8\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__a22o_1
XANTENNA__07225__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08059_ datapath.rf.registers\[19\]\[5\] net944 net856 datapath.rf.registers\[15\]\[5\]
+ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
X_11070_ net1022 _05717_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__nor2_4
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
X_10021_ datapath.PC\[21\] _03583_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08725__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__B1 _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net198 net1653 net581 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_57_clk datapath.multiplication_module.multiplicand_i_n\[28\]
+ net1258 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10296__A1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ _01643_ _01666_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10687__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13642_ clknet_leaf_69_clk _00580_ net1228 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10854_ _01650_ _01669_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10048__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11245__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__C1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13573_ clknet_leaf_87_clk _00523_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ _04116_ _05619_ net846 vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11796__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12524_ net1911 net218 net453 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12455_ net226 net2013 net461 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12407__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11311__S _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11406_ screen.register.currentYbus\[22\] net133 _05888_ net162 vssd1 vssd1 vccd1
+ vccd1 _00380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07216__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ net240 net1892 net470 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14125_ clknet_leaf_119_clk _01012_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11337_ _01511_ net1028 net307 net311 datapath.ru.latched_instruction\[16\] vssd1
+ vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__a32o_1
X_14056_ clknet_leaf_14_clk _00943_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11268_ net1415 net140 net134 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__a21o_1
X_13007_ net2343 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__clkbuf_1
X_10219_ net1277 _04116_ net536 vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__mux2_1
XANTENNA__10451__A _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ net2144 net144 net137 _05236_ vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__a22o_1
XANTENNA__07924__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10287__A1 _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ clknet_leaf_28_clk _00796_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07430_ datapath.rf.registers\[26\]\[19\] net821 net752 datapath.rf.registers\[22\]\[19\]
+ _02356_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11236__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06807__C _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07361_ datapath.rf.registers\[11\]\[21\] net970 _02283_ _02285_ _02287_ vssd1 vssd1
+ vccd1 vccd1 _02288_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08101__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09100_ _04025_ _04026_ net361 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a21o_1
XANTENNA__07455__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07292_ datapath.rf.registers\[23\]\[22\] net788 net724 datapath.rf.registers\[27\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09031_ _03474_ net318 _03957_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_142_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12317__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06823__B _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07207__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold301 datapath.rf.registers\[26\]\[9\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 datapath.rf.registers\[22\]\[28\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 datapath.rf.registers\[5\]\[25\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 datapath.rf.registers\[17\]\[15\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 datapath.rf.registers\[13\]\[25\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold356 datapath.rf.registers\[25\]\[4\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10762__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold367 datapath.rf.registers\[30\]\[12\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 datapath.rf.registers\[22\]\[4\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 datapath.rf.registers\[27\]\[12\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _04858_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__xor2_2
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_4
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_4
Xfanout825 _01740_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
Xfanout836 net838 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
Xfanout847 _01599_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
X_09864_ _04741_ _04743_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06718__A1 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout858 _01853_ vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_4
Xfanout869 _01848_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1105_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 datapath.rf.registers\[24\]\[26\] vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 datapath.rf.registers\[4\]\[5\] vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A2 _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ net706 _03705_ net623 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__a21oi_1
Xhold1023 datapath.rf.registers\[29\]\[31\] vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _04720_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__and2b_1
Xhold1034 datapath.rf.registers\[6\]\[21\] vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout565_A _06465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1045 datapath.rf.registers\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 datapath.rf.registers\[1\]\[30\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 datapath.rf.registers\[6\]\[15\] vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net497 net494 net533 vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__a21o_1
Xhold1078 datapath.rf.registers\[6\]\[3\] vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1089 datapath.rf.registers\[12\]\[3\] vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_37_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _03468_ _03470_ net408 vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__mux2_1
X_07628_ datapath.rf.registers\[2\]\[15\] net921 net862 datapath.rf.registers\[28\]\[15\]
+ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a221o_1
XANTENNA__07694__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ datapath.rf.registers\[6\]\[16\] net815 net785 datapath.rf.registers\[5\]\[16\]
+ _02485_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a221o_1
X_10570_ _01444_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__nand2_1
XANTENNA__07446__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ net334 _04155_ _04146_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12227__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12240_ net286 net2454 net487 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__mux2_1
XANTENNA__09199__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ columns.count\[0\] _06426_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11122_ _05706_ net1020 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_92_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold890 screen.controlBus\[6\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11367__A _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ _05701_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__or2_1
XANTENNA__07906__A0 _02831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ _01432_ net1312 _04928_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_95_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10269__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ net275 net2123 net579 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ net245 datapath.rf.registers\[27\]\[15\] net596 vssd1 vssd1 vccd1 vccd1 _00098_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11886_ net157 _05871_ net150 net2605 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ clknet_leaf_45_clk _00563_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10837_ datapath.mulitply_result\[17\] net428 net662 vssd1 vssd1 vccd1 vccd1 _05664_
+ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ clknet_leaf_88_clk _00506_ net1219 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07437__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ datapath.mulitply_result\[6\] net426 _05603_ _05605_ datapath.MemRead vssd1
+ vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12507_ net1741 net286 net455 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__mux2_1
XANTENNA__10446__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ clknet_leaf_82_clk _00440_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ _01512_ net710 _05546_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12438_ net297 net2356 net460 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10880__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ _05666_ net577 _06450_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__or3_1
XANTENNA__10744__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14108_ clknet_leaf_54_clk _00995_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07070__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09347__C1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ datapath.rf.registers\[5\]\[31\] net853 net849 datapath.rf.registers\[1\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
X_14039_ clknet_leaf_44_clk _00926_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08289__C _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06861_ datapath.rf.registers\[23\]\[31\] net787 net747 datapath.rf.registers\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a22o_1
X_08600_ net393 _03526_ _03520_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__o21a_1
X_06792_ _01595_ _01718_ _01592_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nor3b_1
X_09580_ _03449_ _04107_ _04500_ net679 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__o22a_1
X_08531_ _03288_ _03446_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08322__B1 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08462_ _03181_ _03387_ _03180_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07676__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11209__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ datapath.rf.registers\[30\]\[20\] net911 net882 datapath.rf.registers\[17\]\[20\]
+ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08393_ _02885_ _03318_ _02836_ _02880_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__a211o_1
XANTENNA__06884__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout146_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ datapath.rf.registers\[3\]\[21\] net767 net756 datapath.rf.registers\[24\]\[21\]
+ _02265_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a221o_1
XANTENNA__07428__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07275_ datapath.rf.registers\[9\]\[23\] net886 net878 datapath.rf.registers\[29\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout313_A _05859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1055_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09014_ _02500_ net521 net684 vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold120 net77 vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _00211_ vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1222_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 screen.counter.currentCt\[20\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 net91 vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07061__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 datapath.rf.registers\[0\]\[21\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold175 datapath.rf.registers\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 datapath.rf.registers\[26\]\[3\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 datapath.multiplication_module.multiplicand_i\[12\] vssd1 vssd1 vccd1 vccd1
+ net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
Xfanout611 _03562_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
X_09916_ datapath.PC\[28\] net628 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__or2_1
Xfanout622 _03508_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_2
Xfanout633 _04677_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_1
Xfanout655 _01622_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_2
Xfanout666 _06088_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_2
Xfanout677 _03557_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_2
X_09847_ datapath.PC\[25\] net628 vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__xor2_2
Xfanout688 _03355_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout699 net703 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_2
XANTENNA__08561__A0 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12510__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _01627_ _04678_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08729_ net517 _02742_ net404 vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ screen.counter.ct\[15\] _06084_ _06072_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07667__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11671_ screen.counter.currentCt\[11\] _06120_ net667 vssd1 vssd1 vccd1 vccd1 _06123_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__10965__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13410_ clknet_leaf_88_clk _00366_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10622_ _01602_ _01621_ net839 _01664_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a31o_1
X_14390_ clknet_leaf_24_clk _01277_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ clknet_leaf_97_clk _00326_ net1220 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_10553_ _05458_ _05461_ _01444_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13272_ clknet_leaf_112_clk _00262_ net1094 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
X_10484_ screen.register.controlFill screen.register.xFill _05395_ vssd1 vssd1 vccd1
+ vccd1 screen.screenEdge.enableIn sky130_fd_sc_hd__and3_1
X_12223_ net223 net2597 net575 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__mux2_1
XANTENNA__07052__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _06407_ _06411_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__nand2_1
X_11105_ net1284 net1285 _05271_ _05751_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_9_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12085_ _06353_ _06354_ _06352_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11036_ net1292 net1285 _05686_ net1012 vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a31o_1
XANTENNA__08001__C1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08552__A0 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12420__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10489__D_N net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12987_ net1540 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06638__B _01464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ net152 _05890_ net127 net2585 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06866__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10875__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ net202 _04863_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13608_ clknet_leaf_114_clk _00546_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08607__A1 _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13539_ clknet_leaf_88_clk _00489_ net1211 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08083__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07060_ datapath.rf.registers\[6\]\[28\] net897 net865 datapath.rf.registers\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_136_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07291__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11390__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ datapath.rf.registers\[1\]\[7\] net848 _02888_ net696 vssd1 vssd1 vccd1 vccd1
+ _02889_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09701_ _03440_ _04586_ _04625_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__and3_1
X_06913_ datapath.rf.registers\[14\]\[31\] net893 net889 datapath.rf.registers\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08543__A0 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ datapath.rf.registers\[26\]\[9\] net821 net715 datapath.rf.registers\[29\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09632_ net493 _04543_ _04557_ net677 vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a211o_1
X_06844_ net991 _01733_ _01741_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__and3_1
XANTENNA__12330__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07897__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06829__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09563_ _01717_ _04489_ net493 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a21o_1
X_06775_ datapath.ru.latched_instruction\[29\] _01616_ _01627_ datapath.ru.latched_instruction\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a22o_1
X_08514_ net706 _03440_ net623 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__a21o_1
XANTENNA__07649__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ _02614_ _03326_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10102__B1 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06857__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ _02370_ net523 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10785__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10694__A1_N _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout528_A _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ datapath.rf.registers\[19\]\[0\] net947 net913 datapath.rf.registers\[18\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a22o_1
XANTENNA__06609__B1 _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07327_ _02237_ _02238_ _02251_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__or4_1
XANTENNA__08074__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07282__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ datapath.rf.registers\[6\]\[23\] net814 net806 datapath.rf.registers\[15\]\[23\]
+ _02184_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07821__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12505__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ datapath.rf.registers\[21\]\[25\] net939 net931 datapath.rf.registers\[4\]\[25\]
+ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07034__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 datapath.MUL_EN vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 net443 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_4
Xfanout452 net455 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 _06456_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08534__A0 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2_N net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 net487 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_8
X_12910_ net1549 net260 net545 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
Xfanout496 _03543_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
XANTENNA__12240__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ clknet_leaf_43_clk _00777_ net1185 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07888__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ net270 net2044 net554 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
X_14548__1359 vssd1 vssd1 vccd1 vccd1 net1359 _14548__1359/LO sky130_fd_sc_hd__conb_1
XANTENNA__06560__A2 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ net281 net2132 net561 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14511_ clknet_leaf_3_clk _01398_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11723_ net1293 _06069_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10695__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14442_ clknet_leaf_10_clk _01329_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11654_ _06110_ _06111_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ net1485 net346 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[17\]
+ sky130_fd_sc_hd__and2_1
X_14373_ clknet_leaf_108_clk _01260_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08065__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ _01437_ _01438_ _05266_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__or4b_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ clknet_leaf_75_clk _00314_ net1251 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07273__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10536_ net1025 _05441_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__nor2_1
XANTENNA__07812__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ clknet_leaf_65_clk _00245_ net1268 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12415__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _05373_ _05379_ _05380_ _05381_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__or4_1
XANTENNA__06637__B_N mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ net296 net2272 net574 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__mux2_1
X_13186_ clknet_leaf_43_clk _00178_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10398_ _05298_ _05318_ _05319_ net1281 screen.counter.ct\[11\] vssd1 vssd1 vccd1
+ vccd1 _05320_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__06640__C _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08773__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _06387_ _06391_ _06394_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__a21oi_1
X_12068_ datapath.mulitply_result\[14\] net325 net321 _06341_ vssd1 vssd1 vccd1 vccd1
+ _00589_ sky130_fd_sc_hd__a22o_1
X_11019_ net190 net2564 net585 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__07879__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06560_ datapath.ru.latched_instruction\[29\] _01487_ _01489_ datapath.ru.latched_instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__o22a_1
XANTENNA__08828__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10096__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06491_ net1278 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08230_ datapath.rf.registers\[31\]\[2\] net989 _01746_ vssd1 vssd1 vccd1 vccd1 _03157_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10618__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08161_ net847 _01667_ _01726_ net982 vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a22o_1
XANTENNA__07199__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08056__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07112_ _02018_ net532 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08092_ net509 _03018_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__or2_1
XANTENNA__07803__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07043_ _01955_ _01956_ _01965_ _01969_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__or4_1
XANTENNA__09005__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12325__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07016__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08359__A3 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09556__A2 _02255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08994_ net502 net618 _03543_ net522 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09308__A2 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _02869_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_149_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A _06452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ datapath.rf.registers\[8\]\[9\] net926 net893 datapath.rf.registers\[14\]\[9\]
+ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a221o_1
X_09615_ _03361_ _03362_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__and2b_2
X_06827_ _01638_ net998 net982 _01682_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__and4_2
XFILLER_0_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ _03871_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__nand2_1
X_06758_ _01419_ net1007 _01655_ _01684_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__a31o_1
X_09477_ net640 _04403_ _04397_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a21boi_1
X_06689_ _01612_ _01613_ _01614_ _01616_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__nand4_1
XFILLER_0_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ _01606_ _01607_ _01618_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_82_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08359_ _01583_ net847 _01651_ _01682_ _01723_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a32o_4
XFILLER_0_74_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14559__1332 vssd1 vssd1 vccd1 vccd1 _14559__1332/HI net1332 sky130_fd_sc_hd__conb_1
XFILLER_0_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07255__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ screen.register.currentYbus\[4\] net133 _05870_ net162 vssd1 vssd1 vccd1
+ vccd1 _00362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ _05035_ _05036_ _05246_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__or3_1
XANTENNA__12235__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07007__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ clknet_leaf_1_clk _00032_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10252_ datapath.PC\[3\] net1309 _05176_ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_
+ sky130_fd_sc_hd__a22oi_4
X_10183_ _04787_ _04804_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nand2_1
Xfanout1203 net1222 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
Xfanout1214 net1216 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_2
Xfanout1225 net1226 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_2
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
Xfanout1247 net1249 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 _05638_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1258 net1261 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1269 net1270 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11375__A _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 _05607_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
X_13942_ clknet_leaf_25_clk _00829_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 _05590_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
X_13873_ clknet_leaf_7_clk _00760_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12824_ net196 net2113 net559 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__mux2_1
X_12755_ net217 net2594 net568 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__mux2_1
XANTENNA__09483__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11706_ _05702_ _05718_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__nand2_1
XANTENNA__07494__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11290__B2 mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12686_ net2035 net226 net433 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06635__C mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14425_ clknet_leaf_61_clk _01312_ net1265 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11637_ screen.counter.currentCt\[0\] _06087_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2_1
XANTENNA__08038__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__A_N _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07246__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ clknet_leaf_115_clk _01243_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11568_ _05303_ _05305_ _05781_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__and3_1
XANTENNA__06932__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13307_ clknet_leaf_110_clk _00297_ net1103 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold708 datapath.rf.registers\[20\]\[14\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10519_ net1050 net1026 _05429_ _01444_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__o31a_1
Xhold719 datapath.rf.registers\[15\]\[31\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10454__A _02234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14287_ clknet_leaf_5_clk _01174_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11499_ _05297_ net1014 _05910_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_123_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13238_ clknet_leaf_78_clk _00228_ net1246 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08746__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ clknet_leaf_27_clk _00161_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_07730_ _02634_ net518 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08297__C _01776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ net652 _02587_ net627 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09400_ _03314_ _04311_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__xnor2_1
X_06612_ _01421_ _01459_ _01503_ _01419_ _01541_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__A _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ net695 _02509_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09331_ net391 _04166_ _04167_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__and3_1
X_06543_ net1306 net1302 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ _01473_ sky130_fd_sc_hd__or3b_2
XANTENNA__06826__B _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _03506_ _04173_ _04181_ _04184_ _04127_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__o311a_1
XANTENNA__07485__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06474_ datapath.ru.latched_instruction\[0\] vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XANTENNA__11281__B2 mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06545__C mmio.memload_or_instruction\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08213_ datapath.rf.registers\[23\]\[2\] net932 net880 datapath.rf.registers\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a22o_1
XANTENNA__08029__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ _03307_ net408 _03458_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout226_A _05502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ datapath.rf.registers\[10\]\[3\] net916 net892 datapath.rf.registers\[14\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a22o_1
XANTENNA__07237__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06842__A _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08985__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ datapath.rf.registers\[4\]\[5\] net809 net725 datapath.rf.registers\[27\]\[5\]
+ _03000_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a221o_1
XANTENNA__10792__A0 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14547__1358 vssd1 vssd1 vccd1 vccd1 net1358 _14547__1358/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout1135_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09529__A2 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07026_ datapath.rf.registers\[31\]\[28\] net818 net731 datapath.rf.registers\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__A0 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08201__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 keypad.debounce.debounce\[13\] vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 datapath.multiplication_module.multiplier_i\[7\] vssd1 vssd1 vccd1 vccd1 net1390
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net636 _03889_ _03899_ net612 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__o2bb2a_1
Xhold35 datapath.multiplication_module.multiplier_i\[15\] vssd1 vssd1 vccd1 vccd1
+ net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 net117 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06763__A2 _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 screen.controlBus\[13\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ datapath.rf.registers\[0\]\[8\] net691 _02841_ _02854_ vssd1 vssd1 vccd1
+ vccd1 _02855_ sky130_fd_sc_hd__o22a_2
Xhold68 screen.controlBus\[14\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 net97 vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ net647 _02783_ _02785_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_67_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ net255 net2115 net598 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _02411_ _02432_ net681 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ net283 net2203 net451 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ net299 net2258 net456 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
XANTENNA__10973__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14210_ clknet_leaf_42_clk _01097_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11422_ net2629 net132 _05896_ net161 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__a22o_1
XANTENNA__07228__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14141_ clknet_leaf_24_clk _01028_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11353_ keypad.apps.button\[0\] keypad.apps.button\[2\] keypad.apps.button\[1\] vssd1
+ vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__or3b_1
XFILLER_0_105_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10304_ net334 _03926_ _05230_ _03532_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a22o_1
XANTENNA__06902__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11089__B _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14072_ clknet_leaf_39_clk _00959_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11284_ net4 net1045 net1034 mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1
+ vccd1 _00298_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ clknet_leaf_37_clk _00015_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ _05094_ _05161_ _04447_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a21bo_1
Xfanout1000 _01641_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_1
Xfanout1011 _05308_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_4
Xfanout1022 _05697_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_4
XANTENNA__07400__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1033 net1034 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_2
X_10166_ _04811_ _04809_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__and2b_1
XANTENNA__09940__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 net1045 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_2
XANTENNA__11309__S _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_2
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
Xfanout1077 net1078 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_4
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
X_10097_ _01433_ _03585_ net1274 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a21bo_1
Xfanout1099 net1102 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
X_13925_ clknet_leaf_93_clk _00812_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13856_ clknet_leaf_46_clk _00743_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12807_ net276 net1905 net559 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__mux2_1
XANTENNA__13474__RESET_B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__A _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08259__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09456__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13787_ clknet_leaf_52_clk _00674_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10999_ net277 net1924 net582 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__C net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ net286 net2039 net566 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__mux2_1
XANTENNA__07467__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11263__B2 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10883__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ net2354 net299 net432 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14408_ clknet_leaf_11_clk _01295_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ clknet_leaf_105_clk _01226_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold505 datapath.rf.registers\[6\]\[25\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 datapath.rf.registers\[11\]\[7\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 datapath.rf.registers\[10\]\[28\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 datapath.rf.registers\[5\]\[17\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06812__D _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold549 datapath.rf.registers\[12\]\[13\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08900_ net634 _03810_ _03823_ net610 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06993__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12603__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _04754_ _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08831_ net500 net620 net488 net526 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__o211a_1
Xhold1205 datapath.rf.registers\[19\]\[21\] vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 mmio.memload_or_instruction\[4\] vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 mmio.memload_or_instruction\[16\] vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ _02079_ net532 net353 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__mux2_1
Xhold1238 datapath.rf.registers\[19\]\[15\] vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 screen.register.currentXbus\[7\] vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
X_14558__1331 vssd1 vssd1 vccd1 vccd1 _14558__1331/HI net1331 sky130_fd_sc_hd__conb_1
X_07713_ datapath.rf.registers\[3\]\[13\] net964 net848 datapath.rf.registers\[1\]\[13\]
+ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a221o_1
X_08693_ _03608_ _03610_ _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07644_ datapath.rf.registers\[31\]\[14\] net817 net765 datapath.rf.registers\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07170__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07575_ datapath.rf.registers\[21\]\[16\] net939 net934 datapath.rf.registers\[23\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1085_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09314_ net369 _04131_ _04240_ net382 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a211o_1
X_06526_ mmio.key_data\[3\] mmio.memload_or_instruction\[3\] net1060 vssd1 vssd1 vccd1
+ vccd1 _01456_ sky130_fd_sc_hd__mux2_2
XANTENNA__11254__B2 _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09245_ net397 _04171_ _04168_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_32_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout510_A _02951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ net401 _03897_ _04102_ net336 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o211a_1
XANTENNA__08958__A0 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ datapath.rf.registers\[23\]\[4\] net788 net763 datapath.rf.registers\[17\]\[4\]
+ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08058_ datapath.rf.registers\[30\]\[5\] net908 net896 datapath.rf.registers\[6\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a22o_1
XANTENNA__07630__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout977_A _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
X_07009_ datapath.rf.registers\[25\]\[29\] net874 net863 datapath.rf.registers\[28\]\[29\]
+ _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a221o_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__12513__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
X_10020_ net1052 _03584_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__or2_1
XANTENNA__07394__C1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ net212 net1628 net581 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__mux2_1
XANTENNA__10968__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ clknet_leaf_57_clk datapath.multiplication_module.multiplicand_i_n\[27\]
+ net1257 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net164 net2182 net596 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__mux2_1
XANTENNA__07697__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07161__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ clknet_leaf_70_clk _00579_ net1228 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10853_ net2073 net163 net603 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13572_ clknet_leaf_88_clk _00522_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11245__B2 _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10784_ net1277 _05485_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11796__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ net1773 net223 net454 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12454_ net243 net2050 net461 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11548__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ _02234_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ net248 net2433 net469 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XANTENNA__10756__B1 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14124_ clknet_leaf_32_clk _01011_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11336_ _01461_ net1028 net307 net311 datapath.ru.latched_instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__a32o_1
XANTENNA__07621__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14055_ clknet_leaf_20_clk _00942_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12423__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ net1308 net143 net137 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__a21o_1
X_13006_ net2292 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__clkbuf_1
X_10218_ datapath.PC\[15\] net1251 _05143_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_
+ sky130_fd_sc_hd__o22a_1
X_11198_ _01404_ _05256_ _05838_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10149_ _04792_ _04794_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_128_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10878__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09677__B2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ clknet_leaf_117_clk _00795_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546__1357 vssd1 vssd1 vccd1 vccd1 net1357 _14546__1357/LO sky130_fd_sc_hd__conb_1
XANTENNA__07152__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ clknet_leaf_6_clk _00726_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06807__D net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07360_ datapath.rf.registers\[19\]\[21\] net945 net878 datapath.rf.registers\[29\]\[21\]
+ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a221o_1
XANTENNA__11236__B2 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07291_ datapath.rf.registers\[11\]\[22\] net776 net757 datapath.rf.registers\[24\]\[22\]
+ _02216_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ net335 _03528_ _03956_ net640 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__o211a_1
XANTENNA__06663__A1 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09062__C1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 datapath.rf.registers\[21\]\[16\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 datapath.rf.registers\[12\]\[12\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 datapath.rf.registers\[21\]\[12\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold335 net67 vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 datapath.rf.registers\[12\]\[19\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 datapath.rf.registers\[29\]\[23\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 datapath.rf.registers\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _04850_ _04851_ _04852_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold379 datapath.rf.registers\[20\]\[0\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12333__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout804 _01751_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_8
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_4
Xfanout826 _01740_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_4
X_09863_ _04788_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__nor2_1
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_2
Xfanout848 net851 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout293_A _05590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _01853_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
Xhold1002 datapath.mulitply_result\[29\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ _03339_ _03704_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__a21oi_1
Xhold1013 datapath.rf.registers\[11\]\[23\] vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _01426_ _02906_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__nand2_1
Xhold1024 datapath.rf.registers\[23\]\[19\] vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 datapath.rf.registers\[2\]\[26\] vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__B1 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07391__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 datapath.rf.registers\[16\]\[14\] vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1057 datapath.rf.registers\[13\]\[11\] vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net502 net618 _03543_ _01950_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout460_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 datapath.rf.registers\[4\]\[9\] vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10788__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 datapath.rf.registers\[16\]\[29\] vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _03601_ _03602_ net414 vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__mux2_1
XANTENNA__08876__C1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ datapath.rf.registers\[21\]\[15\] net938 net901 datapath.rf.registers\[20\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07558_ datapath.rf.registers\[15\]\[16\] net807 net736 datapath.rf.registers\[12\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06509_ screen.controlBus\[1\] vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07489_ datapath.rf.registers\[3\]\[18\] net965 net886 datapath.rf.registers\[9\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a22o_1
X_09228_ net380 _04154_ _04148_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07851__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09159_ net688 _04083_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a21o_1
X_12170_ _01446_ _01449_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__nand2_1
XANTENNA__07603__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _05705_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12243__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold880 datapath.rf.registers\[31\]\[31\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 datapath.rf.registers\[20\]\[30\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11367__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ net1300 net1301 vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09118__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08022__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ net208 _04929_ net1312 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a21oi_1
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__A _02721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ net279 net1665 net578 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__mux2_1
XANTENNA__07134__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ net249 net2337 net594 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11885_ net158 _05870_ net150 screen.controlBus\[4\] vssd1 vssd1 vccd1 vccd1 _00483_
+ sky130_fd_sc_hd__a22o_1
X_13624_ clknet_leaf_29_clk _00562_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ _03909_ _05662_ net844 vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__mux2_1
XANTENNA__11769__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13555_ clknet_leaf_88_clk _00505_ net1219 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08095__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12418__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ net840 _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12506_ net1570 net295 net453 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__mux2_1
XANTENNA__07842__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ clknet_leaf_82_clk _00439_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ datapath.mulitply_result\[27\] net427 net660 vssd1 vssd1 vccd1 vccd1 _05547_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10446__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14557__1330 vssd1 vssd1 vccd1 vccd1 _14557__1330/HI net1330 sky130_fd_sc_hd__conb_1
XFILLER_0_63_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12437_ net289 net2414 net460 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XANTENNA__10729__B1 _05572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ net1799 net163 net473 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__mux2_1
X_14107_ clknet_leaf_19_clk _00994_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11319_ datapath.ru.ack_mul_reg _05852_ _05853_ _05858_ _05857_ vssd1 vssd1 vccd1
+ vccd1 _05859_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10462__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net1662 net169 net482 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__mux2_1
X_14038_ clknet_leaf_25_clk _00925_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_06860_ datapath.rf.registers\[13\]\[31\] net793 net749 datapath.rf.registers\[10\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06791_ _01584_ _01593_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08530_ net977 _03446_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__nand2_1
XANTENNA__08322__A1 _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07125__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08322__B2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08461_ _03181_ _03387_ _03180_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07412_ datapath.rf.registers\[19\]\[20\] net946 net879 datapath.rf.registers\[29\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08392_ _02885_ _03318_ _02880_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a21oi_1
X_07343_ datapath.rf.registers\[10\]\[21\] net749 net731 datapath.rf.registers\[16\]\[21\]
+ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12328__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout139_A _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ datapath.rf.registers\[27\]\[23\] net870 net853 datapath.rf.registers\[5\]\[23\]
+ _02200_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09013_ net418 _03646_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_154_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold110 net66 vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold121 datapath.PC\[12\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 net74 vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold143 datapath.multiplication_module.multiplicand_i\[30\] vssd1 vssd1 vccd1 vccd1
+ net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 net57 vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 mmio.memload_or_instruction\[3\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold176 datapath.rf.registers\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 datapath.rf.registers\[31\]\[2\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _05668_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_4
Xhold198 datapath.multiplication_module.multiplicand_i\[26\] vssd1 vssd1 vccd1 vccd1
+ net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _03561_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11187__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09915_ datapath.PC\[28\] net628 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nand2_1
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_4
Xfanout634 _03560_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout656 _01622_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
Xfanout667 _06088_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08010__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _04674_ _04772_ _04671_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a21oi_2
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07364__A2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 _03355_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08561__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__inv_2
X_06989_ datapath.rf.registers\[11\]\[29\] net776 net750 datapath.rf.registers\[10\]\[29\]
+ _01911_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a221o_1
X_08728_ _03653_ _03654_ net408 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07116__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08659_ datapath.PC\[23\] net1274 _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11670_ screen.counter.currentCt\[11\] _06120_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__and2_1
X_10621_ _01643_ _01667_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__nand2_2
XFILLER_0_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08077__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12238__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ clknet_leaf_97_clk _00325_ net1218 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07824__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ _05432_ _05459_ _05460_ _05455_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13271_ clknet_leaf_90_clk _00261_ net1209 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10981__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10483_ _05389_ _05391_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_20_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12222_ net232 net2527 net576 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__mux2_1
XANTENNA__10187__A1 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545__1356 vssd1 vssd1 vccd1 vccd1 net1356 _14545__1356/LO sky130_fd_sc_hd__conb_1
X_12153_ net2469 net327 net323 _06412_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a22o_1
XANTENNA__10282__A _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11104_ screen.counter.ct\[13\] _01439_ net1288 screen.counter.ct\[15\] vssd1 vssd1
+ vccd1 vccd1 _05754_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_9_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12084_ _06352_ _06353_ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__or3_1
X_11035_ net1279 _05323_ _05685_ _05300_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a31o_1
XANTENNA__12701__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10221__S net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ net2417 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07107__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11937_ net153 _05889_ net128 net2636 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11868_ datapath.PC\[30\] net305 _06254_ _06256_ vssd1 vssd1 vccd1 vccd1 _00474_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13607_ clknet_leaf_107_clk _00545_ net1110 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08068__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ datapath.mulitply_result\[14\] net428 _05645_ _05648_ net659 vssd1 vssd1
+ vccd1 vccd1 _05649_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11799_ net833 _04081_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ clknet_leaf_87_clk _00488_ net1219 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13469_ clknet_leaf_80_clk net1384 net1239 vssd1 vssd1 vccd1 vccd1 screen.counter.ack3
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10891__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06670__A _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10178__A1 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08240__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ datapath.rf.registers\[3\]\[7\] net964 net936 datapath.rf.registers\[21\]\[7\]
+ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__a221o_1
X_09700_ net678 _04626_ _03440_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__mux2_1
X_06912_ net1001 net985 net980 _01812_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__and4_1
XANTENNA__12611__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ datapath.rf.registers\[19\]\[9\] net760 net727 datapath.rf.registers\[2\]\[9\]
+ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a221o_1
XANTENNA__07346__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ net674 _04544_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06843_ net990 _01731_ _01742_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__and3_1
XANTENNA__06829__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ net656 _04485_ _04487_ _04488_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__and4_1
X_06774_ datapath.ru.latched_instruction\[9\] _01643_ _01666_ datapath.ru.latched_instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08513_ _01864_ _03439_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__xor2_2
XFILLER_0_148_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09493_ _04007_ _04046_ _04386_ _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout256_A _05644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ _02370_ net523 vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08059__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ datapath.rf.registers\[8\]\[0\] net925 net883 datapath.rf.registers\[17\]\[0\]
+ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07326_ datapath.rf.registers\[10\]\[22\] net918 net887 datapath.rf.registers\[9\]\[22\]
+ _02252_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a221o_1
XANTENNA__07806__B1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09271__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07257_ datapath.rf.registers\[14\]\[23\] net800 net735 datapath.rf.registers\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07188_ datapath.rf.registers\[22\]\[25\] net954 net890 datapath.rf.registers\[12\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
XANTENNA__11366__B1 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07585__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout431 net435 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_4
XANTENNA__10830__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12521__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout464 net467 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07337__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 _06453_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08534__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout486 net487 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_4
X_09829_ _04708_ _04712_ _04755_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__and3_1
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
X_12840_ net275 net2151 net555 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ net286 net1902 net561 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10976__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ clknet_leaf_2_clk _01397_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11722_ screen.counter.ct\[7\] net665 _06154_ net712 vssd1 vssd1 vccd1 vccd1 _00430_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10644__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ screen.counter.currentCt\[5\] _06108_ net666 vssd1 vssd1 vccd1 vccd1 _06111_
+ sky130_fd_sc_hd__o21ai_1
X_14441_ clknet_leaf_13_clk _01328_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10604_ net1551 net346 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[16\]
+ sky130_fd_sc_hd__and2_1
X_14372_ clknet_leaf_104_clk _01259_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11584_ net1290 net1291 screen.counter.ct\[17\] net1285 vssd1 vssd1 vccd1 vccd1 _06048_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_92_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13323_ clknet_leaf_76_clk _00313_ net1248 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_10535_ _05401_ _05406_ _05440_ _05444_ _05404_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a311o_1
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13254_ clknet_leaf_65_clk _00244_ net1268 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
X_10466_ net507 _03087_ _03146_ _03207_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__or4_1
XANTENNA__09014__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ net291 net2271 net574 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
X_13185_ clknet_leaf_42_clk _00177_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10397_ net1301 screen.counter.ct\[3\] net1293 screen.counter.ct\[22\] vssd1 vssd1
+ vccd1 vccd1 _05319_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07576__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12136_ datapath.mulitply_result\[26\] datapath.multiplication_module.multiplicand_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__or2_1
XANTENNA__10580__A1 _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12431__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ _06337_ _06339_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07328__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net192 net2443 net584 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10886__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ net282 net2249 net606 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06490_ datapath.rf.registers\[0\]\[8\] vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
XANTENNA__07500__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09238__C1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ datapath.rf.registers\[0\]\[3\] net690 _03075_ _03086_ vssd1 vssd1 vccd1
+ vccd1 _03087_ sky130_fd_sc_hd__o22a_4
XANTENNA__11045__C1 _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07111_ datapath.rf.registers\[0\]\[27\] net693 _02025_ _02037_ vssd1 vssd1 vccd1
+ vccd1 _02038_ sky130_fd_sc_hd__o22a_2
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _02998_ _03017_ net650 vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_151_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12606__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07042_ datapath.rf.registers\[8\]\[28\] net738 _01966_ _01968_ net832 vssd1 vssd1
+ vccd1 vccd1 _01969_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_141_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06831__C _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07567__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ _02432_ _03545_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nand2_1
XANTENNA__06775__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07944_ datapath.rf.registers\[3\]\[8\] net766 net743 datapath.rf.registers\[1\]\[8\]
+ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a221o_1
XANTENNA__12341__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07319__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ datapath.rf.registers\[21\]\[9\] net938 net853 datapath.rf.registers\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a22o_1
X_06826_ net993 _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__and2_2
X_09614_ _04499_ _04518_ _04540_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor3b_1
X_09545_ _03909_ _04449_ _04471_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__and3_1
X_06757_ _01418_ net1006 _01637_ _01642_ _01412_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a32o_1
XFILLER_0_149_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11823__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ net339 _04399_ _04402_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a21o_1
XANTENNA__06575__A mmio.memload_or_instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14544__1355 vssd1 vssd1 vccd1 vccd1 net1355 _14544__1355/LO sky130_fd_sc_hd__conb_1
X_06688_ datapath.ru.latched_instruction\[29\] net1041 net1008 _01615_ vssd1 vssd1
+ vccd1 vccd1 _01616_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_22_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ _01608_ _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout805_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ datapath.rf.registers\[0\]\[0\] net830 _03279_ _03284_ vssd1 vssd1 vccd1
+ vccd1 _03285_ sky130_fd_sc_hd__o22a_4
XFILLER_0_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07309_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08289_ datapath.rf.registers\[29\]\[1\] net990 _01756_ vssd1 vssd1 vccd1 vccd1 _03216_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12516__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10320_ _05037_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08204__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ net200 _04790_ _05177_ net1243 vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__o31a_1
XANTENNA__07558__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _04417_ _05104_ _05108_ net204 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__a211oi_1
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__clkbuf_4
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_4
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_2
Xfanout1237 net1242 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_2
XANTENNA__12251__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 _05650_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_1
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 net264 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
Xfanout1259 net1261 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout272 _05622_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
Xfanout283 _05602_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
X_13941_ clknet_leaf_29_clk _00828_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10314__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout294 _05596_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
X_13872_ clknet_leaf_4_clk _00759_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07191__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12823_ net212 net2276 net559 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__mux2_1
XANTENNA__11391__A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12754_ net224 net2263 net567 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11705_ net712 net663 net1301 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__mux2_1
X_12685_ net1735 net243 net433 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11636_ screen.counter.currentEnable _06081_ net713 vssd1 vssd1 vccd1 vccd1 _06099_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA__06635__D mmio.memload_or_instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14424_ clknet_leaf_39_clk _01311_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11567_ net1013 _05740_ _05742_ _05747_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__or4_1
XANTENNA__12426__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14355_ clknet_leaf_60_clk _01242_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07797__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13306_ clknet_leaf_112_clk _00296_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_10518_ _05409_ _05422_ net1025 vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__o21ba_1
X_14286_ clknet_leaf_116_clk _01173_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 datapath.rf.registers\[6\]\[12\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11498_ _05305_ _05782_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__nor2_1
XANTENNA__10454__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ clknet_leaf_78_clk _00227_ net1246 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
X_10449_ _02971_ _03017_ _03060_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__or3_1
XANTENNA__07549__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13168_ clknet_leaf_4_clk _00160_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _06382_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__or2_1
X_13099_ clknet_leaf_55_clk _00091_ net1175 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09171__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07660_ datapath.rf.registers\[0\]\[14\] _02586_ net827 vssd1 vssd1 vccd1 vccd1 _02587_
+ sky130_fd_sc_hd__mux2_4
XANTENNA__07182__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07721__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ datapath.ru.latched_instruction\[23\] _01502_ _01513_ datapath.ru.latched_instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07591_ _02511_ _02513_ _02515_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__or4_1
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ net395 _04176_ _04254_ net403 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a211o_1
X_06542_ mmio.memload_or_instruction\[8\] net1062 vssd1 vssd1 vccd1 vccd1 _01472_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08131__C1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ _04157_ _04187_ net615 _04127_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__o211a_1
X_06473_ datapath.ru.zero_multi1 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
X_08212_ datapath.rf.registers\[30\]\[2\] net909 net857 datapath.rf.registers\[15\]\[2\]
+ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a221o_1
X_09192_ _03641_ _03643_ net408 vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08143_ datapath.rf.registers\[2\]\[3\] net923 net861 datapath.rf.registers\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06842__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_A _05519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__A1 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ datapath.rf.registers\[15\]\[5\] net805 net744 datapath.rf.registers\[21\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a22o_1
XANTENNA__06996__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07025_ _01930_ net534 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout588_A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 keypad.debounce.debounce\[3\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _03330_ _03873_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21a_1
Xhold25 keypad.debounce.debounce\[12\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 datapath.multiplication_module.multiplier_i\[13\] vssd1 vssd1 vccd1 vccd1
+ net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 net118 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ _02849_ _02851_ _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or3_1
Xhold58 net64 vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 screen.controlBus\[21\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ net650 _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__or2_1
XANTENNA__07173__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07712__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ _01731_ net973 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__and2_2
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07789_ datapath.rf.registers\[31\]\[11\] net817 net809 datapath.rf.registers\[4\]\[11\]
+ _02703_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ net415 _04392_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09459_ _04116_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12470_ net287 net1522 net456 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11421_ net344 net714 vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12246__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ clknet_leaf_57_clk _01027_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11352_ _01488_ net1030 net310 net314 datapath.ru.latched_instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06987__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ _03552_ net612 vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14071_ clknet_leaf_44_clk _00958_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11283_ net3 net1046 net1035 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1
+ vccd1 _00297_ sky130_fd_sc_hd__a22o_1
X_13022_ clknet_leaf_50_clk _00014_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10234_ net701 _04446_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__nand2_1
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_2
Xfanout1012 _05308_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
X_10165_ datapath.PC\[11\] net1248 _05090_ _05091_ vssd1 vssd1 vccd1 vccd1 _05092_
+ sky130_fd_sc_hd__o22a_1
Xfanout1023 _05697_ vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1034 _05848_ vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_4
Xfanout1045 _05846_ vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_4
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__clkbuf_4
Xfanout1067 net1070 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
X_10096_ net538 _03703_ _05022_ net1057 vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__a211o_1
Xfanout1078 net1085 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
Xfanout1089 net1125 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09153__B2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ clknet_leaf_15_clk _00811_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07164__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13855_ clknet_leaf_38_clk _00742_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12806_ net278 net1851 net557 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10998_ net281 net2208 net582 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__mux2_1
X_13786_ clknet_leaf_22_clk _00673_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10449__B _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12737_ net295 net1642 net567 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ net1856 net289 net432 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XANTENNA__09208__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14407_ clknet_leaf_16_clk _01294_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11619_ _05756_ _06069_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__nand2_1
XANTENNA__10465__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ net2540 net164 net445 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
XANTENNA__08967__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14338_ clknet_leaf_33_clk _01225_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold506 datapath.rf.registers\[13\]\[13\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 datapath.rf.registers\[18\]\[19\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 datapath.rf.registers\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 datapath.rf.registers\[19\]\[8\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14269_ clknet_leaf_33_clk _01156_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14543__1354 vssd1 vssd1 vccd1 vccd1 net1354 _14543__1354/LO sky130_fd_sc_hd__conb_1
X_08830_ _03755_ _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1206 datapath.rf.registers\[24\]\[0\] vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 datapath.rf.registers\[23\]\[22\] vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ _03686_ _03687_ net388 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
Xhold1228 datapath.rf.registers\[17\]\[22\] vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 screen.controlBus\[5\] vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
X_07712_ datapath.rf.registers\[17\]\[13\] net880 net856 datapath.rf.registers\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a22o_1
X_08692_ net421 _03614_ _03618_ net317 vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a211o_1
X_07643_ datapath.rf.registers\[23\]\[14\] net786 net744 datapath.rf.registers\[21\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__B _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07574_ _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__inv_2
XANTENNA__09447__A2 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ _04140_ _04143_ _03538_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__o21a_1
X_06525_ net1306 net1302 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__nor2_2
XANTENNA__11254__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_62_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09244_ net390 _04015_ _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07949__A _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ net401 _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout503_A _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ datapath.rf.registers\[7\]\[4\] net825 net797 datapath.rf.registers\[25\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a22o_1
XANTENNA__08958__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ datapath.rf.registers\[31\]\[5\] net948 net904 datapath.rf.registers\[24\]\[5\]
+ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07008_ datapath.rf.registers\[3\]\[29\] net966 net942 datapath.rf.registers\[26\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a22o_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XANTENNA_fanout872_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__08186__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07933__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _03847_ _03885_ net367 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__mux2_1
X_11970_ net216 net2439 net581 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XANTENNA__07146__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ net168 net2121 net596 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13640_ clknet_leaf_70_clk _00578_ net1229 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10852_ net1589 net170 net604 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11245__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ clknet_leaf_89_clk _00521_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10783_ net2007 net274 net604 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__mux2_1
XANTENNA__10984__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
X_12522_ net2016 net233 net453 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12453_ net236 net1811 net460 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11404_ screen.register.currentYbus\[21\] net133 _05887_ net162 vssd1 vssd1 vccd1
+ vccd1 _00379_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12384_ net251 net1859 net468 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XANTENNA__09071__B1 _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10756__B2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11335_ mmio.memload_or_instruction\[14\] net1063 net309 net313 datapath.ru.latched_instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__a32o_1
X_14123_ clknet_leaf_56_clk _01010_ net1257 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09793__B _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12704__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14054_ clknet_leaf_111_clk _00941_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11266_ net1445 net140 net134 _01799_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__a22o_1
X_10217_ net205 _05136_ net1311 vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a21o_1
X_13005_ net1481 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__clkbuf_1
X_11197_ _01404_ _05256_ _05838_ _05253_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a22o_1
XANTENNA__07385__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10451__C _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net698 _04337_ _05070_ _05074_ net203 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_128_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11844__A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ _04833_ _04835_ _04778_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07137__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ clknet_leaf_59_clk _00794_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13838_ clknet_leaf_2_clk _00725_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10894__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08637__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ clknet_leaf_3_clk _00656_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08101__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07290_ datapath.rf.registers\[9\]\[22\] net780 net736 datapath.rf.registers\[12\]\[22\]
+ _02215_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06663__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11944__B1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 datapath.rf.registers\[3\]\[24\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold314 datapath.rf.registers\[27\]\[7\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 datapath.rf.registers\[17\]\[25\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12614__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 datapath.rf.registers\[31\]\[5\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 datapath.rf.registers\[18\]\[25\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 datapath.rf.registers\[15\]\[16\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 datapath.rf.registers\[15\]\[18\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _04856_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__nand2_1
Xfanout805 net808 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
Xfanout816 _01748_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09862_ _04732_ _04740_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__xnor2_1
Xfanout827 net830 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_6
Xfanout838 _01722_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_2
Xfanout849 net851 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_4
XANTENNA__07915__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1003 datapath.rf.registers\[25\]\[10\] vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net706 _03739_ net491 vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__o21a_1
Xhold1014 columns.count\[2\] vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _01426_ _02906_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nor2_1
Xhold1025 screen.counter.currentCt\[4\] vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout286_A _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1036 datapath.rf.registers\[20\]\[25\] vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 datapath.rf.registers\[6\]\[8\] vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 datapath.rf.registers\[26\]\[11\] vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _01905_ net359 vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__nand2_1
XANTENNA__07128__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 datapath.rf.registers\[20\]\[29\] vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06848__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _03464_ _03467_ net408 vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout453_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1195_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ datapath.rf.registers\[30\]\[15\] net910 _02548_ _02550_ _02552_ vssd1 vssd1
+ vccd1 vccd1 _02553_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_138_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07557_ datapath.rf.registers\[30\]\[16\] net772 net761 datapath.rf.registers\[19\]\[16\]
+ _02482_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
X_06508_ screen.controlBus\[0\] vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07488_ datapath.rf.registers\[20\]\[18\] net901 net897 datapath.rf.registers\[6\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07300__B1 _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09227_ net372 _04150_ _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09158_ net708 _04084_ net624 vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_79_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11935__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08109_ datapath.rf.registers\[8\]\[4\] net926 net853 datapath.rf.registers\[5\]\[4\]
+ _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12524__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _02566_ net356 _04013_ _03522_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__a211o_1
X_11120_ _05753_ _05754_ _05755_ _05757_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__or4_2
Xhold870 datapath.rf.registers\[8\]\[23\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold881 datapath.rf.registers\[31\]\[30\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 datapath.rf.registers\[9\]\[2\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ screen.counter.ct\[3\] net1298 vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__nand2_1
XANTENNA__07367__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _04782_ _04829_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10979__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11383__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ net280 net2060 net578 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__mux2_1
X_10904_ net253 net2092 net594 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ net157 _05869_ net150 net2078 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a22o_1
XANTENNA__08973__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13623_ clknet_leaf_28_clk _00561_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10835_ _05491_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
X_14542__1353 vssd1 vssd1 vccd1 vccd1 net1353 _14542__1353/LO sky130_fd_sc_hd__conb_1
X_13554_ clknet_leaf_88_clk _00504_ net1219 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10766_ _01425_ _05483_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12505_ net1577 net291 net455 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__mux2_1
X_13485_ clknet_leaf_82_clk _00438_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10219__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697_ _04561_ _05545_ net845 vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__mux2_1
X_12436_ net181 net2642 net463 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
XANTENNA__10729__A1 _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11926__B1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12434__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net1805 net167 net474 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14106_ clknet_leaf_23_clk _00993_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11318_ datapath.ru.ack_mul_reg2 net1029 _01601_ datapath.ru.ack_mul_reg vssd1 vssd1
+ vccd1 vccd1 _05858_ sky130_fd_sc_hd__or4b_1
XANTENNA__07070__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12298_ net1708 net172 net483 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__mux2_1
XANTENNA__10462__B _02476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11249_ net1474 net141 net136 _02587_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__a22o_1
XANTENNA__09347__B2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ clknet_leaf_29_clk _00924_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07358__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06790_ _01606_ _01607_ _01618_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__or3_4
XANTENNA__09044__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ _03251_ _03288_ _03308_ _03250_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07411_ datapath.rf.registers\[20\]\[20\] net902 net898 datapath.rf.registers\[6\]\[20\]
+ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08391_ _02932_ _03317_ _02928_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12609__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
X_07342_ datapath.rf.registers\[23\]\[21\] net787 net723 datapath.rf.registers\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06834__C _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07273_ datapath.rf.registers\[22\]\[23\] net953 net949 datapath.rf.registers\[31\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a22o_1
X_09012_ net422 _03659_ net318 vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_154_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 datapath.rf.registers\[0\]\[29\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold111 screen.controlBus\[17\] vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12344__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout201_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 net95 vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 screen.counter.currentEnable vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06850__B _01776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 net100 vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__C1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07061__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 datapath.multiplication_module.multiplicand_i\[24\] vssd1 vssd1 vccd1 vccd1
+ net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 datapath.rf.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 net119 vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 datapath.multiplication_module.multiplicand_i\[27\] vssd1 vssd1 vccd1 vccd1
+ net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 datapath.rf.registers\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net605 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_8
X_09914_ _04837_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__nand2_1
Xfanout613 _03554_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07349__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 _03357_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1208_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net647 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _04771_ _04770_ _04769_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__or3b_1
Xfanout657 _01622_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_2
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10799__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 _03500_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_4
X_09776_ net632 _04701_ datapath.PC\[13\] vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__o21a_1
X_06988_ datapath.rf.registers\[3\]\[29\] net767 net761 datapath.rf.registers\[19\]\[29\]
+ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a221o_1
X_08727_ net519 net518 net404 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout835_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08658_ _01432_ _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_105_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ datapath.rf.registers\[20\]\[15\] net802 net727 datapath.rf.registers\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XANTENNA__12519__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ _03512_ net398 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__nand2_2
XFILLER_0_138_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10620_ _01650_ _01668_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__nand2_2
XFILLER_0_107_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12181__A_N _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10551_ _05405_ _05406_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _05390_ _05392_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__or3_1
X_13270_ clknet_leaf_92_clk _00260_ net1202 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09577__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ net229 net2142 net575 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__mux2_1
XANTENNA__12254__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _06409_ _06410_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__xor2_1
XANTENNA__07052__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ net1295 net1281 net1282 screen.counter.ct\[4\] vssd1 vssd1 vccd1 vccd1 _05753_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_130_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12083_ datapath.mulitply_result\[17\] datapath.multiplication_module.multiplicand_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11034_ net1290 net1288 net1283 vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__and3_1
XANTENNA__08001__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08050__A_N net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12985_ net1516 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
X_11936_ net153 _05888_ net128 net2640 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07512__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06866__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ _05566_ net176 _06255_ net179 vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a22o_1
XANTENNA__12429__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06935__B _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ clknet_leaf_14_clk _00544_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_151_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10818_ net841 _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ net200 _04807_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ clknet_leaf_88_clk _00487_ net1217 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06618__A2 _01473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10749_ _01456_ net709 _05589_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__o21a_2
XFILLER_0_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13468_ clknet_leaf_80_clk net1371 net1239 vssd1 vssd1 vccd1 vccd1 screen.counter.ack2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07291__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12419_ net2077 net240 net466 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
X_13399_ clknet_leaf_77_clk _00000_ net1246 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07579__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ datapath.rf.registers\[7\]\[7\] net956 net912 datapath.rf.registers\[18\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_4_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_06911_ net1001 net985 net978 _01812_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__and4_1
X_07891_ datapath.rf.registers\[18\]\[9\] net790 net763 datapath.rf.registers\[17\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09630_ net615 _04552_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__and3_1
X_06842_ _01738_ net972 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06829__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ datapath.ru.latched_instruction\[11\] _01664_ _01698_ _01699_ vssd1 vssd1
+ vccd1 vccd1 _01700_ sky130_fd_sc_hd__a211o_1
X_09561_ net338 _04180_ net315 vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10638__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ _01908_ _03435_ _03436_ _01907_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__o31a_1
X_09492_ _04081_ _04416_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08700__C1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ _02281_ _02301_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nor2_1
XANTENNA__06857__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12339__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06845__B _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ datapath.rf.registers\[28\]\[0\] net861 net851 datapath.rf.registers\[1\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07022__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07325_ datapath.rf.registers\[18\]\[22\] net915 net874 datapath.rf.registers\[25\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1060_A _01455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1158_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ _02179_ _02181_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_59_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07282__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07187_ datapath.rf.registers\[24\]\[25\] net906 net894 datapath.rf.registers\[14\]\[25\]
+ _02113_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07034__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout785_A _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 _03455_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07990__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_2
XFILLER_0_10_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 _06463_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 _06461_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_4
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout952_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net467 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_8
Xfanout476 _06452_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_8
X_09828_ _04714_ _04717_ _04752_ _04713_ _04711_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a311o_1
Xfanout487 _06447_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout498 _03542_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
X_09759_ _01676_ _04678_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ net294 net1656 net562 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _06069_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__nor2_1
XANTENNA__12249__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ clknet_leaf_13_clk _01327_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11652_ screen.counter.currentCt\[5\] _06108_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ net1528 net520 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[15\]
+ sky130_fd_sc_hd__mux2_1
X_14371_ clknet_leaf_105_clk _01258_ net1101 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10992__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11583_ net1279 screen.counter.ct\[22\] _05705_ net1280 vssd1 vssd1 vccd1 vccd1 _06047_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10801__B1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ clknet_leaf_75_clk _00312_ net1250 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_10534_ net1048 _05442_ _05443_ _05434_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a22o_1
XANTENNA__07273__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11389__A _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13253_ clknet_leaf_76_clk _00243_ net1248 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
X_10465_ net533 net532 _02997_ _03307_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__or4_1
X_12204_ net300 net1894 net573 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
X_10396_ screen.counter.ct\[6\] screen.counter.ct\[12\] net1284 net1280 vssd1 vssd1
+ vccd1 vccd1 _05318_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ clknet_leaf_48_clk _00176_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12135_ datapath.mulitply_result\[26\] datapath.multiplication_module.multiplicand_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_131_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12712__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__A _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ _06337_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nand2b_1
X_11017_ net199 net1972 net585 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
XANTENNA__12013__A datapath.mulitply_result\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ net285 net2097 net606 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__mux2_1
XANTENNA__10096__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net153 _05871_ net128 net2149 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__a22o_1
XANTENNA__11293__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12899_ net2033 net287 net548 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14569_ net1339 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ net695 _02027_ _02036_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__or3_1
X_08090_ datapath.rf.registers\[0\]\[5\] net827 _03009_ _03016_ vssd1 vssd1 vccd1
+ vccd1 _03017_ sky130_fd_sc_hd__o22a_4
XANTENNA__06681__A _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07041_ datapath.rf.registers\[6\]\[28\] net814 net735 datapath.rf.registers\[12\]\[28\]
+ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11348__A1 _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07016__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12622__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ net523 net359 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__or2_1
XANTENNA__06775__B2 datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07943_ datapath.rf.registers\[14\]\[8\] net799 net774 datapath.rf.registers\[11\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a22o_1
XANTENNA__06551__C_N mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout199_A _05537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06527__A1 mmio.memload_or_instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ datapath.rf.registers\[3\]\[9\] net965 net849 datapath.rf.registers\[1\]\[9\]
+ _02800_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a221o_1
XANTENNA__07724__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ _04535_ _04539_ _03558_ _04521_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__o2bb2a_1
X_06825_ _01639_ _01646_ net982 net977 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__and4_2
XFILLER_0_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout366_A _03540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ net673 _04450_ _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o21a_1
X_06756_ _01409_ _01597_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10087__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11284__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06687_ mmio.memload_or_instruction\[29\] net1063 net1029 vssd1 vssd1 vccd1 vccd1
+ _01615_ sky130_fd_sc_hd__and3_1
X_09475_ net335 _04400_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout533_A _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08426_ _01606_ _01618_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout700_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ _03280_ _03281_ _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07308_ net649 _02234_ net626 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07255__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08288_ datapath.rf.registers\[21\]\[1\] net745 _03212_ _03213_ _03214_ vssd1 vssd1
+ vccd1 vccd1 _03215_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07239_ _02161_ _02163_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__or3_1
XANTENNA__11339__B2 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ _04788_ _04789_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__and2_1
XANTENNA__07007__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ net1055 _05105_ _05107_ net833 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__o211a_1
XANTENNA__12532__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1222 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_2
XANTENNA__07963__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1216 net1222 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_2
Xfanout1227 net1255 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_2
Xfanout1238 net1239 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
Xfanout1249 net1253 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_2
Xfanout251 _05650_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xfanout262 net264 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13940_ clknet_leaf_115_clk _00827_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout273 net276 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout284 _05602_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_1
XANTENNA__10314__A2 _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07715__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _05596_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10987__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ clknet_leaf_7_clk _00758_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12822_ net216 net2226 net559 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__mux2_1
XANTENNA__09468__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11391__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ net232 net2538 net568 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__mux2_1
X_11704_ net1404 _06142_ _06144_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12684_ net2068 net237 net431 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
XANTENNA__07494__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14423_ clknet_leaf_45_clk _01310_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11635_ _06087_ _06096_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12707__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09750__B1_N _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07246__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ clknet_leaf_42_clk _01241_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _05300_ _05730_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__nand2_1
XANTENNA__09640__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13305_ clknet_leaf_110_clk _00295_ net1104 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10517_ _05421_ _05424_ _05427_ keypad.alpha vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__and4b_1
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08994__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14285_ clknet_leaf_119_clk _01172_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11497_ net1011 _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__nand2_1
XANTENNA__12008__A datapath.mulitply_result\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10454__C net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13236_ clknet_leaf_78_clk _00226_ net1246 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
X_10448_ _02410_ _02456_ _02499_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__or3_1
XANTENNA__11847__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12442__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ clknet_leaf_5_clk _00159_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10379_ _05279_ _05284_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__nor2_1
X_12118_ datapath.mulitply_result\[23\] datapath.multiplication_module.multiplicand_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__nor2_1
X_13098_ clknet_leaf_9_clk _00090_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ datapath.mulitply_result\[12\] datapath.multiplication_module.multiplicand_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__nand2_1
XANTENNA__10897__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ _01416_ _01479_ _01481_ datapath.ru.latched_instruction\[10\] _01539_ vssd1
+ vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__a221o_1
X_07590_ datapath.rf.registers\[11\]\[16\] net971 net898 datapath.rf.registers\[6\]\[16\]
+ _02516_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__a221o_1
XANTENNA__06676__A _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06541_ _01411_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11266__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11805__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06472_ datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
X_09260_ _03506_ _04173_ _04181_ net611 vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__o31a_1
XFILLER_0_146_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ datapath.rf.registers\[26\]\[2\] net943 net875 datapath.rf.registers\[25\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09191_ net671 _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__or2_1
XANTENNA__12617__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08142_ datapath.rf.registers\[22\]\[3\] net955 net903 datapath.rf.registers\[20\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07237__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ datapath.rf.registers\[28\]\[5\] net718 net717 datapath.rf.registers\[29\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a22o_1
XANTENNA__08985__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07024_ _01930_ net534 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12352__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _03330_ _03873_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a21oi_1
Xhold15 keypad.debounce.debounce\[7\] vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _06449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 screen.register.cFill2 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 datapath.multiplication_module.multiplier_i\[8\] vssd1 vssd1 vccd1 vccd1 net1403
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ datapath.rf.registers\[11\]\[8\] net969 net885 datapath.rf.registers\[9\]\[8\]
+ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a221o_1
Xhold48 net60 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 screen.controlBus\[12\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ _01607_ _01727_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout650_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06808_ _01646_ net977 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__nor2_2
X_07788_ datapath.rf.registers\[14\]\[11\] net799 net766 datapath.rf.registers\[3\]\[11\]
+ _02714_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11257__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ net419 _04453_ net318 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06739_ mmio.memload_or_instruction\[10\] net1061 net1006 datapath.ru.latched_instruction\[10\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__a32oi_4
XANTENNA_fanout915_A _01830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09458_ _04360_ _04383_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__nand2_1
XANTENNA__07476__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__B1_N net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ _02349_ _03335_ _02345_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__o21a_1
XANTENNA__12527__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net361 _04198_ _04199_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11420_ screen.register.currentYbus\[29\] net133 _05895_ net162 vssd1 vssd1 vccd1
+ vccd1 _00387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07228__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__C1 datapath.MemRead vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11351_ mmio.memload_or_instruction\[30\] net1063 net310 net314 datapath.ru.latched_instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08025__B net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__A1 datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10302_ net380 _04365_ _05228_ net331 vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__o211a_1
X_14070_ clknet_leaf_32_clk _00957_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ net33 net1044 net1033 mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1
+ vccd1 _00296_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13021_ clknet_leaf_32_clk _00013_ net1143 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10233_ _05157_ _05158_ _05159_ net1056 net701 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a221o_1
XANTENNA__12262__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06739__A1 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 _01640_ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_2
X_10164_ net203 _05083_ net1310 vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1013 _05729_ vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07400__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_2
Xfanout1057 _03567_ vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_4
X_10095_ net1274 net538 vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__nor2_1
Xfanout1068 net1070 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1085 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_4
X_13923_ clknet_leaf_105_clk _00810_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__B1 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ clknet_leaf_50_clk _00741_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11248__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ net281 net1900 net557 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ clknet_leaf_60_clk _00672_ net1265 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10997_ net285 net2165 net582 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__mux2_1
XANTENNA__10449__C _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ net293 net1537 net566 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07467__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10471__B2 datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ net1581 net181 net432 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XANTENNA__12437__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14406_ clknet_leaf_108_clk _01293_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11618_ net1279 net1280 screen.counter.ct\[22\] _06080_ vssd1 vssd1 vccd1 vccd1 _06081_
+ sky130_fd_sc_hd__and4_1
XANTENNA__09613__B1 _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10465__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ net1673 net167 net445 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
X_14337_ clknet_leaf_45_clk _01224_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11549_ screen.register.currentYbus\[14\] _05736_ _06013_ _06015_ vssd1 vssd1 vccd1
+ vccd1 _06016_ sky130_fd_sc_hd__a211o_1
Xhold507 datapath.rf.registers\[0\]\[28\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 datapath.rf.registers\[10\]\[1\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold529 datapath.rf.registers\[4\]\[21\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ clknet_leaf_52_clk _01155_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09377__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13219_ clknet_leaf_97_clk datapath.multiplication_module.zero_multi net1220 vssd1
+ vssd1 vccd1 vccd1 datapath.ru.zero_multi1 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07774__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ clknet_leaf_45_clk _01086_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1207 datapath.rf.registers\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12900__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08760_ net533 net534 net353 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1218 datapath.rf.registers\[1\]\[29\] vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 screen.register.currentXbus\[20\] vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
X_07711_ datapath.rf.registers\[7\]\[13\] net956 net892 datapath.rf.registers\[14\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a22o_1
X_08691_ net422 _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nor2_1
X_07642_ datapath.rf.registers\[30\]\[14\] net770 net718 datapath.rf.registers\[28\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11239__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07573_ net651 _02499_ _01729_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a21o_1
XANTENNA__08104__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ net506 net505 net360 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__mux2_1
X_06524_ _01405_ datapath.multiplication_module.mul_prev _01453_ vssd1 vssd1 vccd1
+ vccd1 _01454_ sky130_fd_sc_hd__a21o_1
XANTENNA__09510__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06666__B1 _01456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09243_ net516 net356 _04169_ net385 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12347__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout231_A _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06853__B _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09174_ _03991_ _04100_ net396 vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10214__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ datapath.rf.registers\[24\]\[4\] net755 net719 datapath.rf.registers\[28\]\[4\]
+ _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1140_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07091__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ datapath.rf.registers\[7\]\[5\] net956 net888 datapath.rf.registers\[12\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07630__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07007_ datapath.rf.registers\[11\]\[29\] net971 net894 datapath.rf.registers\[14\]\[29\]
+ _01933_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__07918__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout865_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _02431_ net522 net359 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XANTENNA__07904__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ net514 _02833_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__and2_1
X_08889_ net526 net357 _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a21o_1
X_10920_ net172 net2601 net597 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__mux2_1
XANTENNA__07697__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ net1891 net173 net604 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13570_ clknet_leaf_89_clk _00520_ net1214 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07449__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ _01472_ net658 _05616_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06657__B1 _01464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ net2331 net228 net454 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12257__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12452_ net238 net1802 net462 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10285__B _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ net342 net714 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12383_ net254 net1841 net468 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ clknet_leaf_9_clk _01009_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11334_ datapath.ru.latched_instruction\[13\] net314 net309 _01628_ vssd1 vssd1 vccd1
+ vccd1 _00336_ sky130_fd_sc_hd__a22o_1
XANTENNA__07082__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07621__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11397__A _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ clknet_leaf_108_clk _00940_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07594__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ net344 _05844_ net147 net2602 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__a2bb2o_1
X_13004_ net1579 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__clkbuf_1
X_10216_ net701 _04448_ _05137_ _05142_ net205 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a311oi_1
X_11196_ mmio.wishbone.curr_state\[0\] _05252_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__nand2_2
XANTENNA__08582__A0 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10451__D _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12720__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ net1055 _05073_ _05072_ net698 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_128_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ net836 _05002_ _05004_ net206 _05000_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a311o_1
X_13906_ clknet_leaf_34_clk _00793_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10141__B1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__A1_N _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13837_ clknet_leaf_0_clk _00724_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06896__B1 _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13768_ clknet_leaf_13_clk _00655_ net1115 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ net228 net1921 net571 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13699_ clknet_leaf_68_clk datapath.multiplication_module.multiplicand_i_n\[16\]
+ net1226 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13664__RESET_B net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11944__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07073__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 datapath.rf.registers\[22\]\[22\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 datapath.rf.registers\[5\]\[19\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold326 datapath.rf.registers\[5\]\[27\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 datapath.rf.registers\[23\]\[18\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 datapath.rf.registers\[25\]\[6\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ datapath.PC\[30\] _01728_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__or2_1
Xhold359 datapath.rf.registers\[23\]\[16\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout806 net808 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_4
X_09861_ _04735_ _04739_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__xnor2_1
Xfanout817 _01747_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_4
Xfanout828 net830 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_8
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_2
X_08812_ net654 _03732_ _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__or3_1
XANTENNA__12630__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1004 datapath.rf.registers\[2\]\[29\] vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ datapath.PC\[8\] _02877_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and2_1
Xhold1015 datapath.rf.registers\[2\]\[10\] vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 datapath.rf.registers\[23\]\[21\] vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 datapath.rf.registers\[11\]\[12\] vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _01860_ net360 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__or2_1
Xhold1048 datapath.rf.registers\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 datapath.rf.registers\[17\]\[6\] vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout181_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout279_A _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__A2_N _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _03461_ _03463_ net409 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ datapath.rf.registers\[7\]\[15\] net957 net914 datapath.rf.registers\[18\]\[15\]
+ _02551_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07556_ datapath.rf.registers\[24\]\[16\] net757 net721 datapath.rf.registers\[28\]\[16\]
+ _02481_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06507_ net1291 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07487_ datapath.rf.registers\[16\]\[18\] net962 net889 datapath.rf.registers\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ net375 _04151_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07851__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ _03400_ _04082_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12805__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ datapath.rf.registers\[14\]\[4\] net893 net873 datapath.rf.registers\[25\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08800__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07603__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ net517 net518 net356 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ datapath.rf.registers\[19\]\[6\] net759 net722 datapath.rf.registers\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_55_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold860 datapath.rf.registers\[19\]\[23\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold871 datapath.rf.registers\[23\]\[15\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold882 datapath.rf.registers\[1\]\[26\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net1022 _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__nor2_4
Xhold893 datapath.rf.registers\[5\]\[5\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ net837 _04925_ _04927_ net208 _04923_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a311o_1
XANTENNA__12540__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ net285 net1702 net578 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ net257 net1755 net594 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__mux2_1
XANTENNA__10995__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ net157 _05868_ net150 net2387 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13622_ clknet_leaf_115_clk _00560_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10834_ datapath.PC\[17\] _05490_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ clknet_leaf_87_clk _00503_ net1219 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ net839 _04191_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__nand2_1
XANTENNA__08095__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12504_ net2281 net297 net452 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13484_ clknet_leaf_82_clk _00437_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07842__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10696_ datapath.PC\[27\] _05538_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12435_ _05478_ _05479_ net577 vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12715__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11926__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10729__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07055__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_73_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12366_ net1943 net171 net474 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14105_ clknet_leaf_48_clk _00992_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11317_ _01671_ _05855_ _05853_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12297_ net2349 net186 net482 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__mux2_1
XANTENNA__10462__C net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ clknet_leaf_113_clk _00923_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09347__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ net1486 net141 net135 _02633_ vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__a22o_1
XANTENNA__12450__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ keypad.decode.sticky_n\[2\] keypad.decode.sticky_n\[3\] _05827_ vssd1 vssd1
+ vccd1 vccd1 _05828_ sky130_fd_sc_hd__nor3_4
XANTENNA__08307__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09044__B _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08858__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07410_ datapath.rf.registers\[18\]\[20\] net915 net866 datapath.rf.registers\[13\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08390_ _02978_ _03019_ _03315_ _02973_ net510 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09060__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ datapath.rf.registers\[14\]\[21\] net800 net779 datapath.rf.registers\[9\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
XANTENNA__08086__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07294__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ datapath.rf.registers\[3\]\[23\] net966 net945 datapath.rf.registers\[19\]\[23\]
+ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a221o_1
XANTENNA__07833__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _03552_ net635 _03927_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_154_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12625__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07046__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 screen.controlBus\[11\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 screen.controlBus\[16\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 screen.counter.currentCt\[9\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _00478_ vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 net115 vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 datapath.rf.registers\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 net120 vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 keypad.apps.app_c\[0\] vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _04838_ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__xnor2_1
Xhold189 datapath.rf.registers\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout603 net604 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout614 _03554_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout625 _03356_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _03559_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_2
Xfanout647 net649 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_4
X_09844_ datapath.PC\[23\] net629 vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12360__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_4
Xfanout669 _05695_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_2
X_09775_ datapath.PC\[13\] net632 _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout563_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ datapath.rf.registers\[22\]\[29\] net753 net732 datapath.rf.registers\[16\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
XANTENNA__06578__B _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ net521 net520 net404 vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__mux2_1
XANTENNA__08849__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ datapath.PC\[21\] _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout730_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07608_ datapath.rf.registers\[14\]\[15\] net800 net756 datapath.rf.registers\[24\]\[15\]
+ _02528_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a221o_1
X_08588_ _01657_ _03121_ _03507_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ datapath.rf.registers\[7\]\[17\] net956 net924 datapath.rf.registers\[8\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10550_ _05415_ _05455_ net1025 vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07824__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ net498 net495 net510 vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__a21o_1
XANTENNA__09026__A1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ screen.register.currentYbus\[17\] screen.register.currentYbus\[16\] screen.register.currentYbus\[19\]
+ screen.register.currentYbus\[18\] vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__or4_1
XANTENNA__12535__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07037__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12220_ net242 net1885 net575 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08785__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _06409_ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__or2_1
X_11102_ net1296 net1295 vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__nand2_2
X_12082_ datapath.mulitply_result\[17\] datapath.multiplication_module.multiplicand_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__and2_1
Xhold690 datapath.rf.registers\[7\]\[27\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__A0 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11033_ _05314_ _05321_ _05328_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__and4_1
XANTENNA__12270__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__A2 _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12984_ net1593 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11935_ net153 _05887_ net128 net2634 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ net705 _04860_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13605_ clknet_leaf_107_clk _00543_ net1110 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10817_ _05489_ _05646_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__nor2_1
XANTENNA__08068__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ datapath.PC\[10\] net302 _06203_ _06205_ vssd1 vssd1 vccd1 vccd1 _00454_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ clknet_leaf_80_clk _00486_ net1234 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07276__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07112__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07815__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ datapath.mulitply_result\[3\] net426 _05587_ _05588_ net659 vssd1 vssd1 vccd1
+ vccd1 _05589_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13467_ clknet_leaf_80_clk net714 net1239 vssd1 vssd1 vccd1 vccd1 screen.counter.ack1
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09017__A1 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12445__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ _01473_ net660 _05529_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07028__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12418_ net2036 net245 net465 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
X_13398_ clknet_leaf_92_clk _00003_ net1202 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12349_ net1999 net258 net472 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__mux2_1
XANTENNA__08240__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14019_ clknet_leaf_104_clk _00906_ net1115 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_06910_ datapath.rf.registers\[2\]\[31\] net921 net897 datapath.rf.registers\[6\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
X_07890_ datapath.rf.registers\[11\]\[9\] net775 net756 datapath.rf.registers\[24\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a22o_1
X_06841_ datapath.rf.registers\[3\]\[31\] net768 net764 datapath.rf.registers\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ _03529_ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__nand2_1
X_06772_ datapath.ru.latched_instruction\[4\] _01593_ _01624_ datapath.ru.latched_instruction\[14\]
+ _01683_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a221o_1
XANTENNA__06829__D _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08511_ _01909_ _03437_ _01907_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a21bo_1
X_09491_ _04047_ _04081_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__or3_1
XANTENNA__10638__B2 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08442_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08373_ datapath.rf.registers\[7\]\[0\] net956 net891 datapath.rf.registers\[12\]\[0\]
+ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a221o_1
XANTENNA__08059__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout144_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07267__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ _02244_ _02246_ _02248_ _02250_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07806__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07255_ datapath.rf.registers\[5\]\[23\] net784 net763 datapath.rf.registers\[17\]\[23\]
+ _02173_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout311_A _05859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12355__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1053_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07019__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07186_ datapath.rf.registers\[16\]\[25\] net963 net934 datapath.rf.registers\[23\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout400 _03515_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout778_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _03450_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 net435 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_8
Xfanout444 net447 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_8
Xfanout455 _06458_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_8
X_09827_ _04714_ _04717_ _04752_ _04713_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a31o_1
Xfanout477 _06452_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_107_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 net490 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
XANTENNA_fanout945_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_2
X_09758_ _04683_ _04684_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__nor2_1
XANTENNA__06950__C1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _03600_ _03632_ _03633_ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a31o_1
X_09689_ _02932_ _02978_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ net1294 _06068_ screen.counter.ct\[7\] vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_120_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11651_ _06108_ _06109_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10602_ net1547 net519 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[14\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ clknet_leaf_33_clk _01257_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11582_ net1287 net1288 screen.counter.ct\[19\] net1282 vssd1 vssd1 vccd1 vccd1 _06046_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13321_ clknet_leaf_111_clk _00311_ net1103 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_10533_ _05413_ _05440_ _05423_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a21o_1
XANTENNA__12265__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_65_clk _00242_ net1269 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ _02079_ net531 net529 net528 vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ net287 net2217 net573 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__mux2_1
XANTENNA__08758__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ clknet_leaf_37_clk _00175_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ screen.counter.ct\[6\] net1291 net1284 net1280 _05298_ vssd1 vssd1 vccd1
+ vccd1 _05317_ sky130_fd_sc_hd__a41o_1
XANTENNA__07430__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ datapath.mulitply_result\[25\] net327 net323 _06396_ vssd1 vssd1 vccd1 vccd1
+ _00600_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12065_ _06331_ _06338_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__or2_1
X_11016_ net210 net2275 net585 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA__09306__C net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11817__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ net294 net2504 net606 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11918_ net153 _05870_ net128 screen.register.currentXbus\[4\] vssd1 vssd1 vccd1
+ vccd1 _00515_ sky130_fd_sc_hd__a22o_1
X_12898_ net1529 net182 net545 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ _06242_ datapath.PC\[25\] net304 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14568_ net1338 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_16_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13519_ clknet_leaf_64_clk _00469_ net1270 vssd1 vssd1 vccd1 vccd1 datapath.PC\[25\]
+ sky130_fd_sc_hd__dfstp_2
X_14499_ clknet_leaf_105_clk _01386_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06681__B net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07040_ datapath.rf.registers\[7\]\[28\] net825 net784 datapath.rf.registers\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08213__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12903__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08991_ net372 _03805_ _03806_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_10_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07942_ datapath.rf.registers\[15\]\[8\] net808 net726 datapath.rf.registers\[2\]\[8\]
+ _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_149_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A2 _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ datapath.rf.registers\[30\]\[9\] net910 net886 datapath.rf.registers\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__a22o_1
X_09612_ net673 _04536_ _04538_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__and3_1
X_06824_ net987 _01734_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__and2_1
X_09543_ _04451_ _04465_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__o21ai_1
X_06755_ datapath.ru.latched_instruction\[20\] net1039 net1006 _01680_ vssd1 vssd1
+ vccd1 vccd1 _01682_ sky130_fd_sc_hd__a22o_4
XANTENNA__09477__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06856__B _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07488__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net396 _04171_ _04264_ net399 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06686_ _01488_ net1030 net1008 net1041 datapath.ru.latched_instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a32oi_4
XANTENNA__11284__B2 mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08425_ _01864_ _03351_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1170_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_A _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ datapath.rf.registers\[24\]\[0\] net758 _03256_ _03257_ _03267_ vssd1 vssd1
+ vccd1 vccd1 _03283_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_82_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07307_ datapath.rf.registers\[0\]\[22\] net829 _02233_ vssd1 vssd1 vccd1 vccd1 _02234_
+ sky130_fd_sc_hd__o21ai_4
X_08287_ datapath.rf.registers\[9\]\[1\] net995 _01754_ vssd1 vssd1 vccd1 vccd1 _03214_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_117_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07238_ datapath.rf.registers\[19\]\[24\] net946 net942 datapath.rf.registers\[26\]\[24\]
+ _02164_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08204__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12813__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07169_ datapath.rf.registers\[15\]\[25\] net807 net776 datapath.rf.registers\[11\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a22o_1
XANTENNA__07412__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _03575_ _05106_ net1051 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a21o_1
Xfanout1206 net1208 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_4
Xfanout1217 net1218 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_4
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout230 _05508_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 _05660_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xfanout1239 net1242 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
Xfanout252 _05650_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_89_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
Xfanout274 net276 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_89_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout285 _05602_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
Xfanout296 _05596_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ clknet_leaf_1_clk _00757_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07191__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net219 net2353 net559 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12752_ net226 net2342 net565 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__mux2_1
XANTENNA__11275__B2 mmio.memload_or_instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ net1404 _06142_ net666 vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__o21ai_1
X_12683_ net1724 net239 net434 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14422_ clknet_leaf_32_clk _01309_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11634_ screen.counter.ct\[22\] _06074_ net1019 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_37_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14353_ clknet_leaf_9_clk _01240_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11565_ net1533 _05901_ _06030_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__o21a_1
XANTENNA__07597__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ clknet_leaf_112_clk _00294_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10516_ _05425_ _05426_ net1050 _05401_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_122_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07651__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14284_ clknet_leaf_30_clk _01171_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11496_ screen.register.currentYbus\[27\] _05777_ _05954_ _05963_ _05965_ vssd1 vssd1
+ vccd1 vccd1 _05966_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire697 _01828_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_1
X_13235_ clknet_leaf_76_clk _00225_ net1248 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
X_10447_ _02587_ _02633_ _02677_ _02721_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12723__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ clknet_leaf_118_clk _00158_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09943__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10378_ _05294_ _05297_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__or2_2
X_12117_ datapath.mulitply_result\[23\] datapath.multiplication_module.multiplicand_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__and2_1
X_13097_ clknet_leaf_3_clk _00089_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08221__B net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ net321 _06323_ _06324_ net325 net1804 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a32o_1
XANTENNA__07706__A1 _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07182__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06676__B net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ clknet_leaf_7_clk _00886_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_06540_ mmio.memload_or_instruction\[7\] net1058 vssd1 vssd1 vccd1 vccd1 _01470_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10069__A2 _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11266__B2 _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10198__B _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08210_ datapath.rf.registers\[4\]\[2\] net929 net861 datapath.rf.registers\[28\]\[2\]
+ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09190_ _02978_ _03397_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07890__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ _03064_ _03066_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ datapath.rf.registers\[7\]\[5\] net824 net817 datapath.rf.registers\[31\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
XANTENNA__07642__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06996__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ datapath.rf.registers\[0\]\[29\] net693 _01937_ _01949_ vssd1 vssd1 vccd1
+ vccd1 _01950_ sky130_fd_sc_hd__o22a_2
XFILLER_0_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07727__S net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08974_ net708 _03900_ net491 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__o21a_1
Xhold16 keypad.debounce.debounce\[1\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold27 datapath.ru.n_memread vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ datapath.rf.registers\[4\]\[8\] net929 net923 datapath.rf.registers\[2\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a22o_1
Xhold38 screen.counter.currentCt\[22\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 net110 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13359__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A _06452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _02767_ _02768_ _02782_ net827 datapath.rf.registers\[0\]\[10\] vssd1 vssd1
+ vccd1 vccd1 _02783_ sky130_fd_sc_hd__o32a_4
XANTENNA__07173__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ _01639_ net998 _01656_ net977 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__and4_4
X_07787_ datapath.rf.registers\[7\]\[11\] net824 net820 datapath.rf.registers\[26\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ _04430_ _04452_ net412 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__mux2_1
X_06738_ _01664_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09457_ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__inv_2
X_06669_ _01592_ _01593_ _01595_ _01596_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__and4_2
XANTENNA_fanout810_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12808__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_A _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06684__A1 _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ _02390_ _03334_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ net317 _03753_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07881__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08339_ datapath.rf.registers\[9\]\[0\] net995 _01754_ vssd1 vssd1 vccd1 vccd1 _03266_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_151_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ datapath.ru.latched_instruction\[29\] net314 net310 _01615_ vssd1 vssd1 vccd1
+ vccd1 _00352_ sky130_fd_sc_hd__a22o_1
XANTENNA__07633__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06987__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ net380 _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__nand2_1
X_11281_ net32 net1046 net1035 mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1
+ vccd1 _00295_ sky130_fd_sc_hd__a22o_1
XANTENNA__12543__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13020_ clknet_leaf_53_clk _00012_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10232_ datapath.PC\[14\] _03577_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ _05085_ _05089_ net200 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__o21a_1
Xfanout1014 _05727_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__buf_2
Xfanout1025 _05417_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
Xfanout1036 _05847_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input37_A gpio_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 _05845_ vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10998__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _04833_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__or2_1
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_2
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_2
X_13922_ clknet_leaf_43_clk _00809_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13853_ clknet_leaf_24_clk _00740_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ net285 net2002 net557 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
XANTENNA__11248__B2 _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ clknet_leaf_39_clk _00671_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10996_ net296 net1699 net583 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08992__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08113__B2 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12735_ net298 net1607 net566 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12718__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12666_ _05669_ _05671_ net577 vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__nor3_2
XFILLER_0_154_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10746__B _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ net1284 net1281 net1282 _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__and4_1
X_14405_ clknet_leaf_107_clk _01292_ net1110 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ net2493 net171 net446 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12019__A datapath.mulitply_result\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10465__C _02997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07624__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ screen.register.currentXbus\[14\] net1016 _06014_ vssd1 vssd1 vccd1 vccd1
+ _06015_ sky130_fd_sc_hd__a21o_1
X_14336_ clknet_leaf_46_clk _01223_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold508 datapath.rf.registers\[15\]\[27\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12453__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14267_ clknet_leaf_19_clk _01154_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold519 datapath.rf.registers\[1\]\[18\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ net1017 _05949_ _05931_ _05918_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a211o_1
X_13218_ clknet_leaf_33_clk _00210_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14198_ clknet_leaf_26_clk _01085_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13149_ clknet_leaf_32_clk _00141_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1208 datapath.rf.registers\[31\]\[20\] vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 screen.register.currentXbus\[24\] vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ datapath.rf.registers\[31\]\[13\] net948 net860 datapath.rf.registers\[28\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
X_08690_ _03615_ _03616_ net414 vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__mux2_1
XANTENNA__06687__A mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__C1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07641_ _02546_ net520 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11239__B2 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07572_ datapath.rf.registers\[0\]\[16\] _02498_ net829 vssd1 vssd1 vccd1 vccd1 _02499_
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09311_ net498 net495 net508 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__a21o_1
X_06523_ datapath.ru.n_memread datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 _01453_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_146_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ net500 net621 net489 net515 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09173_ _04098_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__nand2_1
X_08124_ datapath.rf.registers\[21\]\[4\] net744 net725 datapath.rf.registers\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07615__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ datapath.rf.registers\[2\]\[5\] net923 net916 datapath.rf.registers\[10\]\[5\]
+ _02981_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12363__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ datapath.rf.registers\[6\]\[29\] net898 net887 datapath.rf.registers\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout593_A _05673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08040__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08591__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ net375 _03766_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout858_A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__inv_2
X_08888_ net500 net621 net489 net524 vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__o211a_1
XANTENNA__07146__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ datapath.rf.registers\[17\]\[10\] net765 net726 datapath.rf.registers\[2\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a22o_1
X_10850_ net1608 net185 net603 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06564__C_N mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09509_ _03484_ _04433_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12538__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ datapath.mulitply_result\[8\] net426 net658 vssd1 vssd1 vccd1 vccd1 _05617_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12520_ net1979 net243 net454 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net247 net1985 net461 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XANTENNA__10058__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ screen.register.currentYbus\[20\] net132 _05886_ net161 vssd1 vssd1 vccd1
+ vccd1 _00378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07606__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ net259 net2075 net468 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14121_ clknet_leaf_2_clk _01008_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11333_ _01509_ net1031 net308 net312 datapath.ru.latched_instruction\[12\] vssd1
+ vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12273__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ clknet_leaf_14_clk _00939_ net1115 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11397__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ net535 _05844_ net147 net94 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__a2bb2o_1
X_13003_ net2607 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__clkbuf_1
X_10215_ net701 _05141_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__nor2_1
XANTENNA__08031__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ net2251 _05828_ _05837_ vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__a21o_1
XANTENNA__07385__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ datapath.PC\[5\] _03571_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ _03588_ _05003_ net1052 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a21o_1
XANTENNA__07137__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ clknet_leaf_8_clk _00792_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10141__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13836_ clknet_leaf_31_clk _00723_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08098__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12448__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13767_ clknet_leaf_18_clk _00654_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08637__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ net230 net2579 net588 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07845__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ net243 net2453 net569 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13698_ clknet_leaf_68_clk datapath.multiplication_module.multiplicand_i_n\[15\]
+ net1223 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09047__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12649_ net247 net2327 net437 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold305 datapath.rf.registers\[22\]\[3\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ clknet_leaf_3_clk _01206_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08270__B1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 datapath.rf.registers\[4\]\[16\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 datapath.rf.registers\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 datapath.rf.registers\[28\]\[15\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 datapath.rf.registers\[23\]\[24\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
X_09860_ _04715_ _04753_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__xor2_1
Xfanout807 net808 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12911__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08897__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 _01747_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_4
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_6
X_08811_ net319 _03733_ _03734_ _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__a31o_1
X_09791_ net1277 _02832_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__and2_1
Xhold1005 datapath.rf.registers\[26\]\[20\] vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 datapath.rf.registers\[14\]\[5\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 datapath.rf.registers\[23\]\[5\] vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ net317 _03668_ _03652_ _03650_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__o211a_1
Xhold1038 datapath.rf.registers\[11\]\[22\] vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 datapath.rf.registers\[30\]\[17\] vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08673_ net689 _03597_ _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__a21o_1
XANTENNA__10132__A1 _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_A _05562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07624_ datapath.rf.registers\[11\]\[15\] net970 net865 datapath.rf.registers\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07025__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07555_ datapath.rf.registers\[26\]\[16\] net822 net791 datapath.rf.registers\[18\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ net1294 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ datapath.rf.registers\[22\]\[18\] net953 net853 datapath.rf.registers\[5\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a22o_1
XANTENNA__08137__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07300__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ _03679_ _03680_ net368 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _03319_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_79_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08107_ datapath.rf.registers\[22\]\[4\] net953 net905 datapath.rf.registers\[24\]\[4\]
+ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a221o_1
XANTENNA__08261__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ net520 net357 _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_110_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_2_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08038_ datapath.rf.registers\[10\]\[6\] net748 net726 datapath.rf.registers\[2\]\[6\]
+ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold850 datapath.rf.registers\[26\]\[6\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 datapath.rf.registers\[18\]\[12\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08303__C _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08013__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 datapath.rf.registers\[30\]\[8\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 datapath.rf.registers\[24\]\[6\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12821__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 datapath.rf.registers\[7\]\[29\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07367__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ _03585_ _04926_ net1057 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__o21ai_1
X_09989_ _04914_ _04915_ net208 _04913_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a211o_1
XANTENNA__07119__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ net296 net1955 net579 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ net263 net2211 net594 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__mux2_1
X_11882_ net157 _05867_ net150 screen.controlBus\[1\] vssd1 vssd1 vccd1 vccd1 _00480_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13621_ clknet_leaf_48_clk _00559_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10833_ net2446 net240 net604 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ clknet_leaf_79_clk _00502_ net1233 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07827__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ net1800 net283 net602 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08047__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ net1884 net287 net452 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13483_ clknet_leaf_82_clk _00436_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net192 net2367 net607 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12434_ net2109 net165 net465 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12365_ net2082 net184 net473 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_101_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11316_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__inv_2
X_14104_ clknet_leaf_37_clk _00991_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ net1850 net191 net483 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__mux2_1
X_14035_ clknet_leaf_59_clk _00922_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10462__D _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ net1559 net142 net134 _02677_ vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__a22o_1
XANTENNA__12731__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ keypad.decode.sticky\[1\] keypad.decode.sticky\[2\] _01450_ keypad.decode.push
+ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__or4b_1
X_10129_ _04799_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__nand2_1
XANTENNA__11311__A0 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A1 _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10665__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__A2 _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ clknet_leaf_55_clk _00706_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10487__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07340_ datapath.rf.registers\[30\]\[21\] net771 net720 datapath.rf.registers\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__B _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07271_ datapath.rf.registers\[17\]\[23\] net882 net850 datapath.rf.registers\[1\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12906__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11810__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09010_ _03513_ _03936_ _03928_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08243__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold102 net99 vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 datapath.rf.registers\[0\]\[18\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 datapath.multiplication_module.multiplicand_i\[23\] vssd1 vssd1 vccd1 vccd1
+ net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 datapath.rf.registers\[27\]\[0\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 datapath.multiplication_module.multiplicand_i\[19\] vssd1 vssd1 vccd1 vccd1
+ net1512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 datapath.rf.registers\[11\]\[0\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 screen.counter.currentCt\[12\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 net81 vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09912_ datapath.PC\[27\] net628 vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12641__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07349__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_2
Xfanout626 _01730_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
X_09843_ datapath.PC\[22\] net629 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__xnor2_2
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_2
Xfanout648 net649 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11550__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 datapath.MemRead vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_4
X_09774_ _01631_ _04678_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nor2_1
X_06986_ datapath.rf.registers\[17\]\[29\] net764 net716 datapath.rf.registers\[29\]\[29\]
+ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a221o_1
X_08725_ _02169_ net686 net678 _02172_ _03651_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__o221a_1
XANTENNA__11302__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ datapath.PC\[20\] _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ datapath.rf.registers\[26\]\[15\] net821 net720 datapath.rf.registers\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a22o_1
X_08587_ _01656_ _03120_ _03507_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout723_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07538_ datapath.rf.registers\[11\]\[17\] net968 net940 datapath.rf.registers\[26\]\[17\]
+ _02464_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a221o_1
XANTENNA__07809__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07469_ datapath.rf.registers\[9\]\[18\] net779 net771 datapath.rf.registers\[30\]\[18\]
+ _02395_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12816__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ net502 net618 net496 net512 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10480_ screen.register.currentYbus\[21\] screen.register.currentYbus\[20\] screen.register.currentYbus\[23\]
+ screen.register.currentYbus\[22\] vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09139_ _02698_ net516 _03545_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__mux2_1
XANTENNA__09431__C1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _06402_ _06404_ _06403_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10592__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ net1280 screen.counter.ct\[22\] net1279 vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__or3b_1
X_12081_ _06347_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12551__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 datapath.rf.registers\[1\]\[23\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 datapath.rf.registers\[12\]\[24\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ net1299 _05307_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07760__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ net1472 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__clkbuf_1
X_11934_ net153 _05886_ net128 net2595 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__a22o_1
XANTENNA__07512__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11865_ net705 _04608_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13604_ clknet_leaf_97_clk net659 net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memread
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ datapath.PC\[14\] _05488_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nor2_1
X_11796_ _05625_ net175 _06204_ net177 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13535_ clknet_leaf_80_clk _00485_ net1234 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ net840 _05170_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or2_1
XANTENNA__12726__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13466_ clknet_leaf_81_clk _00422_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10678_ datapath.mulitply_result\[24\] net427 net660 vssd1 vssd1 vccd1 vccd1 _05530_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_136_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12417_ net1588 net252 net464 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__mux2_1
X_13397_ clknet_leaf_92_clk net1378 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08224__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07579__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ net1834 net262 net472 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__mux2_1
XANTENNA__10583__A1 _02721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net2358 net267 net480 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__mux2_1
XANTENNA__12461__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08528__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ clknet_leaf_43_clk _00905_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06840_ _01735_ net972 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__and2_2
XFILLER_0_156_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__A2 _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06771_ datapath.ru.latched_instruction\[15\] _01653_ _01662_ datapath.ru.latched_instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a22o_1
X_08510_ _03435_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__nor2_1
X_09490_ _04386_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08441_ _02281_ _02301_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08372_ datapath.rf.registers\[29\]\[0\] net877 net857 datapath.rf.registers\[15\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07323_ datapath.rf.registers\[7\]\[22\] net958 net882 datapath.rf.registers\[17\]\[22\]
+ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a221o_1
XANTENNA__12636__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout137_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07254_ datapath.rf.registers\[25\]\[23\] net797 net756 datapath.rf.registers\[24\]\[23\]
+ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08216__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ datapath.rf.registers\[30\]\[25\] net911 net854 datapath.rf.registers\[5\]\[25\]
+ _02107_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout304_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12371__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout401 net403 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
XANTENNA__07990__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 _03454_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout434 _06463_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
Xfanout445 net447 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_4
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout456 net459 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_6
X_09826_ _04717_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__nand2_1
Xfanout467 _06455_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_4
Xfanout478 _06452_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout840_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ net1275 net633 _04682_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__nor3_1
X_06969_ datapath.rf.registers\[19\]\[30\] net945 net914 datapath.rf.registers\[18\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout938_A _01817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08708_ net615 _03620_ _03634_ net493 _03597_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a32o_1
X_09688_ _03127_ _03182_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _03440_ net673 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__or2_1
X_11650_ net2391 _06106_ net666 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_25_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ net1563 net518 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[13\]
+ sky130_fd_sc_hd__mux2_1
X_11581_ _06041_ screen.dcx _06045_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12546__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ _05416_ net1025 _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__or3b_1
X_13320_ clknet_leaf_113_clk _00310_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10801__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08207__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13251_ clknet_leaf_65_clk _00241_ net1268 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
X_10463_ _05374_ _05375_ _05376_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_118_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09404__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ net180 net2058 net574 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__mux2_1
X_13182_ clknet_leaf_51_clk _00174_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10394_ net1296 screen.counter.ct\[10\] net1287 _05294_ vssd1 vssd1 vccd1 vccd1 _05316_
+ sky130_fd_sc_hd__and4_1
X_12133_ _06392_ _06395_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12281__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07981__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _06330_ _06332_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__nor2_1
X_11015_ net213 net2463 net584 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
XANTENNA__07194__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 net991 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07733__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06941__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ net293 net1896 net609 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__mux2_1
X_11917_ net151 _05869_ net126 net2614 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__a22o_1
XANTENNA__08694__A0 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ net631 _05666_ _06450_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__nor3_1
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11848_ _04663_ _05534_ _06241_ _04940_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_138_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13477__RESET_B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14567_ net1337 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA__12456__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ net698 _04796_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13518_ clknet_leaf_64_clk _00468_ net1268 vssd1 vssd1 vccd1 vccd1 datapath.PC\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_14498_ clknet_leaf_51_clk _01385_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13449_ clknet_leaf_81_clk _00405_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08990_ net369 _03676_ _03683_ net380 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_71_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07941_ datapath.rf.registers\[18\]\[8\] net789 net730 datapath.rf.registers\[16\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a22o_1
XANTENNA__10308__A1 _05234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ datapath.rf.registers\[25\]\[9\] net873 _02794_ _02796_ _02798_ vssd1 vssd1
+ vccd1 vccd1 _02799_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09713__A3 _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07185__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ net614 _04530_ _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__or3_1
X_06823_ net993 _01746_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__and2_1
X_06754_ datapath.ru.latched_instruction\[20\] net1039 net1006 _01680_ vssd1 vssd1
+ vccd1 vccd1 _01681_ sky130_fd_sc_hd__a22oi_4
X_09542_ _04464_ _04466_ _04468_ net673 vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__o211a_1
XANTENNA__09477__A2 _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09154__A1_N net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06685_ mmio.memload_or_instruction\[26\] net1063 net1010 datapath.ru.latched_instruction\[26\]
+ net1041 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a32oi_4
XANTENNA__11284__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ net391 _04178_ _04255_ net402 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_90_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08424_ _01910_ _01952_ _03349_ _01906_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_22_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08355_ datapath.rf.registers\[6\]\[0\] net816 _03269_ _03272_ _03273_ vssd1 vssd1
+ vccd1 vccd1 _03282_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_82_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1163_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout519_A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _02217_ _02218_ _02232_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08286_ datapath.rf.registers\[27\]\[1\] net990 _01763_ vssd1 vssd1 vccd1 vccd1 _03213_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_117_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06999__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07237_ datapath.rf.registers\[3\]\[24\] net966 net958 datapath.rf.registers\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07168_ datapath.rf.registers\[23\]\[25\] net788 net757 datapath.rf.registers\[24\]\[25\]
+ _02094_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout790_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07099_ datapath.rf.registers\[18\]\[27\] net915 net890 datapath.rf.registers\[12\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
XANTENNA__07963__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1207 net1208 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_2
Xfanout1218 net1222 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_2
Xfanout220 _04662_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_4
Xfanout1229 net1255 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_2
Xfanout231 _05508_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_1
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
Xfanout253 net256 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
Xfanout264 _05634_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_89_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
XANTENNA__07715__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 _05602_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_1
Xfanout297 net300 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
X_09809_ _03208_ _03209_ datapath.PC\[1\] vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__o21a_1
X_12820_ net222 net2571 net558 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__mux2_1
X_12751_ net244 net2221 net567 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_81_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
X_11702_ net666 _06141_ _06143_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__and3_1
X_12682_ net1830 net246 net433 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
X_14421_ clknet_leaf_27_clk _01308_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11633_ _06089_ _06090_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nor3_1
XANTENNA__12276__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ clknet_leaf_4_clk _01239_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ _05987_ _06024_ _06029_ net1017 _05902_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__a221o_1
XANTENNA__07100__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire643 _03294_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_1
XFILLER_0_64_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13303_ clknet_leaf_112_clk _00293_ net1104 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ net1026 _05423_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__or2_1
X_11495_ screen.register.currentYbus\[11\] _05776_ _05964_ vssd1 vssd1 vccd1 vccd1
+ _05965_ sky130_fd_sc_hd__a21o_1
X_14283_ clknet_leaf_18_clk _01170_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10446_ net424 net530 vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__nand2_1
X_13234_ clknet_leaf_77_clk _00224_ net1247 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ clknet_leaf_119_clk _00157_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10377_ _05294_ _05297_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12116_ net323 _06380_ _06381_ net327 net1991 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__a32o_1
X_13096_ clknet_leaf_13_clk _00088_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12047_ _06320_ _06321_ _06322_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__or3_1
XANTENNA__07167__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_148_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ clknet_leaf_116_clk _00885_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11266__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ _05496_ net1703 net543 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08131__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10495__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10226__B1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08140_ _03064_ _03066_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__or2_1
XANTENNA__10777__A1 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08071_ net847 _01726_ _01606_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12914__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07022_ net695 _01939_ _01948_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__or3_1
XFILLER_0_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09395__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap976 _01803_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_1
XFILLER_0_140_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap998 _01645_ vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__buf_4
X_08973_ net653 _03882_ _03890_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__or4_1
Xhold17 screen.screenEdge.enable2 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold28 datapath.pc_module.i_ack1 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ datapath.rf.registers\[7\]\[8\] net958 net946 datapath.rf.registers\[19\]\[8\]
+ _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a221o_1
Xhold39 net54 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _02770_ _02772_ _02775_ _02781_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or4_1
XANTENNA__06905__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__A2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06806_ _01638_ net982 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nor2_1
X_07786_ _02707_ _02708_ _02710_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ _03653_ _03661_ net341 vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06737_ _01518_ net1031 net1007 net1043 datapath.ru.latched_instruction\[11\] vssd1
+ vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_94_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08122__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06668_ _01595_ _01596_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__nand2_1
X_09456_ net670 _04361_ _04378_ _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o22a_2
XFILLER_0_148_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08407_ _02437_ _02478_ _03331_ _02433_ _02391_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__o311a_1
X_06599_ _01467_ _01469_ _01525_ _01528_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__or4b_1
X_09387_ _03020_ net687 net679 _04311_ _04313_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ datapath.rf.registers\[13\]\[0\] net994 _01756_ vssd1 vssd1 vccd1 vccd1 _03265_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09083__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__A1 datapath.mulitply_result\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08269_ datapath.rf.registers\[4\]\[1\] net929 net920 datapath.rf.registers\[2\]\[1\]
+ _03191_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a221o_1
XANTENNA__12824__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10300_ net369 _04283_ _04284_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net31 net1044 net1033 net2608 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__o22a_1
XANTENNA__08603__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08189__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ datapath.PC\[14\] net537 net1051 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07397__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ net1055 _05086_ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__o21ba_1
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
Xfanout1015 _05727_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_2
Xfanout1026 _05416_ vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_2
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_4
X_10093_ _04780_ _04832_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__nor2_1
XANTENNA__07149__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1060 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_2
X_13921_ clknet_leaf_42_clk _00808_ net1162 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08361__A2 _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ clknet_leaf_54_clk _00739_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12803_ net296 net1688 net559 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__mux2_1
X_13783_ clknet_leaf_45_clk _00670_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ net292 net1756 net583 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12734_ net287 net1867 net565 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07321__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12665_ net164 net2470 net437 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
X_14404_ clknet_leaf_16_clk _01291_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11616_ net1287 net1289 net1286 _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_13_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__B1 _03998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ net1640 net185 net445 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10465__D _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14335_ clknet_leaf_38_clk _01222_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11547_ screen.register.currentYbus\[6\] _05737_ _05742_ screen.register.currentYbus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__a22o_1
XANTENNA__12734__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold509 datapath.rf.registers\[9\]\[14\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ clknet_leaf_23_clk _01153_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11478_ screen.register.currentYbus\[26\] _05742_ _05945_ _05947_ _05948_ vssd1 vssd1
+ vccd1 vccd1 _05949_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_40_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13217_ clknet_leaf_45_clk _00209_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ _05345_ _05347_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__or2_1
X_14197_ clknet_leaf_28_clk _01084_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07388__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06595__A2_N _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ clknet_leaf_57_clk _00140_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13079_ clknet_leaf_45_clk _00071_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1209 mmio.memload_or_instruction\[31\] vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11487__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07640_ _02546_ net520 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07560__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07571_ datapath.rf.registers\[9\]\[16\] net780 _02494_ _02496_ _02497_ vssd1 vssd1
+ vccd1 vccd1 _02498_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12909__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08104__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06522_ datapath.ru.n_memread datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 _01452_
+ sky130_fd_sc_hd__nor2_1
X_09310_ net509 net360 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07312__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _04166_ _04167_ net391 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09172_ _02698_ net354 _04057_ net390 vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _03043_ _03045_ _03047_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__or4_1
XANTENNA__12644__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ datapath.rf.registers\[20\]\[5\] net900 _02980_ net696 vssd1 vssd1 vccd1
+ vccd1 _02981_ sky130_fd_sc_hd__a211o_1
XANTENNA__07091__A2 _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ datapath.rf.registers\[2\]\[29\] net922 net915 datapath.rf.registers\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07379__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout586_A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08956_ net362 _03621_ _03622_ net371 vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o211a_1
X_07907_ net514 _02833_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__or2_2
XANTENNA__11478__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10135__C1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net500 net621 net489 net527 vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o211a_1
XANTENNA__06597__B _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10686__B1 _05535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07000__C1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ datapath.rf.registers\[15\]\[10\] net805 net799 datapath.rf.registers\[14\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout920_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _02689_ _02691_ _02693_ _02695_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__or4_1
XANTENNA__12819__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
X_09508_ _02610_ net687 net679 _02614_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__o221a_1
X_10780_ _04384_ _05615_ net844 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__mux2_1
XANTENNA__07303__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09439_ _03925_ _04365_ net380 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12450_ net250 net2170 net461 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ net525 screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11402__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ net262 net2598 net468 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__mux2_1
XANTENNA__12554__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14120_ clknet_leaf_12_clk _01007_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11332_ _01518_ net1027 net308 net312 datapath.ru.latched_instruction\[11\] vssd1
+ vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__a32o_1
XANTENNA__09429__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07082__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ clknet_leaf_104_clk _00938_ net1115 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ net425 _05844_ net147 net93 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__a2bb2o_1
X_13002_ net1530 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__clkbuf_1
X_10214_ net1056 _05138_ _05139_ _05140_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__o22a_1
X_11194_ mmio.key_data\[6\] net220 _05829_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__and3_1
X_10145_ datapath.PC\[5\] net536 net1051 _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__o211a_1
XANTENNA__10802__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06788__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07790__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10076_ datapath.PC\[26\] _03587_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ clknet_leaf_1_clk _00791_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07542__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13835_ clknet_leaf_101_clk _00722_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12729__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
X_13766_ clknet_leaf_114_clk _00653_ net1098 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ net226 net1957 net587 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12717_ net237 net1836 net570 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__mux2_1
X_13697_ clknet_leaf_101_clk datapath.multiplication_module.multiplicand_i_n\[14\]
+ net1223 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ net252 net1930 net436 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11929__B1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11869__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12464__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ net2232 net262 net444 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14318_ clknet_leaf_2_clk _01205_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07073__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 datapath.rf.registers\[4\]\[15\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold317 datapath.rf.registers\[26\]\[15\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold328 datapath.rf.registers\[5\]\[15\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 datapath.rf.registers\[24\]\[1\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ clknet_leaf_2_clk _01136_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 _01750_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_4
Xfanout819 _01747_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_4
X_08810_ net680 _03704_ _03736_ _03448_ _03735_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__a221o_1
X_09790_ net1277 _02832_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__or2_1
XANTENNA__07781__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 datapath.rf.registers\[18\]\[20\] vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 datapath.rf.registers\[21\]\[10\] vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net418 _03659_ _03663_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a2bb2o_1
Xhold1028 datapath.rf.registers\[11\]\[4\] vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 datapath.rf.registers\[12\]\[9\] vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
X_08672_ net706 _03598_ net623 vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a21o_1
XANTENNA__07533__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ datapath.rf.registers\[16\]\[15\] net962 net941 datapath.rf.registers\[26\]\[15\]
+ _02549_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12639__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
X_07554_ datapath.rf.registers\[7\]\[16\] net826 net798 datapath.rf.registers\[25\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a22o_1
X_06505_ screen.counter.ct\[7\] vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
XANTENNA__10159__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07485_ datapath.rf.registers\[29\]\[18\] net878 net862 datapath.rf.registers\[28\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1076_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08137__B _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09224_ _03801_ _03802_ net363 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09589__A1 _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09155_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or2_1
XANTENNA__12374__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout501_A _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08106_ datapath.rf.registers\[7\]\[4\] net957 net901 datapath.rf.registers\[20\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a22o_1
XANTENNA__07064__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09086_ net500 net621 net489 net519 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08037_ datapath.rf.registers\[23\]\[6\] net786 net734 datapath.rf.registers\[12\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold840 datapath.rf.registers\[16\]\[26\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 datapath.rf.registers\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 datapath.rf.registers\[21\]\[23\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 datapath.rf.registers\[29\]\[11\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold884 datapath.rf.registers\[9\]\[30\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A _01848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 datapath.rf.registers\[30\]\[22\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ net837 _04498_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__nor2_1
X_08939_ net614 _03842_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11950_ net293 net1899 net578 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ net265 net2542 net594 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__mux2_1
X_11881_ net157 _05866_ net149 screen.controlBus\[0\] vssd1 vssd1 vccd1 vccd1 _00479_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12549__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13620_ clknet_leaf_34_clk _00558_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10832_ _01511_ net710 _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__o21a_1
X_13551_ clknet_leaf_79_clk _00501_ net1233 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10763_ _01501_ net709 _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__o21a_2
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08047__B _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ net2017 net181 net455 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__mux2_1
XANTENNA__10831__B1 _05655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ clknet_leaf_82_clk _00435_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10694_ _01466_ net660 _05542_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_152_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12433_ net2025 net168 net465 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
XANTENNA__12284__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07055__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12364_ net1692 net191 net474 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__mux2_1
X_14103_ clknet_leaf_44_clk _00990_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11315_ net1308 _05696_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12295_ net1731 net193 net482 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__mux2_1
X_14034_ clknet_leaf_33_clk _00921_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11246_ net1789 net142 net134 _02721_ vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ _05826_ screen.screenLogic.currentWrx _05824_ vssd1 vssd1 vccd1 vccd1 _00213_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07763__B1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ _04798_ _04797_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_145_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08307__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ _01429_ _04985_ net1251 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__mux2_1
XANTENNA__07515__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A2 _04277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12459__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13818_ clknet_leaf_51_clk _00705_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10487__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13749_ clknet_leaf_29_clk _00636_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07270_ datapath.rf.registers\[11\]\[23\] net970 net938 datapath.rf.registers\[21\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__a22o_1
XANTENNA__07294__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07046__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold103 net79 vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 net104 vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold125 net101 vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 screen.counter.ct\[20\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12922__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold147 net102 vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 net51 vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ datapath.PC\[26\] net628 _04776_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a21oi_1
Xhold169 net114 vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06554__C_N mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 _05576_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
Xfanout616 _03553_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_2
Xfanout627 _01729_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
X_09842_ _04767_ _04768_ _04676_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__and3b_1
Xfanout638 _03530_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
Xfanout649 _01725_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_2
XANTENNA__07754__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_1
X_06985_ datapath.rf.registers\[25\]\[29\] net798 net772 datapath.rf.registers\[30\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout284_A _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _02148_ _02168_ net681 vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a21o_1
X_08655_ datapath.PC\[19\] _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1193_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ datapath.rf.registers\[11\]\[15\] net775 net760 datapath.rf.registers\[19\]\[15\]
+ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ net337 _03512_ _01717_ _03504_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07537_ datapath.rf.registers\[12\]\[17\] net888 net848 datapath.rf.registers\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout716_A _01783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10813__B1 _05642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ datapath.rf.registers\[28\]\[18\] net720 net715 datapath.rf.registers\[29\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
XANTENNA__07285__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ net498 net495 net513 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07399_ datapath.rf.registers\[8\]\[20\] net927 net918 datapath.rf.registers\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07037__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09138_ _04055_ _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_20_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08314__C _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12832__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ _02656_ net683 net679 _03978_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ net1293 screen.counter.ct\[11\] screen.counter.ct\[10\] screen.counter.ct\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__or4b_1
XANTENNA__07993__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ net321 _06350_ _06351_ net325 net1843 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__a32o_1
Xhold670 datapath.rf.registers\[7\]\[15\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 datapath.rf.registers\[22\]\[23\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 datapath.rf.registers\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _05680_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_9_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06548__A1 mmio.memload_or_instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__C1 _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ net2526 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ net151 _05885_ net126 screen.register.currentXbus\[19\] vssd1 vssd1 vccd1
+ vccd1 _00530_ sky130_fd_sc_hd__a22o_1
XANTENNA__12279__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__A _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11864_ _06253_ datapath.PC\[29\] net305 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__mux2_1
XANTENNA__06720__A1 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ clknet_leaf_97_clk net1393 net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memread2
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ net841 _04446_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11795_ net700 _04787_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13534_ clknet_leaf_80_clk _00484_ net1234 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10746_ net839 _04232_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__nand2_1
XANTENNA__07276__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10280__A1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13465_ clknet_leaf_81_clk _00421_ net1241 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ net842 _03703_ _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_153_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07028__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ net2467 net253 net464 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13396_ clknet_leaf_92_clk net1379 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06577__C_N mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08224__C _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__A1 _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ net2194 net265 net472 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__mux2_1
XANTENNA__12742__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__S net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12278_ net1603 net272 net482 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14017_ clknet_leaf_43_clk _00904_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11229_ net1414 net146 net139 _04898_ vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07736__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06770_ datapath.ru.latched_instruction\[2\] _01595_ _01650_ datapath.ru.latched_instruction\[7\]
+ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a221o_1
XANTENNA__06695__B _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ _02193_ _02212_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08371_ datapath.rf.registers\[10\]\[0\] net919 net875 datapath.rf.registers\[25\]\[0\]
+ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12917__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07322_ datapath.rf.registers\[13\]\[22\] net866 net850 datapath.rf.registers\[1\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XANTENNA__07267__A2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07253_ datapath.rf.registers\[8\]\[23\] net738 net715 datapath.rf.registers\[29\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
X_07184_ datapath.rf.registers\[26\]\[25\] net942 net887 datapath.rf.registers\[9\]\[25\]
+ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07019__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__A1 _03785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12652__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07975__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1039_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_4
X_09825_ _04748_ _04749_ _04718_ _04719_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211o_1
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net459 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
Xfanout468 net471 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_8
Xfanout479 _06452_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ net633 _04682_ net1275 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o21a_1
XANTENNA__10900__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ datapath.rf.registers\[22\]\[30\] net954 net894 datapath.rf.registers\[14\]\[30\]
+ _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a221o_1
X_08707_ net635 _03624_ _03632_ net610 vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a22o_1
X_09687_ _04613_ _04082_ _02886_ _04612_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and4b_1
XANTENNA__08152__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06899_ net1001 net985 net978 net976 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout833_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _03442_ _03551_ net676 _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_120_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08309__C _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12827__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ datapath.ru.latched_instruction\[12\] net1040 net1008 _01626_ _01631_ vssd1
+ vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_25_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ net1420 net517 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[12\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07258__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _05763_ _06044_ _06035_ _05798_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10531_ _05415_ _05439_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__or2_1
XANTENNA__12539__A0 _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13250_ clknet_leaf_65_clk _00240_ net1269 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ _02431_ _02476_ net521 _02566_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_118_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ _05575_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__or3_4
XANTENNA__11211__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ clknet_leaf_32_clk _00173_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12562__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ screen.counter.ct\[4\] screen.counter.ct\[10\] net1287 _05294_ vssd1 vssd1
+ vccd1 vccd1 _05315_ sky130_fd_sc_hd__nor4_1
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07966__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12132_ _06393_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__or2_1
XANTENNA__07430__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12063_ _06335_ _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nand2_1
XANTENNA__07718__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ _05519_ net2261 net585 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
XANTENNA__09183__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_2
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
X_12965_ net300 net2066 net609 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__mux2_1
XANTENNA__08143__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ net151 _05868_ net126 net2639 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__a22o_1
XANTENNA__08694__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ net165 net2431 net551 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ net201 _04835_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__nor2_1
XANTENNA__12737__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ net1336 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__07249__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ net698 _04191_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__B _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13517_ clknet_leaf_66_clk _00467_ net1270 vssd1 vssd1 vccd1 vccd1 datapath.PC\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11450__B1 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10729_ _01488_ net710 _05572_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o22a_2
XFILLER_0_153_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14497_ clknet_leaf_41_clk _01384_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13448_ clknet_leaf_81_clk _00404_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11202__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12472__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13379_ clknet_leaf_89_clk net1471 net1210 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07940_ datapath.rf.registers\[30\]\[8\] net773 net739 datapath.rf.registers\[8\]\[8\]
+ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a221o_1
X_07871_ datapath.rf.registers\[11\]\[9\] net970 net941 datapath.rf.registers\[26\]\[9\]
+ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__a221o_1
XANTENNA__10005__B _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ net635 _04531_ _04533_ _03561_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__o2bb2a_1
X_06822_ net993 _01734_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ net614 _04459_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__or3b_1
X_06753_ datapath.ru.latched_instruction\[20\] _01505_ net1027 vssd1 vssd1 vccd1 vccd1
+ _01680_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_69_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07488__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _03516_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and2_1
X_06684_ _01459_ net1030 net1008 net1041 datapath.ru.latched_instruction\[28\] vssd1
+ vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _01910_ _01952_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12647__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ datapath.rf.registers\[22\]\[0\] net751 _03263_ _03265_ _03270_ vssd1 vssd1
+ vccd1 vccd1 _03281_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_82_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10244__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ _02220_ _02223_ _02224_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__or4_1
X_08285_ datapath.rf.registers\[7\]\[1\] net995 _01739_ vssd1 vssd1 vccd1 vccd1 _03212_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_132_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07236_ datapath.rf.registers\[8\]\[24\] net927 net863 datapath.rf.registers\[28\]\[24\]
+ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12382__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ datapath.rf.registers\[18\]\[25\] net791 net739 datapath.rf.registers\[8\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07948__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09257__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07412__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ datapath.rf.registers\[5\]\[27\] net854 _02020_ _02022_ _02024_ vssd1 vssd1
+ vccd1 vccd1 _02025_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout783_A _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1222 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_2
Xfanout210 _05531_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_1
Xfanout1219 net1221 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_4
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
Xfanout243 _05496_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net256 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout950_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 _05628_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08373__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 _05618_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
Xfanout287 net290 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
X_09808_ _04733_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__nor2_1
Xfanout298 net300 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10180__B1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ net843 net220 net704 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a21o_1
XANTENNA__08125__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ net234 net2197 net566 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__mux2_1
X_11701_ _06142_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__inv_2
X_12681_ net1792 net249 net431 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XANTENNA__12557__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ clknet_leaf_117_clk _01307_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11632_ _06091_ _06092_ _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11432__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ clknet_leaf_5_clk _01238_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11563_ screen.register.currentYbus\[7\] _05737_ _06026_ _06028_ vssd1 vssd1 vccd1
+ vccd1 _06029_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13302_ clknet_leaf_111_clk _00292_ net1103 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10786__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10514_ _05396_ _05408_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__nor2_1
Xwire644 _03201_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_1
XFILLER_0_123_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14282_ clknet_leaf_10_clk _01169_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11494_ screen.register.currentXbus\[19\] _05707_ _05772_ screen.register.currentYbus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07651__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13233_ clknet_leaf_75_clk _00223_ net1250 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
X_10445_ _01799_ net344 net535 net425 vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__and4b_1
XANTENNA__12292__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11801__A2_N net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ clknet_leaf_30_clk _00156_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07403__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ screen.controlBus\[4\] _05291_ _05296_ screen.controlBus\[5\] vssd1 vssd1
+ vccd1 vccd1 _05298_ sky130_fd_sc_hd__or4bb_2
X_12115_ _06373_ _06379_ _06378_ _06377_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__o211ai_2
X_13095_ clknet_leaf_15_clk _00087_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12046_ _06321_ _06322_ _06320_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08364__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07415__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13997_ clknet_leaf_0_clk _00884_ net1070 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08116__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12948_ net237 net1990 net544 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__mux2_1
XANTENNA__08667__A1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12879_ net250 net1753 net549 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
XANTENNA__12467__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14532__1319 vssd1 vssd1 vccd1 vccd1 _14532__1319/HI net1319 sky130_fd_sc_hd__conb_1
XFILLER_0_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07890__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14549_ net1360 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_83_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ datapath.rf.registers\[0\]\[5\] net690 _02982_ _02996_ vssd1 vssd1 vccd1
+ vccd1 _02997_ sky130_fd_sc_hd__o22a_4
XANTENNA__07642__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07021_ _01941_ _01943_ _01945_ _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__or4_1
XFILLER_0_114_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08972_ net337 _03898_ net315 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06633__D_N mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ datapath.rf.registers\[31\]\[8\] net950 net911 datapath.rf.registers\[30\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__a22o_1
Xhold18 screen.counter.ack2 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 datapath.ru.ack_mul_reg vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout197_A _05537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ datapath.rf.registers\[25\]\[10\] net796 _02777_ _02779_ _02780_ vssd1 vssd1
+ vccd1 vccd1 _02781_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06805_ _01638_ net996 _01656_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__and3_1
X_07785_ datapath.rf.registers\[19\]\[11\] net759 net722 datapath.rf.registers\[27\]\[11\]
+ _02711_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a221o_1
XANTENNA__08107__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ _02437_ _03332_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__xnor2_1
X_06736_ datapath.ru.latched_instruction\[16\] net1037 net1004 _01661_ vssd1 vssd1
+ vccd1 vccd1 _01663_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09455_ net653 _04379_ _04381_ net675 vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a31o_1
X_06667_ _01596_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__inv_2
XANTENNA__12377__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_A _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1273_A _00004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08406_ _02437_ _02478_ _03331_ _02433_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o31a_1
XFILLER_0_148_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09386_ _03019_ net684 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nand2_1
X_06598_ _01410_ _01457_ _01478_ _01408_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__o22a_1
XANTENNA__07881__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13368__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ datapath.rf.registers\[26\]\[0\] net988 _01743_ vssd1 vssd1 vccd1 vccd1 _03264_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10768__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07094__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ _03186_ _03189_ _03190_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nor3_1
XANTENNA__07633__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07219_ _02139_ _02141_ _02143_ _02145_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__or4_1
XANTENNA__06841__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__inv_2
X_10230_ net537 _04446_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ net1055 _03576_ _05087_ net700 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a31o_1
XANTENNA__12840__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1005 _01581_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_2
Xfanout1016 _05726_ vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
Xfanout1027 net1031 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
Xfanout1038 net1043 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
X_10092_ net1311 _05018_ _05010_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__o21a_1
X_13920_ clknet_leaf_44_clk _00807_ net1195 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ clknet_leaf_22_clk _00738_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12802_ net291 net2561 net560 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__mux2_1
X_13782_ clknet_leaf_24_clk _00669_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ net299 net2219 net583 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12733_ net180 net2560 net565 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__mux2_1
XANTENNA__12287__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12664_ net169 net2124 net438 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XANTENNA__07872__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14403_ clknet_leaf_104_clk _01290_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11615_ screen.counter.ct\[11\] net1290 net1291 _06077_ vssd1 vssd1 vccd1 vccd1 _06078_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ net1842 net188 net446 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07085__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14334_ clknet_leaf_51_clk _01221_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11546_ screen.register.currentXbus\[6\] _05720_ _05735_ screen.register.currentYbus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07624__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14265_ clknet_leaf_47_clk _01152_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11477_ screen.register.currentYbus\[10\] _05736_ _05737_ screen.register.currentYbus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13216_ clknet_leaf_46_clk _00208_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ net37 net38 vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__or2_1
X_14196_ clknet_leaf_114_clk _01083_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08232__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13147_ clknet_leaf_52_clk _00139_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12750__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10359_ screen.controlBus\[17\] screen.controlBus\[16\] screen.controlBus\[19\] screen.controlBus\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__or4_1
X_13078_ clknet_leaf_26_clk _00070_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_146_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _06305_ _06306_ _06307_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or3_1
XANTENNA__06687__C net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ _02483_ _02484_ _02491_ _02493_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_66_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ net1309 vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__inv_2
X_09240_ net389 _04164_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09171_ net515 net354 _04097_ net386 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_32_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12925__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ datapath.rf.registers\[13\]\[4\] net794 net760 datapath.rf.registers\[19\]\[4\]
+ _03048_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a221o_1
XANTENNA__07076__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07615__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ datapath.rf.registers\[21\]\[5\] net936 net912 datapath.rf.registers\[18\]\[5\]
+ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11250__A1_N net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ _01930_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08040__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1119_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11265__A1_N net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _03877_ _03878_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout481_A _06449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _02831_ _02832_ net647 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold1227_A mmio.memload_or_instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ net393 _03688_ _03520_ net398 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o211a_1
XANTENNA__10686__A1 _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07837_ net515 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout746_A _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ datapath.rf.registers\[16\]\[12\] net960 net956 datapath.rf.registers\[7\]\[12\]
+ _02694_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ _02588_ net519 net684 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06719_ mmio.memload_or_instruction\[21\] net1061 net1006 datapath.ru.latched_instruction\[21\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a32o_4
XFILLER_0_149_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout913_A _01830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ datapath.rf.registers\[14\]\[13\] net799 net734 datapath.rf.registers\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ net370 _04285_ _04286_ _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_149_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07854__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09369_ _02997_ net357 _04260_ net385 vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a211o_1
XANTENNA__12835__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ screen.register.currentYbus\[19\] net130 _05885_ net159 vssd1 vssd1 vccd1
+ vccd1 _00377_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07606__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12380_ net265 net2452 net468 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11331_ mmio.memload_or_instruction\[10\] net1061 net308 net312 datapath.ru.latched_instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14050_ clknet_leaf_43_clk _00937_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11262_ net1560 net142 net135 _02017_ vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13001_ net1542 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__clkbuf_1
X_10213_ net1056 _03578_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__nand2_1
XANTENNA__12570__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ net1544 _05828_ _05836_ vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__a21o_1
XANTENNA__08031__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14531__1318 vssd1 vssd1 vccd1 vccd1 _14531__1318/HI net1318 sky130_fd_sc_hd__conb_1
X_10144_ net536 _04336_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10075_ net539 _04540_ _05001_ net1057 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_128_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ clknet_leaf_6_clk _00790_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13834_ clknet_leaf_15_clk _00721_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06750__C1 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ clknet_leaf_95_clk _00652_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08098__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ net242 net2338 net587 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__mux2_1
X_12716_ net239 net2048 net571 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07845__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13696_ clknet_leaf_101_clk datapath.multiplication_module.multiplicand_i_n\[13\]
+ net1223 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08227__C _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ net253 net2518 net436 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09047__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12745__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11929__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07058__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12578_ net1995 net266 net444 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10601__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14317_ clknet_leaf_1_clk _01204_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11529_ screen.register.currentYbus\[13\] _05776_ _05777_ screen.register.currentYbus\[29\]
+ _05962_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08270__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold307 datapath.rf.registers\[12\]\[30\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 datapath.rf.registers\[22\]\[14\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ clknet_leaf_13_clk _01135_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold329 datapath.rf.registers\[5\]\[16\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08558__A0 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14179_ clknet_leaf_103_clk _01066_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12480__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net812 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07230__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ net411 _03666_ net422 vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a21oi_1
Xhold1007 datapath.rf.registers\[28\]\[23\] vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 datapath.rf.registers\[8\]\[31\] vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 datapath.rf.registers\[28\]\[25\] vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ _03434_ _03595_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08730__A0 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ datapath.rf.registers\[17\]\[15\] net881 net873 datapath.rf.registers\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07553_ _02479_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06504_ screen.register.cFill2 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__inv_2
XANTENNA__07297__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ net651 _02410_ net627 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ net368 _03677_ _03678_ _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12655__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07049__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ net670 _04049_ _04076_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_79_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08105_ _03027_ _03029_ _03030_ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_79_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09085_ net392 _03931_ _03932_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__and3_1
XANTENNA__08261__A2 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1236_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ datapath.rf.registers\[15\]\[6\] net805 net737 datapath.rf.registers\[8\]\[6\]
+ _02960_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold830 datapath.multiplication_module.multiplicand_i\[9\] vssd1 vssd1 vccd1 vccd1
+ net2196 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A0 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold841 datapath.rf.registers\[17\]\[7\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold852 datapath.rf.registers\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 datapath.rf.registers\[9\]\[25\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12390__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 datapath.rf.registers\[23\]\[30\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10903__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold885 keypad.apps.app_c\[1\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 datapath.rf.registers\[8\]\[21\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09265__A _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _03747_ _04497_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout863_A _01851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net635 _03851_ _03863_ net610 vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a22o_1
X_08869_ net413 _03645_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ net269 net2096 net596 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__mux2_1
X_11880_ _05037_ _05258_ _05689_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_123_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ datapath.mulitply_result\[16\] net428 _05655_ _05658_ net662 vssd1 vssd1
+ vccd1 vccd1 _05659_ sky130_fd_sc_hd__a221o_1
XANTENNA__09277__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08328__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ clknet_leaf_79_clk _00500_ net1233 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07288__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ datapath.mulitply_result\[5\] net430 _05597_ _05600_ net659 vssd1 vssd1 vccd1
+ vccd1 _05601_ sky130_fd_sc_hd__a221o_1
XANTENNA__07827__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12501_ _05667_ net577 vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ clknet_leaf_83_clk _00434_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10831__B2 _05658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ datapath.mulitply_result\[26\] net427 net660 vssd1 vssd1 vccd1 vccd1 _05543_
+ sky130_fd_sc_hd__a21o_1
X_12432_ net2260 net173 net466 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08237__C1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12363_ net1950 net194 net473 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14102_ clknet_leaf_24_clk _00989_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11314_ datapath.pc_module.i_ack1 datapath.i_ack vssd1 vssd1 vccd1 vccd1 _05854_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07460__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12294_ net1596 net196 net483 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14033_ clknet_leaf_27_clk _00920_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11245_ net1498 net142 net135 _02783_ vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07212__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _05682_ _05786_ _05794_ net1012 _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a221o_1
X_10127_ net835 _04360_ _05053_ _05052_ net200 vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__o311a_1
XFILLER_0_145_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10058_ _04977_ _04984_ net202 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08519__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13817_ clknet_leaf_47_clk _00704_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09268__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10487__C net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_114_clk _00635_ net1096 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07818__A2 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12475__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ clknet_leaf_110_clk _00614_ net1103 vssd1 vssd1 vccd1 vccd1 columns.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__A2 _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold104 keypad.decode.sticky\[2\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07451__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold115 datapath.rf.registers\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold126 datapath.rf.registers\[25\]\[1\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10008__B net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold137 datapath.rf.registers\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 screen.counter.currentCt\[6\] vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 datapath.multiplication_module.multiplier_i\[4\] vssd1 vssd1 vccd1 vccd1
+ net1525 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _04778_ _04833_ _04835_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 net609 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_4
X_09841_ _01431_ net629 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07203__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_4
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
Xfanout639 _03529_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08951__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ datapath.PC\[14\] net632 _04697_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__nor3_1
X_06984_ datapath.rf.registers\[7\]\[29\] net826 net787 datapath.rf.registers\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
X_08723_ net420 _03646_ _03649_ _03448_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__o211ai_1
XANTENNA__11302__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08654_ net1275 _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ datapath.rf.registers\[21\]\[15\] net746 net715 datapath.rf.registers\[29\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout444_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ datapath.rf.registers\[17\]\[17\] net883 net861 datapath.rf.registers\[28\]\[17\]
+ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a221o_1
XANTENNA__07809__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07467_ datapath.rf.registers\[20\]\[18\] net802 net787 datapath.rf.registers\[23\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a22o_1
XANTENNA__12385__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout709_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09206_ net502 net618 net496 net514 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07690__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ datapath.rf.registers\[11\]\[20\] net971 net871 datapath.rf.registers\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09137_ net338 _04056_ _04063_ _03504_ _01717_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08234__A2 _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ net319 _03607_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08019_ datapath.rf.registers\[7\]\[6\] net956 net920 datapath.rf.registers\[2\]\[6\]
+ _02945_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a221o_1
XANTENNA__06635__A_N mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 datapath.rf.registers\[14\]\[28\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 datapath.rf.registers\[10\]\[9\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ _01440_ _05284_ _05348_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__or3_2
Xhold682 datapath.rf.registers\[16\]\[16\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 datapath.rf.registers\[31\]\[13\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08330__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ net2522 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
X_11932_ net151 _05884_ net126 screen.register.currentXbus\[18\] vssd1 vssd1 vccd1
+ vccd1 _00529_ sky130_fd_sc_hd__a22o_1
XANTENNA__10588__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ net836 _03637_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10814_ net1647 net255 net602 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ clknet_leaf_72_clk datapath.MemWrite net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memwrite
+ sky130_fd_sc_hd__dfrtp_4
X_11794_ net700 _04416_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13533_ clknet_leaf_80_clk _00483_ net1234 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10745_ net1585 net299 net605 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__mux2_1
XANTENNA__12295__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09670__A1 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13464_ clknet_leaf_82_clk _00420_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10280__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ net842 _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12415_ net2286 net257 net464 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13395_ clknet_leaf_109_clk net1391 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12346_ net1774 net269 net473 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
XANTENNA__11780__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ net1734 net275 net481 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09186__B1 _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ clknet_leaf_50_clk _00903_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11228_ net1428 net146 net139 _04909_ vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ _05748_ _05752_ _05805_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__nor3_1
XANTENNA__09489__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__B2 mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__A _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08161__B2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__A _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06711__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08370_ datapath.rf.registers\[16\]\[0\] net961 net885 datapath.rf.registers\[9\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09110__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10256__C1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ datapath.rf.registers\[12\]\[22\] net890 net859 datapath.rf.registers\[15\]\[22\]
+ _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11403__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07252_ datapath.rf.registers\[2\]\[23\] net727 net723 datapath.rf.registers\[27\]\[23\]
+ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a221o_1
XANTENNA__07672__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12933__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07183_ datapath.rf.registers\[13\]\[25\] net866 _02109_ net695 vssd1 vssd1 vccd1
+ vccd1 _02110_ sky130_fd_sc_hd__a211o_1
XANTENNA__10019__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07424__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08431__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 _03514_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_2
Xfanout414 _03453_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_2
XANTENNA__07727__A1 _02653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 net439 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_6
XFILLER_0_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09824_ _04748_ _04749_ _04719_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a21o_1
Xfanout447 _06460_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1101_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_4
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _01679_ _04678_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nor2_1
X_06967_ datapath.rf.registers\[31\]\[30\] net949 net874 datapath.rf.registers\[25\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout561_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A datapath.MemRead vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net637 _03624_ _03620_ net657 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o211a_1
XANTENNA__11287__B2 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ _02792_ _04048_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__or2_1
X_06898_ net1002 net986 net981 _01801_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__and4_2
XFILLER_0_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07063__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _03503_ net616 _03563_ net492 _03352_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout826_A _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ net1003 _03493_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07519_ datapath.rf.registers\[22\]\[17\] net751 net744 datapath.rf.registers\[21\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08455__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09652__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ _03366_ _03425_ _03367_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__o21ai_1
X_10530_ _05439_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__inv_2
XANTENNA__07663__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ _01860_ _01904_ net534 net511 vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or4_1
XANTENNA__08207__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12843__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12200_ _05478_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__o21bai_4
XTAP_TAPCELL_ROW_118_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13180_ clknet_leaf_55_clk _00172_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10392_ net1299 _05307_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11762__A2 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ datapath.mulitply_result\[25\] datapath.multiplication_module.multiplicand_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_131_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12062_ datapath.mulitply_result\[14\] datapath.multiplication_module.multiplicand_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__or2_1
Xhold490 datapath.rf.registers\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ net223 net2491 net584 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
XANTENNA__11514__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11983__A datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout970 _01802_ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_4
XANTENNA__07194__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout981 _01662_ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_2
Xfanout992 _01648_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06796__B net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06941__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__B2 mmio.memload_or_instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ net288 net1705 net609 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__mux2_1
Xhold1190 datapath.rf.registers\[16\]\[27\] vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
X_11915_ net151 _05867_ net126 net2649 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__a22o_1
X_12895_ net168 net1750 net551 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11846_ _06239_ _06240_ net1274 net304 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ net1335 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_11777_ datapath.PC\[5\] net302 _06188_ _06190_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08516__B _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07654__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13516_ clknet_leaf_66_clk _00466_ net1268 vssd1 vssd1 vccd1 vccd1 datapath.PC\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_10728_ datapath.mulitply_result\[31\] net427 net661 vssd1 vssd1 vccd1 vccd1 _05573_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07420__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14496_ clknet_leaf_46_clk _01383_ net1195 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12753__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13447_ clknet_leaf_82_clk _00403_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10659_ net842 _04496_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07406__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13378_ clknet_leaf_92_clk keypad.decode.d1 net1204 vssd1 vssd1 vccd1 vccd1 keypad.decode.d2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ net2095 net199 net479 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07870_ datapath.rf.registers\[18\]\[9\] net914 net862 datapath.rf.registers\[28\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__a22o_1
XANTENNA__07185__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ net996 _01733_ _01741_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__and3_1
X_09540_ net635 _04460_ _04463_ net610 vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a22o_1
X_06752_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nor2_2
XANTENNA__08134__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ net395 _04176_ _04254_ net399 vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a211o_1
X_06683_ datapath.ru.latched_instruction\[27\] net1041 _01609_ vssd1 vssd1 vccd1 vccd1
+ _01611_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_69_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12928__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ _01996_ _02040_ _03346_ _01992_ _01951_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o311a_1
XANTENNA__06696__A1 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__B _03210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08353_ datapath.rf.registers\[5\]\[0\] net783 _03253_ _03255_ _03268_ vssd1 vssd1
+ vccd1 vccd1 _03280_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_22_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout142_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07304_ _02226_ _02228_ _02230_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07330__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07645__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ net651 _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07235_ datapath.rf.registers\[21\]\[24\] net939 net859 datapath.rf.registers\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12663__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1149_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ datapath.rf.registers\[7\]\[25\] net826 net728 datapath.rf.registers\[2\]\[25\]
+ _02087_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07097_ datapath.rf.registers\[30\]\[27\] net911 net898 datapath.rf.registers\[6\]\[27\]
+ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout200 net202 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_4
Xfanout1209 net1212 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 _05531_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
Xfanout222 net225 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
Xfanout233 _05508_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout244 _05496_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10911__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 _05628_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_1
X_09807_ net1278 _03147_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nor2_1
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
Xfanout288 net290 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
X_07999_ datapath.rf.registers\[0\]\[7\] net827 _02921_ _02925_ vssd1 vssd1 vccd1
+ vccd1 _02926_ sky130_fd_sc_hd__o22a_4
X_09738_ net841 net220 net699 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12838__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net418 _04480_ _04595_ net318 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_139_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12209__A0 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ screen.counter.currentCt\[21\] screen.counter.currentCt\[20\] _06138_ vssd1
+ vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__and3_1
X_12680_ net1786 net254 net431 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XANTENNA__08617__A _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ screen.counter.currentCt\[21\] screen.counter.currentCt\[20\] screen.counter.currentCt\[22\]
+ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__or4_1
XANTENNA__09086__C1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11562_ screen.register.currentXbus\[23\] net1015 _05742_ screen.register.currentYbus\[31\]
+ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a221o_1
X_14350_ clknet_leaf_118_clk _01237_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07636__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07100__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ clknet_leaf_112_clk _00291_ net1096 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_10513_ _05399_ net1026 _05422_ _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__or4_1
XFILLER_0_80_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14281_ clknet_leaf_3_clk _01168_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11493_ screen.register.currentXbus\[3\] _05704_ _05775_ screen.register.currentYbus\[19\]
+ _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a221o_1
XANTENNA__12573__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ clknet_leaf_73_clk _00222_ net1245 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10444_ _05352_ _05353_ _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 screen.register.xFill
+ sky130_fd_sc_hd__or4_1
XFILLER_0_150_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08061__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ clknet_leaf_56_clk _00155_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10375_ screen.controlBus\[4\] _05291_ _05296_ screen.controlBus\[5\] vssd1 vssd1
+ vccd1 vccd1 _05297_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _06377_ _06378_ _06379_ _06373_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__a211o_1
X_13094_ clknet_leaf_108_clk _00086_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ datapath.mulitply_result\[11\] datapath.multiplication_module.multiplicand_i\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__and2_1
XANTENNA__10821__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13996_ clknet_leaf_31_clk _00883_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12947_ net238 net1725 net542 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__mux2_1
XANTENNA__12748__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ net255 net2512 net549 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09077__C1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ net704 _03871_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__C net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07627__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ net1359 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_43_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14479_ clknet_leaf_6_clk _01366_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07020_ datapath.rf.registers\[27\]\[29\] net871 net854 datapath.rf.registers\[5\]\[29\]
+ _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14555__1366 vssd1 vssd1 vccd1 vccd1 net1366 _14555__1366/LO sky130_fd_sc_hd__conb_1
XFILLER_0_51_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08052__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08254__A_N net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08971_ _03891_ _03897_ net401 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__mux2_1
X_07922_ _02842_ _02844_ _02846_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__or4_1
Xhold19 screen.register.xFill2 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ datapath.rf.registers\[9\]\[10\] net778 net734 datapath.rf.registers\[12\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a22o_1
XANTENNA__10162__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06905__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ _01646_ _01682_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_2
X_07784_ datapath.rf.registers\[25\]\[11\] net796 net795 datapath.rf.registers\[13\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06735_ datapath.ru.latched_instruction\[16\] net1037 net1004 _01661_ vssd1 vssd1
+ vccd1 vccd1 _01662_ sky130_fd_sc_hd__a22oi_4
X_09523_ _02437_ _03417_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12658__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1099_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ net611 _04375_ _04376_ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06666_ datapath.ru.latched_instruction\[3\] net1042 _01456_ net1009 vssd1 vssd1
+ vccd1 vccd1 _01596_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08405_ _02478_ _03331_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__nor2_1
XANTENNA__10178__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09385_ _03393_ _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06597_ _01406_ _01458_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout524_A _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ datapath.rf.registers\[20\]\[0\] net988 _01734_ vssd1 vssd1 vccd1 vccd1 _03263_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_35_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11798__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ _03192_ _03193_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__or2_1
XANTENNA__12393__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10906__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ datapath.rf.registers\[13\]\[24\] net794 _02144_ _01736_ vssd1 vssd1 vccd1
+ vccd1 _02145_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_115_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ net506 _03120_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout893_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07149_ datapath.rf.registers\[31\]\[26\] net949 net945 datapath.rf.registers\[19\]\[26\]
+ _02075_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a221o_1
XANTENNA__07397__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ datapath.PC\[11\] _03575_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__nand2_1
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_4
Xfanout1017 _05682_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
X_10091_ _05015_ _05017_ net205 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__mux2_1
Xfanout1028 net1031 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_2
Xfanout1039 net1043 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07149__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ clknet_leaf_51_clk _00737_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ net297 net2544 net557 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__mux2_1
XANTENNA__12568__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ net290 datapath.rf.registers\[30\]\[1\] net583 vssd1 vssd1 vccd1 vccd1 _00180_
+ sky130_fd_sc_hd__mux2_1
X_13781_ clknet_leaf_28_clk _00668_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12732_ net630 _05575_ _06443_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__or3_4
XFILLER_0_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ net171 net2461 net438 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
X_14402_ clknet_leaf_33_clk _01289_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07609__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11614_ screen.counter.ct\[10\] _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ net1686 net192 net445 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ clknet_leaf_32_clk _01220_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11545_ net1011 _06011_ _06006_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14264_ clknet_leaf_39_clk _01151_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11476_ screen.register.currentXbus\[26\] net1013 _05946_ vssd1 vssd1 vccd1 vccd1
+ _05947_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ clknet_leaf_39_clk _00207_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10427_ net37 net38 vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__nor2_1
XANTENNA__08034__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ clknet_leaf_50_clk _01082_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07388__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ screen.controlBus\[21\] screen.controlBus\[20\] screen.controlBus\[23\] screen.controlBus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__or4_1
X_13146_ clknet_leaf_51_clk _00138_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06596__B1 _01492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ clknet_leaf_29_clk _00069_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10289_ net391 _04296_ _04297_ net399 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _06305_ _06306_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07560__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12478__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ clknet_leaf_22_clk _00866_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06520_ net34 net39 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07312__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ net499 net620 net488 net514 vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_32_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08121_ datapath.rf.registers\[14\]\[4\] net801 net750 datapath.rf.registers\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08273__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11411__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ datapath.rf.registers\[3\]\[5\] net964 net880 datapath.rf.registers\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07003_ net648 net535 net626 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12941__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07379__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08720__A _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08954_ _02478_ net681 _03880_ _03449_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__o22a_1
X_07905_ _01616_ _01727_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__nor2_1
XANTENNA__10135__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ net393 _03688_ _03520_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout474_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ datapath.rf.registers\[0\]\[10\] _02762_ net690 vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__mux2_4
XANTENNA__10686__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ datapath.rf.registers\[14\]\[12\] net892 net888 datapath.rf.registers\[12\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout641_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ net419 _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07839__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06718_ mmio.memload_or_instruction\[21\] net1061 net1006 datapath.ru.latched_instruction\[21\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a32oi_4
X_07698_ _02620_ _02622_ _02624_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07303__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06649_ datapath.ru.n_memwrite2 _01578_ net1042 datapath.ru.zero_multi1 vssd1 vssd1
+ vccd1 vccd1 _01579_ sky130_fd_sc_hd__a211o_1
X_09437_ _04027_ _04028_ net373 vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ net402 _04018_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08264__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ net649 _03244_ _03211_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_113_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10636__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09299_ _03127_ _03312_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ _01514_ net1027 net308 net312 datapath.ru.latched_instruction\[9\] vssd1
+ vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__a32o_1
XANTENNA__08333__C _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08016__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ net1519 net142 net134 _02059_ vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12851__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ datapath.PC\[14\] _03577_ datapath.PC\[15\] vssd1 vssd1 vccd1 vccd1 _05139_
+ sky130_fd_sc_hd__o21a_1
X_13000_ net2008 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__clkbuf_1
X_11192_ mmio.key_data\[5\] net220 _05829_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__and3_1
X_10143_ _04310_ _04336_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or2_1
XANTENNA__08319__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09516__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07790__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ datapath.PC\[26\] net539 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ clknet_leaf_117_clk _00789_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07542__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ clknet_leaf_3_clk _00720_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12298__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ clknet_leaf_14_clk _00651_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10976_ net235 net2502 net586 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__mux2_1
X_14554__1365 vssd1 vssd1 vccd1 vccd1 net1365 _14554__1365/LO sky130_fd_sc_hd__conb_1
XFILLER_0_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12715_ net246 net2567 net571 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__mux2_1
X_13695_ clknet_leaf_101_clk datapath.multiplication_module.multiplicand_i_n\[12\]
+ net1223 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12646_ net257 net1977 net436 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12577_ net2405 net271 net445 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ clknet_leaf_30_clk _01203_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11528_ _05303_ _05784_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 datapath.rf.registers\[20\]\[1\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08007__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold319 datapath.multiplication_module.multiplicand_i\[8\] vssd1 vssd1 vccd1 vccd1
+ net1685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12761__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14247_ clknet_leaf_18_clk _01134_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11459_ _05303_ _05782_ net975 vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09074__A2_N _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08558__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ clknet_leaf_43_clk _01065_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11562__B1 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ clknet_leaf_2_clk _00121_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07781__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09507__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 datapath.rf.registers\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 datapath.rf.registers\[9\]\[13\] vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _03348_ _03596_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07533__A2 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ datapath.rf.registers\[31\]\[15\] net949 net889 datapath.rf.registers\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ _02457_ net522 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__and2_1
X_06503_ screen.register.xFill2 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07483_ datapath.rf.registers\[0\]\[18\] _02409_ net828 vssd1 vssd1 vccd1 vccd1 _02410_
+ sky130_fd_sc_hd__mux2_8
XANTENNA__12936__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ net362 _03672_ _03673_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09153_ _04074_ _04077_ _04079_ net613 net670 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08246__B1 _01777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08104_ datapath.rf.registers\[11\]\[4\] net970 net934 datapath.rf.registers\[23\]\[4\]
+ _03024_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__a221o_1
XANTENNA__08434__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09084_ net688 _04008_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ datapath.rf.registers\[6\]\[6\] net813 net809 datapath.rf.registers\[4\]\[6\]
+ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12671__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold820 datapath.rf.registers\[9\]\[21\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 datapath.rf.registers\[17\]\[17\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 datapath.rf.registers\[30\]\[6\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 datapath.rf.registers\[30\]\[2\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 columns.count\[1\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A _05673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 datapath.rf.registers\[27\]\[18\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold886 datapath.rf.registers\[24\]\[23\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold897 datapath.rf.registers\[17\]\[21\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__S net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ net1052 _04912_ _04911_ net837 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o211a_1
X_08937_ net653 _03842_ _03852_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout856_A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ net410 _03647_ net414 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07524__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ datapath.rf.registers\[22\]\[10\] net952 net884 datapath.rf.registers\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a22o_1
X_08799_ net501 net622 net490 net528 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__o211a_1
X_10830_ net841 _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08328__C _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10761_ net840 _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__or2_1
XANTENNA__12846__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ net163 net2279 net457 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__mux2_1
X_13480_ clknet_leaf_83_clk _00433_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10831__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10692_ net843 _04540_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13352__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08237__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12431_ net2000 net184 net465 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10044__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ net1689 net199 net474 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__mux2_1
XANTENNA__10595__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14101_ clknet_leaf_28_clk _00988_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11313_ datapath.ru.n_memwrite datapath.MemWrite net659 datapath.ru.n_memread vssd1
+ vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a22o_1
XANTENNA__12581__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ net1669 net210 net483 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__mux2_1
X_11244_ net1480 net142 net135 _02831_ vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__a22o_1
X_14032_ clknet_leaf_4_clk _00919_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net975 _05822_ _05300_ _05769_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10126_ _04338_ _04359_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nor2_1
XANTENNA__07763__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _04981_ _04983_ net702 vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__mux2_1
XANTENNA__08465__A_N net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07515__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13816_ clknet_leaf_40_clk _00703_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09268__A2 _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13747_ clknet_leaf_59_clk _00634_ net1267 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10959_ net181 net2198 net586 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12756__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ clknet_leaf_110_clk _00613_ net1103 vssd1 vssd1 vccd1 vccd1 columns.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11264__A1_N net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12629_ net1618 net184 net441 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__mux2_1
XANTENNA__08254__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10035__B1 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__A1 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold105 keypad.decode.sticky_n\[1\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold116 screen.controlBus\[26\] vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 keypad.apps.button\[0\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 datapath.rf.registers\[0\]\[8\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 net103 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09366__A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _04680_ _04766_ _04681_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__o21ai_2
Xfanout607 net609 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout618 _03531_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_4
Xfanout629 _01728_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10305__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07754__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ net632 _04697_ datapath.PC\[14\] vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__o21a_1
X_06983_ _01907_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__and2_2
XANTENNA__06962__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ net420 _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand2_1
X_08653_ datapath.PC\[17\] _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08429__B _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07604_ datapath.rf.registers\[31\]\[15\] net818 net810 datapath.rf.registers\[4\]\[15\]
+ _02527_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _01860_ net622 vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_105_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09113__D1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07535_ datapath.rf.registers\[29\]\[17\] net876 _02461_ net696 vssd1 vssd1 vccd1
+ vccd1 _02462_ sky130_fd_sc_hd__a211o_1
XFILLER_0_147_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout437_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ datapath.rf.registers\[14\]\[18\] net800 net775 datapath.rf.registers\[11\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09205_ _04129_ _04131_ net373 vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07397_ net648 net525 net626 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10026__B1 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ net400 _03858_ _03859_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__a31oi_2
XANTENNA__10577__A1 _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07442__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ net401 _03762_ _03993_ net336 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__o211a_1
XANTENNA__10914__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08018_ datapath.rf.registers\[18\]\[6\] net912 net868 datapath.rf.registers\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a22o_1
XANTENNA__07993__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold650 datapath.rf.registers\[10\]\[20\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 datapath.rf.registers\[26\]\[8\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09707__C _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14553__1364 vssd1 vssd1 vccd1 vccd1 net1364 _14553__1364/LO sky130_fd_sc_hd__conb_1
Xhold672 datapath.rf.registers\[21\]\[8\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 datapath.rf.registers\[19\]\[20\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 datapath.rf.registers\[31\]\[6\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07745__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _04841_ _04848_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__xor2_1
XANTENNA__06953__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ net236 net2040 net606 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__mux2_1
X_11931_ net151 _05883_ net126 screen.register.currentXbus\[17\] vssd1 vssd1 vccd1
+ vccd1 _00528_ sky130_fd_sc_hd__a22o_1
XANTENNA__08170__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07243__B net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11862_ net207 _04854_ _06251_ net705 vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__a211o_1
X_13601_ clknet_leaf_79_clk net1399 net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memwrite2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _01516_ net658 _05642_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12576__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ _06202_ net1650 net302 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ clknet_leaf_86_clk _00482_ net1231 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10744_ _01478_ net709 _05584_ _05585_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_41_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13463_ clknet_leaf_77_clk _00419_ net1249 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10280__A3 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ net1274 _05520_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12414_ net1822 net263 net464 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13394_ clknet_leaf_92_clk net1370 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12345_ net1727 net275 net475 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07984__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ net1632 net279 net480 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__mux2_1
XANTENNA__09186__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09186__B2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14015_ clknet_leaf_37_clk _00902_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11227_ net1419 net145 net139 _05009_ vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__a22o_1
XANTENNA__07736__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__inv_2
XANTENNA__10740__A1 _01464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06944__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ datapath.PC\[31\] net1313 _04867_ _04878_ _04898_ vssd1 vssd1 vccd1 vccd1
+ _05036_ sky130_fd_sc_hd__a2111o_2
X_11089_ _05678_ _05705_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08249__B _03175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12486__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07320_ datapath.rf.registers\[30\]\[22\] net911 net894 datapath.rf.registers\[14\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07251_ datapath.rf.registers\[13\]\[23\] net793 net749 datapath.rf.registers\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11403__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07182_ datapath.rf.registers\[7\]\[25\] net958 net946 datapath.rf.registers\[19\]\[25\]
+ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07975__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout404 net407 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07188__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 net417 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_2
Xfanout426 net430 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09823_ _04719_ _04749_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__nand2b_1
Xfanout437 net439 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_4
Xfanout448 net451 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_8
Xfanout459 _06457_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
XANTENNA__10192__C1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ datapath.PC\[19\] net633 _04679_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_107_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06966_ datapath.rf.registers\[21\]\[30\] net938 net881 datapath.rf.registers\[17\]\[30\]
+ _01892_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a221o_1
X_08705_ net335 _03631_ net316 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_61_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09685_ _02614_ _02702_ _03947_ _03978_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__and4_1
X_06897_ net986 net978 _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08152__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _03548_ net636 net610 _03550_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07360__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout721_A _01782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net1003 _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__nor2_4
XANTENNA__10909__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout819_A _01747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ datapath.rf.registers\[5\]\[17\] net782 net740 datapath.rf.registers\[1\]\[17\]
+ _02444_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08498_ _02259_ _03422_ _03423_ _02257_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o31a_1
XFILLER_0_147_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07449_ datapath.rf.registers\[24\]\[19\] net905 _02375_ net694 vssd1 vssd1 vccd1
+ vccd1 _02376_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _02763_ _02812_ _02855_ _02905_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_70_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ net675 _04008_ _04041_ _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_150_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10391_ _05309_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nand2_1
XANTENNA__11211__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12130_ datapath.mulitply_result\[25\] datapath.multiplication_module.multiplicand_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__and2_1
XANTENNA__08341__C _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__D_N net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ datapath.mulitply_result\[14\] datapath.multiplication_module.multiplicand_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_131_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 datapath.rf.registers\[7\]\[26\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 datapath.mulitply_result\[19\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ net233 net2549 net585 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
XANTENNA__11983__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 _01806_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_8
Xfanout971 _01802_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 _01657_ vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_51_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ net180 net2572 net609 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_84_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 datapath.rf.registers\[23\]\[26\] vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08143__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1191 datapath.rf.registers\[11\]\[26\] vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ net155 _05866_ _06265_ net2509 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12894_ net171 net2365 net552 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
X_11845_ net704 _03703_ net208 _04780_ net304 vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ net1334 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ _05599_ net175 _06189_ net177 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07103__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13515_ clknet_leaf_66_clk _00465_ net1270 vssd1 vssd1 vccd1 vccd1 datapath.PC\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_10727_ net845 _05571_ _05570_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_109_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14495_ clknet_leaf_38_clk _01382_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11450__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13446_ clknet_leaf_82_clk _00402_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10658_ net222 net2294 net607 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13377_ clknet_leaf_91_clk net1396 net1204 vssd1 vssd1 vccd1 vccd1 keypad.decode.q2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10589_ datapath.multiplication_module.multiplicand_i\[0\] _03207_ net349 vssd1 vssd1
+ vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[1\] sky130_fd_sc_hd__mux2_1
XFILLER_0_140_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ net1557 net211 net479 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
XANTENNA__09159__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12259_ net211 net2346 net486 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__mux2_1
XANTENNA__07709__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_118_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11910__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ net990 _01746_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__and2_2
XANTENNA__07590__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06751_ datapath.ru.latched_instruction\[18\] net1037 vssd1 vssd1 vccd1 vccd1 _01678_
+ sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_75_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08134__A2 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06682_ net1041 _01609_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__nor2_1
X_09470_ _02793_ net679 _04394_ _04396_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_69_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08421_ _01996_ _02040_ _03346_ _01992_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14552__1363 vssd1 vssd1 vccd1 vccd1 net1363 _14552__1363/LO sky130_fd_sc_hd__conb_1
X_08352_ _03274_ _03275_ _03277_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__or4bb_1
XPHY_EDGE_ROW_127_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ datapath.rf.registers\[3\]\[22\] net768 net742 datapath.rf.registers\[1\]\[22\]
+ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12944__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ _03208_ _03209_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__or2_1
XANTENNA__08842__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ _02154_ _02156_ _02158_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ datapath.rf.registers\[4\]\[25\] net811 net742 datapath.rf.registers\[1\]\[25\]
+ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout302_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ datapath.rf.registers\[11\]\[27\] net971 net934 datapath.rf.registers\[23\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout212 _05531_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_1
Xfanout223 net225 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xfanout234 _05665_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout671_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06908__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 _05644_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_1
Xfanout267 _05628_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08373__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ net1278 _03147_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 _05613_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
X_07998_ _02917_ _02918_ _02923_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__or4_1
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07581__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ net843 net220 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__nand2_4
X_06949_ datapath.rf.registers\[31\]\[30\] net818 net760 datapath.rf.registers\[19\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout936_A _01817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08125__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
X_09668_ _03453_ _04527_ _04592_ _04594_ net422 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a221o_1
X_08619_ _01860_ net360 vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nand2_1
XANTENNA__10639__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ _02079_ net531 net405 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
X_11630_ screen.counter.currentCt\[17\] screen.counter.currentCt\[16\] screen.counter.currentCt\[19\]
+ screen.counter.currentCt\[18\] vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__or4_1
XANTENNA__08336__C _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11561_ screen.register.currentXbus\[15\] net1016 _05736_ screen.register.currentYbus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12854__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13300_ clknet_leaf_91_clk _00290_ net1209 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10512_ _05414_ net1025 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14280_ clknet_leaf_14_clk _01167_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11492_ _05773_ _05780_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ clknet_leaf_76_clk _00221_ net1248 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
X_10443_ _05350_ _05351_ _05354_ _05355_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07939__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ clknet_leaf_3_clk _00154_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ _05278_ _05285_ _05292_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nor3_1
X_12113_ _06372_ _06374_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nor2_1
X_13093_ clknet_leaf_108_clk _00085_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12044_ datapath.mulitply_result\[11\] datapath.multiplication_module.multiplicand_i\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08364__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout790 net792 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
X_13995_ clknet_leaf_56_clk _00882_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_57_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08116__A2 _01747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12946_ net245 net2237 net543 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12877_ net260 net1690 net549 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
XANTENNA__11234__A datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11828_ net1275 net303 _06228_ _04966_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ net1358 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_64_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11759_ datapath.ru.n_memwrite2 datapath.ru.n_memread2 _01601_ _05856_ vssd1 vssd1
+ vccd1 vccd1 _06176_ sky130_fd_sc_hd__o31a_1
XANTENNA__12764__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09639__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14478_ clknet_leaf_1_clk _01365_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13429_ clknet_leaf_88_clk _00385_ net1216 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08970_ _03761_ _03896_ net394 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07921_ datapath.rf.registers\[3\]\[8\] net967 net943 datapath.rf.registers\[26\]\[8\]
+ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__a221o_1
XANTENNA__08355__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ datapath.rf.registers\[31\]\[10\] net817 net759 datapath.rf.registers\[19\]\[10\]
+ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a221o_1
XANTENNA__07563__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ _01614_ net651 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__or2_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
X_07783_ datapath.rf.registers\[20\]\[11\] net804 net734 datapath.rf.registers\[12\]\[11\]
+ _02709_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a221o_1
XANTENNA__12939__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08107__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _03977_ _04420_ _04446_ _03946_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__and4b_1
XFILLER_0_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06734_ datapath.ru.latched_instruction\[16\] _01511_ net1028 vssd1 vssd1 vccd1 vccd1
+ _01661_ sky130_fd_sc_hd__mux2_1
XANTENNA__07315__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08574__A2_N net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ net636 _04367_ _04375_ net613 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a31o_1
X_06665_ datapath.ru.latched_instruction\[2\] net1042 _01478_ net1009 vssd1 vssd1
+ vccd1 vccd1 _01595_ sky130_fd_sc_hd__a22oi_4
XANTENNA_fanout252_A _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ _02526_ _02568_ _03328_ _02521_ _02480_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__o311a_1
X_09384_ _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand2_1
X_06596_ datapath.ru.latched_instruction\[11\] _01519_ _01492_ datapath.ru.latched_instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08335_ datapath.rf.registers\[19\]\[0\] _01738_ net972 vssd1 vssd1 vccd1 vccd1 _03262_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12674__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout517_A _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1259_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ datapath.rf.registers\[24\]\[1\] net907 net883 datapath.rf.registers\[17\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a22o_1
XANTENNA__07094__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07217_ datapath.rf.registers\[31\]\[24\] net819 net764 datapath.rf.registers\[17\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06841__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ net506 _03120_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07148_ datapath.rf.registers\[14\]\[26\] net893 net878 datapath.rf.registers\[29\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout886_A _01841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ datapath.rf.registers\[2\]\[27\] net728 net723 datapath.rf.registers\[27\]\[27\]
+ _02003_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a221o_1
XANTENNA__10922__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1007 _01581_ vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
X_10090_ _04822_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__nor2_1
XANTENNA__10138__C1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1029 net1031 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07554__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_12800_ net288 net1586 net560 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_153_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13780_ clknet_leaf_117_clk _00667_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ net183 net1655 net583 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__mux2_1
XANTENNA__08628__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12731_ net166 net2580 net571 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12662_ net185 net2026 net437 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ clknet_leaf_40_clk _01288_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11613_ screen.counter.ct\[9\] net1293 _06075_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__and3_1
XANTENNA__12584__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ net1776 net197 net446 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332_ clknet_leaf_53_clk _01219_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11544_ screen.register.currentXbus\[14\] _05709_ _06008_ _06010_ vssd1 vssd1 vccd1
+ vccd1 _06011_ sky130_fd_sc_hd__a211o_1
XANTENNA__09459__A _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07085__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14263_ clknet_leaf_45_clk _01150_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11475_ screen.register.currentXbus\[2\] _05720_ _05735_ screen.register.currentYbus\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13214_ clknet_leaf_50_clk _00206_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ net35 net36 vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__or2_1
X_14194_ clknet_leaf_33_clk _01081_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13145_ clknet_leaf_47_clk _00137_ net1197 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10357_ _05275_ _05276_ _05277_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__or4_1
X_13076_ clknet_leaf_105_clk _00068_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14551__1362 vssd1 vssd1 vccd1 vccd1 net1362 _14551__1362/LO sky130_fd_sc_hd__conb_1
X_10288_ _04259_ _05214_ net388 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__mux2_1
X_12027_ _06301_ _06303_ _06300_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11341__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12759__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ clknet_leaf_51_clk _00865_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12929_ net2305 net165 net546 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12494__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08120_ datapath.rf.registers\[4\]\[4\] net812 net777 datapath.rf.registers\[11\]\[4\]
+ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a221o_1
XANTENNA__07076__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__B1 _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11411__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ _02974_ _02975_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__and2_2
XFILLER_0_153_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07002_ datapath.rf.registers\[0\]\[29\] net829 _01919_ _01928_ vssd1 vssd1 vccd1
+ vccd1 _01929_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06557__C_N mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07617__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ net415 _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nand2_1
XANTENNA__06521__A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07904_ datapath.rf.registers\[0\]\[9\] _02830_ net828 vssd1 vssd1 vccd1 vccd1 _02831_
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_138_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ net639 _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nand2_1
XANTENNA__07536__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ _02751_ _02755_ _02756_ _02761_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__or4_1
XANTENNA__07000__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12669__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A2 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ datapath.rf.registers\[31\]\[12\] net948 net912 datapath.rf.registers\[18\]\[12\]
+ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a221o_1
X_09505_ net415 _04123_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ _01643_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__inv_2
XANTENNA__10189__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ datapath.rf.registers\[11\]\[13\] net774 net730 datapath.rf.registers\[16\]\[13\]
+ _02623_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout634_A _03560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ _04361_ _04362_ net688 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
X_06648_ datapath.pc_module.i_ack1 datapath.pc_module.i_ack2 vssd1 vssd1 vccd1 vccd1
+ _01578_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09367_ net641 _04279_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout801_A _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ mmio.memload_or_instruction\[12\] net1061 vssd1 vssd1 vccd1 vccd1 _01509_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10917__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ net646 _03210_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09298_ _04210_ _04224_ net616 _04197_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08249_ _03148_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ net424 _05844_ net140 net1454 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a2bb2o_1
X_10211_ datapath.PC\[15\] _03977_ net537 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11191_ _05834_ _05835_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10142_ _05065_ _05068_ datapath.PC\[6\] net1243 vssd1 vssd1 vccd1 vccd1 _05069_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08319__A2 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _04934_ _04999_ _04541_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07527__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ clknet_leaf_119_clk _00788_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12579__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_15_clk _00719_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13763_ clknet_leaf_105_clk _00650_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10975_ net238 net2020 net588 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ net250 net2412 net569 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__mux2_1
XANTENNA__10295__D1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ clknet_leaf_100_clk datapath.multiplication_module.multiplicand_i_n\[11\]
+ net1223 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12645_ net264 net1920 net436 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07058__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ net2021 net275 net446 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14315_ clknet_leaf_17_clk _01202_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11527_ _05745_ _05993_ _05680_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14246_ clknet_leaf_105_clk _01133_ net1101 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold309 datapath.rf.registers\[24\]\[8\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ _05303_ _05712_ _05898_ _05306_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_123_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _05048_ _05179_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14177_ clknet_leaf_43_clk _01064_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11389_ _02587_ net669 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__and2_1
XANTENNA__07766__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ clknet_leaf_13_clk _00120_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07230__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ clknet_leaf_105_clk _00051_ net1101 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 datapath.rf.registers\[28\]\[24\] vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07518__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12489__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _02546_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__inv_2
XANTENNA__06741__A1 mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14087__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ _02457_ net522 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06502_ net1 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__inv_2
XANTENNA__10825__B1 _05652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07482_ _02403_ _02406_ _02407_ _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__or4_1
XANTENNA__07297__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09221_ net380 _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07049__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ net612 _04065_ _04078_ _04055_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__o22a_1
X_08103_ datapath.rf.registers\[4\]\[4\] net928 net856 datapath.rf.registers\[15\]\[4\]
+ _03021_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11250__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12952__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _03323_ _04009_ net641 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_79_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout215_A _05526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ datapath.rf.registers\[14\]\[6\] net799 net774 datapath.rf.registers\[11\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a22o_1
Xhold810 datapath.rf.registers\[29\]\[10\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold821 datapath.rf.registers\[23\]\[25\] vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 datapath.rf.registers\[29\]\[0\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 datapath.rf.registers\[15\]\[7\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 datapath.mulitply_result\[23\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07757__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 datapath.rf.registers\[21\]\[26\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 datapath.rf.registers\[6\]\[6\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold887 datapath.rf.registers\[5\]\[3\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 datapath.rf.registers\[20\]\[4\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07221__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ datapath.PC\[23\] _03585_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout584_A _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ net315 _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__or2_1
XANTENNA__09562__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _02345_ net685 net678 _02349_ _03793_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__o221a_1
XANTENNA__12399__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ datapath.rf.registers\[21\]\[10\] net936 net880 datapath.rf.registers\[17\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
X_08798_ net501 net622 net490 net531 vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07749_ datapath.rf.registers\[2\]\[12\] net726 _02663_ _02672_ _02675_ vssd1 vssd1
+ vccd1 vccd1 _02676_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_123_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10760_ _05483_ _05598_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nor2_1
XANTENNA__07288__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09419_ net381 _03965_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__or2_1
X_10691_ net843 _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__nor2_1
X_14550__1361 vssd1 vssd1 vccd1 vccd1 net1361 _14550__1361/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_43_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12430_ net2056 net190 net466 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XANTENNA__13739__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08344__C _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net1612 net211 net474 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12862__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14100_ clknet_leaf_115_clk _00987_ net1075 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11792__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ _01636_ datapath.ack_mul vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07460__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12292_ net2064 net215 net482 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ clknet_leaf_5_clk _00918_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ net1515 net141 net136 _02876_ vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _05785_ _05796_ _05798_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a211o_1
XANTENNA__07212__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ net1055 _05049_ _05051_ net835 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__o211ai_1
X_10056_ _04449_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__nor2_1
XANTENNA__07920__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ clknet_leaf_45_clk _00702_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13746_ clknet_leaf_33_clk _00633_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10958_ net630 _05575_ _05671_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__or3_1
X_13677_ clknet_leaf_110_clk _00612_ net1106 vssd1 vssd1 vccd1 vccd1 columns.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ _01651_ _01669_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__nand2_2
XFILLER_0_143_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12628_ net2167 net189 net442 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11232__B1 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ net211 net1634 net450 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__mux2_1
XANTENNA__07987__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold106 datapath.rf.registers\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07451__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 screen.controlBus\[8\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 net62 vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 datapath.rf.registers\[13\]\[0\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ clknet_leaf_28_clk _01116_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07739__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_4
XANTENNA__07203__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10305__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 _03531_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _01624_ _04678_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__nor2_1
XANTENNA__08951__A2 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06982_ _01885_ _01905_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ net413 net410 _03647_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__or3_1
XANTENNA__11299__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1190 net1198 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_4
X_08652_ datapath.PC\[16\] _03578_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__or2_1
XANTENNA__10321__A _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06714__A1 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07911__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ datapath.rf.registers\[8\]\[15\] net739 net731 datapath.rf.registers\[16\]\[15\]
+ _02529_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a221o_1
X_08583_ net997 _03062_ _03507_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12947__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07534_ datapath.rf.registers\[23\]\[17\] net935 net885 datapath.rf.registers\[9\]\[17\]
+ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07465_ datapath.rf.registers\[15\]\[18\] net806 net727 datapath.rf.registers\[2\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a22o_1
XANTENNA__08445__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09204_ net366 _04023_ _04024_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07690__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ datapath.rf.registers\[0\]\[20\] net829 _02313_ _02322_ vssd1 vssd1 vccd1
+ vccd1 _02323_ sky130_fd_sc_hd__o22ai_2
XANTENNA__08164__C _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ net401 _04060_ _04061_ net340 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__a31o_1
XANTENNA__12682__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ net401 _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__nand2_1
XANTENNA__07442__A2 _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ _02936_ _02941_ _02942_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout799_A _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 datapath.rf.registers\[29\]\[8\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold651 datapath.rf.registers\[10\]\[0\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 datapath.rf.registers\[21\]\[28\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold673 datapath.rf.registers\[17\]\[5\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 datapath.rf.registers\[8\]\[18\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 datapath.rf.registers\[2\]\[16\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _04879_ _04894_ _04893_ net206 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a211o_1
X_08919_ net363 _03768_ _03769_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _04823_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08155__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ net151 _05882_ net126 screen.register.currentXbus\[16\] vssd1 vssd1 vccd1
+ vccd1 _00527_ sky130_fd_sc_hd__a22o_1
XANTENNA__07902__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08339__C _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ net206 _05558_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nor2_1
XANTENNA__12857__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ clknet_leaf_97_clk datapath.ack_mul net1221 vssd1 vssd1 vccd1 vccd1 datapath.ru.ack_mul_reg
+ sky130_fd_sc_hd__dfrtp_1
X_10812_ datapath.mulitply_result\[13\] net428 net658 vssd1 vssd1 vccd1 vccd1 _05643_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ net833 _06200_ _06201_ _05149_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__a31o_1
X_13531_ clknet_leaf_86_clk _00481_ net1231 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10265__A1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10743_ datapath.mulitply_result\[2\] net426 net659 vssd1 vssd1 vccd1 vccd1 _05585_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_41_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13462_ clknet_leaf_77_clk _00418_ net1249 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07681__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ net213 net2252 net607 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__mux2_1
X_12413_ net1771 net267 net464 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
XANTENNA__11214__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09958__A1 _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13393_ clknet_leaf_109_clk net1389 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12592__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07969__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12344_ net1582 net278 net472 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__mux2_1
XANTENNA__07433__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12275_ net2290 net281 net480 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__mux2_1
XANTENNA__11517__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ clknet_leaf_50_clk _00901_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11226_ net1520 net145 net139 _04943_ vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__a22o_1
XANTENNA__09186__A2 _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ _05711_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__or2_1
XANTENNA__10840__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10740__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _04888_ _04932_ _05032_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__or4_2
X_11088_ _05720_ _05735_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__or4_1
XANTENNA__08146__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ net701 _04471_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__nand2_1
XANTENNA__12767__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10256__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09110__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13729_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[14\] net1206
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07250_ datapath.rf.registers\[18\]\[23\] net790 net752 datapath.rf.registers\[22\]\[23\]
+ _02174_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07672__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11205__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ datapath.rf.registers\[10\]\[25\] net918 net879 datapath.rf.registers\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07424__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout405 net407 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_4
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09822_ datapath.PC\[8\] _02877_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__or2_1
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_2
XANTENNA__10750__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_4
Xfanout449 net451 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_8
X_09753_ net633 _04679_ datapath.PC\[19\] vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o21a_1
X_06965_ datapath.rf.registers\[2\]\[30\] net921 net858 datapath.rf.registers\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout282_A _05607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ net398 _03630_ _03516_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__o21ai_1
X_09684_ _03570_ _03594_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06896_ net984 net981 _01676_ net1002 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__o211a_1
X_08635_ _03504_ _03560_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12677__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _01627_ _01631_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__or2_2
XANTENNA__09637__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07517_ datapath.rf.registers\[20\]\[17\] net804 net795 datapath.rf.registers\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08497_ _03422_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07448_ datapath.rf.registers\[18\]\[19\] net914 net849 datapath.rf.registers\[1\]\[19\]
+ _02374_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a221o_1
XANTENNA__07663__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07379_ datapath.rf.registers\[3\]\[20\] net768 net732 datapath.rf.registers\[16\]\[20\]
+ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09118_ net672 _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ net1290 _05310_ _05311_ net1295 vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__or4b_1
XANTENNA__08612__A1 _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06704__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09049_ _03969_ _03974_ _03975_ net677 vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09119__A1_N net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ net321 _06333_ _06334_ net325 net1785 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold470 datapath.rf.registers\[16\]\[17\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 datapath.rf.registers\[19\]\[12\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__B1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 datapath.mulitply_result\[15\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net227 net1795 net582 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XANTENNA__14119__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net951 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_4
Xfanout961 _01806_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__buf_2
XANTENNA__11263__A1_N net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout972 _01758_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_2
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08128__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout994 net997 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_51_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ net165 net2357 net542 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__mux2_1
Xhold1170 screen.register.currentYbus\[5\] vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _05247_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__nor2_2
Xhold1181 datapath.rf.registers\[24\]\[31\] vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 datapath.rf.registers\[6\]\[5\] vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12587__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ net187 net2028 net551 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11844_ _04664_ _05527_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__nor2_1
X_14563_ screen.screenLogic.currentWrx vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11775_ net698 _04794_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_155_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ clknet_leaf_66_clk _00464_ net1270 vssd1 vssd1 vccd1 vccd1 datapath.PC\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_10726_ datapath.PC\[31\] _05563_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__xor2_1
XANTENNA__07654__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14494_ clknet_leaf_50_clk _01381_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13445_ clknet_leaf_82_clk _00401_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06862__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ _01507_ net660 _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_152_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ clknet_leaf_91_clk keypad.decode.button_n\[4\] net1205 vssd1 vssd1 vccd1
+ vccd1 keypad.apps.button\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07406__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10588_ _03308_ net346 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[0\]
+ sky130_fd_sc_hd__nor2_1
X_12327_ net1827 net214 net478 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
X_12258_ net216 net2475 net486 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11209_ net1539 net143 net137 _05113_ vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__a22o_1
X_12189_ _06436_ _06437_ _05851_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08119__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _01453_ _01576_ _01580_ _01495_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__o211a_2
XANTENNA__09660__A _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06681_ _01512_ net1031 net1007 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08420_ _01996_ _02040_ _03346_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_102_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08276__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ datapath.rf.registers\[8\]\[0\] _01775_ _03258_ _03259_ _03260_ vssd1 vssd1
+ vccd1 vccd1 _03278_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_129_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07302_ datapath.rf.registers\[7\]\[22\] net826 net807 datapath.rf.registers\[15\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ _01599_ _01669_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07645__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__A1 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07233_ datapath.rf.registers\[10\]\[24\] net918 net882 datapath.rf.registers\[17\]\[24\]
+ _02159_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a221o_1
XANTENNA__10745__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07164_ datapath.rf.registers\[6\]\[25\] net815 net750 datapath.rf.registers\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12960__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07095_ datapath.rf.registers\[22\]\[27\] net954 net887 datapath.rf.registers\[9\]\[27\]
+ _02021_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout202 _04666_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_2
Xfanout213 _05526_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
Xfanout235 _05665_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_1
Xfanout246 net248 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07030__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _04730_ _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nand2b_1
Xfanout257 net260 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout268 _05628_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_1
Xfanout279 _05613_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
X_07997_ _02911_ _02912_ _02914_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__or3_1
X_09736_ net846 _04661_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__nor2_2
X_06948_ _01871_ _01872_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__or3_1
X_09667_ net409 _04593_ net411 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21a_1
X_06879_ net999 net985 net980 net976 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__and4_4
XANTENNA_fanout831_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A _01820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ net497 net494 vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__nand2_2
XFILLER_0_139_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09598_ _02081_ net685 net678 _02085_ _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__o221ai_4
XANTENNA__07090__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ net528 net527 net406 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ screen.register.currentXbus\[31\] _05729_ _06025_ vssd1 vssd1 vccd1 vccd1
+ _06026_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08833__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07636__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _05396_ _05413_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11491_ _05927_ _05959_ _05681_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10655__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ clknet_leaf_77_clk net1308 net1247 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ _05356_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_133_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ clknet_leaf_13_clk _00153_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10373_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__inv_2
XANTENNA__08061__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12870__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ datapath.mulitply_result\[22\] datapath.multiplication_module.multiplicand_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13092_ clknet_leaf_16_clk _00084_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12043_ _06317_ _06318_ _06315_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_148_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_4
Xfanout791 net792 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_4
X_13994_ clknet_leaf_3_clk _00881_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12945_ net250 net2051 net541 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12876_ net261 net2213 net549 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09077__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ _05493_ net175 _06227_ net178 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11758_ screen.counter.ct\[22\] net667 net1019 _06175_ vssd1 vssd1 vccd1 vccd1 _00445_
+ sky130_fd_sc_hd__a22o_1
X_14546_ net1357 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XANTENNA__07627__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ datapath.PC\[29\] _05549_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14477_ clknet_leaf_0_clk _01364_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ screen.counter.currentCt\[17\] _06132_ net666 vssd1 vssd1 vccd1 vccd1 _06135_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13428_ clknet_leaf_89_clk _00384_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08588__A0 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13359_ clknet_leaf_99_clk _00344_ net1227 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12780__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08052__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07260__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ datapath.rf.registers\[21\]\[8\] net937 net855 datapath.rf.registers\[5\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__a22o_1
XANTENNA__07012__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ datapath.rf.registers\[11\]\[10\] net774 net717 datapath.rf.registers\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a22o_1
XANTENNA__11895__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__A0 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ _01614_ net650 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__nor2_2
X_07782_ datapath.rf.registers\[9\]\[11\] net778 net765 datapath.rf.registers\[17\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_09521_ _03977_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__or2_1
X_06733_ _01609_ _01610_ datapath.ru.latched_instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ _01660_ sky130_fd_sc_hd__mux2_1
XANTENNA__09304__A2 _04209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ net616 _04362_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__or2_1
X_06664_ _01477_ net1030 net1010 net1040 datapath.ru.latched_instruction\[4\] vssd1
+ vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a32o_1
X_08403_ _02521_ _03329_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__and2_1
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09383_ _04232_ _04277_ _04309_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__and3_1
X_06595_ _01415_ _01511_ _01519_ datapath.ru.latched_instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 _01525_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12955__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ datapath.rf.registers\[15\]\[0\] net995 _01746_ vssd1 vssd1 vccd1 vccd1 _03261_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07079__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08265_ datapath.rf.registers\[7\]\[1\] net959 net955 datapath.rf.registers\[22\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1154_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07216_ datapath.rf.registers\[4\]\[24\] net811 net724 datapath.rf.registers\[27\]\[24\]
+ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_99_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08196_ net506 _03120_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08172__C _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12690__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ datapath.rf.registers\[22\]\[26\] net953 net914 datapath.rf.registers\[18\]\[26\]
+ _02073_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07251__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ datapath.rf.registers\[8\]\[27\] net739 net716 datapath.rf.registers\[29\]\[27\]
+ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout879_A _01844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1008 net1010 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_4
XANTENNA__07003__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13346__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _03405_ _04645_ _04612_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__o21a_1
X_10991_ net631 _05666_ _05671_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__or3_4
XANTENNA__08628__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ net168 net2080 net571 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12661_ net189 net2457 net438 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XANTENNA__12865__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14400_ clknet_leaf_46_clk _01287_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11612_ screen.counter.ct\[7\] net1294 _06068_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and3_1
XANTENNA__07609__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12592_ net2057 net210 net446 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ screen.register.currentYbus\[6\] _05772_ _05777_ screen.register.currentYbus\[30\]
+ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_13_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ clknet_leaf_22_clk _01218_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14262_ clknet_leaf_26_clk _01149_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11474_ screen.register.currentXbus\[10\] net1016 net1014 screen.register.currentXbus\[18\]
+ _05733_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a221o_1
XANTENNA__07490__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ clknet_leaf_32_clk _00205_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ _05341_ _05342_ _05343_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08034__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14193_ clknet_leaf_27_clk _01080_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09231__A1 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ clknet_leaf_39_clk _00136_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10356_ screen.controlBus\[7\] screen.controlBus\[6\] vssd1 vssd1 vccd1 vccd1 _05278_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_148_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ clknet_leaf_61_clk _00067_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ _03307_ _03207_ net353 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__mux2_1
X_12026_ datapath.mulitply_result\[8\] datapath.multiplication_module.multiplicand_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__nor2_1
XANTENNA__09565__A1_N _03560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ clknet_leaf_60_clk _00864_ net1266 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12928_ net2009 net169 net546 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__mux2_1
XANTENNA__07848__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12775__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ net190 net2471 net555 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14529_ net1351 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ net510 _02973_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07481__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07001_ _01921_ _01923_ _01925_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__or4_1
XANTENNA__08516__A_N _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07233__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06802__A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10324__A _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net412 net341 _03471_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_110_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ _02826_ _02827_ _02828_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__or4_1
X_08883_ net376 _03808_ _03809_ net330 vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o211a_1
XANTENNA__08733__A0 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A _05544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ datapath.rf.registers\[26\]\[10\] net940 net904 datapath.rf.registers\[24\]\[10\]
+ _02760_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07765_ datapath.rf.registers\[24\]\[12\] net904 net872 datapath.rf.registers\[25\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
XANTENNA__09289__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06716_ datapath.ru.latched_instruction\[9\] net1039 _01642_ vssd1 vssd1 vccd1 vccd1
+ _01643_ sky130_fd_sc_hd__a21oi_4
X_09504_ _04391_ _04430_ net412 vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07696_ datapath.rf.registers\[31\]\[13\] net817 net782 datapath.rf.registers\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
XANTENNA__07839__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__C _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09435_ _02885_ _03318_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__xnor2_1
X_06647_ net1018 _01551_ _01575_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a21o_1
XANTENNA__12685__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09366_ net688 _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nand2_1
X_06578_ datapath.ru.latched_instruction\[21\] _01507_ vssd1 vssd1 vccd1 vccd1 _01508_
+ sky130_fd_sc_hd__nor2_1
X_08317_ datapath.rf.registers\[0\]\[1\] net827 _03228_ _03243_ vssd1 vssd1 vccd1
+ vccd1 _03244_ sky130_fd_sc_hd__o22a_4
XANTENNA__08264__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ net611 _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ _03163_ _03169_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or3_2
XANTENNA__07472__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08016__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ datapath.rf.registers\[15\]\[3\] net808 net795 datapath.rf.registers\[13\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__a22o_1
XANTENNA__10933__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _03977_ _04447_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nand2_1
XANTENNA__07224__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net1426 _05828_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10141_ net203 _05067_ net1309 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10072_ net705 _04540_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__and2_1
XANTENNA__08724__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13900_ clknet_leaf_35_clk _00787_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13831_ clknet_leaf_20_clk _00718_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13762_ clknet_leaf_51_clk _00649_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10974_ net245 net1954 net587 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12713_ net256 net1919 net569 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__mux2_1
XANTENNA__12595__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13693_ clknet_leaf_100_clk datapath.multiplication_module.multiplicand_i_n\[10\]
+ net1224 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12644_ net265 net2503 net436 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12575_ net1649 net278 net444 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__mux2_1
XANTENNA__10409__A _05048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11004__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14314_ clknet_leaf_15_clk _01201_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11526_ _05752_ _05807_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14245_ clknet_leaf_107_clk _01132_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11457_ _05680_ _05926_ _05928_ _05681_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__o22ai_1
XANTENNA__08007__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10408_ _05313_ _05314_ _05321_ _05329_ _05290_ vssd1 vssd1 vccd1 vccd1 screen.counter.ack
+ sky130_fd_sc_hd__a41o_2
XANTENNA__07215__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14176_ clknet_leaf_44_clk _01063_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11388_ screen.register.currentYbus\[13\] net132 _05879_ net161 vssd1 vssd1 vccd1
+ vccd1 _00371_ sky130_fd_sc_hd__a22o_1
X_10339_ net1470 keypad.decode.sticky\[1\] net1032 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky_n\[1\]
+ sky130_fd_sc_hd__mux2_1
X_13127_ clknet_leaf_25_clk _00119_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10144__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09507__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ clknet_leaf_33_clk _00050_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12009_ datapath.mulitply_result\[5\] datapath.multiplication_module.multiplicand_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__and2_1
X_07550_ net522 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06501_ datapath.PC\[23\] vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
XANTENNA__10825__A1 _01461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07481_ datapath.rf.registers\[3\]\[18\] net767 net741 datapath.rf.registers\[1\]\[18\]
+ _02393_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a221o_1
X_09220_ net373 net365 _03670_ _03671_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__nand4_1
XFILLER_0_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08284__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ net636 _04072_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__nand2_1
XANTENNA__08246__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ datapath.rf.registers\[10\]\[4\] net917 net913 datapath.rf.registers\[18\]\[4\]
+ _03022_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09082_ _02743_ _03322_ _02702_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07454__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08033_ datapath.rf.registers\[31\]\[6\] net817 net778 datapath.rf.registers\[9\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a22o_1
Xhold800 datapath.rf.registers\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold811 datapath.rf.registers\[5\]\[4\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout208_A _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07206__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 datapath.rf.registers\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 datapath.rf.registers\[8\]\[25\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 datapath.rf.registers\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 datapath.rf.registers\[17\]\[18\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 datapath.rf.registers\[12\]\[11\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold877 datapath.rf.registers\[1\]\[22\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 datapath.rf.registers\[18\]\[31\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _01433_ _01715_ _03567_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__a211o_1
Xhold899 datapath.rf.registers\[16\]\[25\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08935_ _03860_ _03861_ net340 vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21oi_1
X_08866_ _02324_ _02344_ net681 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a21o_1
XANTENNA__08459__A _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07817_ _02722_ net516 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__and2_1
X_08797_ net393 _03722_ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout744_A _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ _02662_ _02669_ _02673_ _02674_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_123_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10928__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ _02594_ _02601_ _02603_ _02605_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout911_A _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ net372 _04067_ _04343_ net377 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07693__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ _05538_ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__nor2_1
XANTENNA__06707__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08237__A2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09349_ net491 _04271_ net671 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_101_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07445__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12360_ net1925 net213 net474 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__mux2_1
XANTENNA__11241__B2 _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11311_ net124 _05398_ _05851_ vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XANTENNA__10638__A2_N _05494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12291_ net1971 _05519_ net483 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__mux2_1
XANTENNA__09737__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14030_ clknet_leaf_118_clk _00917_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09198__B1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11242_ net1513 net140 net134 _02926_ vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__a22o_1
X_11173_ _05769_ _05799_ _05818_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a2bb2o_1
X_10124_ _03573_ _05050_ net1051 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a21o_1
XANTENNA__13361__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ _03946_ _04448_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_3_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ clknet_leaf_26_clk _00701_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ clknet_leaf_15_clk _00632_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10957_ net163 net2348 net592 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__mux2_1
XANTENNA__09673__B2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ clknet_leaf_109_clk _00611_ net1106 vssd1 vssd1 vccd1 vccd1 columns.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ net165 net2451 net600 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__mux2_1
X_12627_ net2300 net192 net441 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07436__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12558_ net215 net2379 net449 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__mux2_1
X_11509_ _05681_ _05741_ _05968_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_151_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold107 screen.controlBus\[19\] vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ net230 net2222 net458 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__mux2_1
Xhold118 screen.controlBus\[27\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold129 datapath.multiplication_module.multiplicand_i\[18\] vssd1 vssd1 vccd1 vccd1
+ net1495 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ clknet_leaf_115_clk _01115_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ clknet_leaf_7_clk _01046_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 _05481_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_4
XANTENNA__10743__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10305__C net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06981_ _01885_ _01905_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__and2_1
XANTENNA__06962__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _03307_ _03458_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__nand2_1
XANTENNA__11299__B2 mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__A _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1199 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_2
X_08651_ datapath.PC\[14\] datapath.PC\[15\] _03577_ vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__or3_1
Xfanout1191 net1198 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11417__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__B _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ datapath.rf.registers\[13\]\[15\] net793 net735 datapath.rf.registers\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08582_ net992 _03061_ _03507_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07533_ datapath.rf.registers\[21\]\[17\] net936 net868 datapath.rf.registers\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08321__D1 _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07675__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ _02369_ net523 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ net363 _03921_ _03922_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12963__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08219__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07395_ _02315_ _02317_ _02319_ _02321_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__or4_1
XFILLER_0_146_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09134_ _03952_ _03953_ net396 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a21o_1
XANTENNA__07427__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09065_ _03895_ _03991_ net396 vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08016_ datapath.rf.registers\[12\]\[6\] net888 net884 datapath.rf.registers\[9\]\[6\]
+ _02940_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a221o_1
Xhold630 datapath.rf.registers\[0\]\[11\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 datapath.rf.registers\[25\]\[8\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 datapath.rf.registers\[11\]\[11\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 datapath.rf.registers\[18\]\[22\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 datapath.rf.registers\[24\]\[17\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 datapath.rf.registers\[23\]\[14\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 datapath.rf.registers\[4\]\[18\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_A _01851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ net221 _04562_ _04584_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a21o_1
XANTENNA__06953__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net371 _03710_ _03843_ net378 vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__o211a_1
XANTENNA__12203__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ _04766_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__xnor2_2
X_08849_ net639 _03773_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11860_ datapath.PC\[28\] net305 _06248_ _06250_ vssd1 vssd1 vccd1 vccd1 _00472_
+ sky130_fd_sc_hd__a22o_1
X_10811_ net841 _04007_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a21oi_2
X_11791_ net204 _05619_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__or2_1
XANTENNA__10658__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ clknet_leaf_86_clk _00480_ net1231 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07666__B1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10742_ _01423_ _04278_ net840 vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13461_ clknet_leaf_77_clk _00417_ net1249 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12873__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ _01503_ net660 _05524_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a22o_2
XANTENNA__09407__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ net1816 net270 net465 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__mux2_1
X_13392_ clknet_leaf_92_clk net1369 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12343_ net1718 net282 net472 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12274_ net1824 net286 net481 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11225_ net1465 net145 net139 _05030_ vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__a22o_1
X_14013_ clknet_leaf_24_clk _00900_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ _05266_ _05748_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_8_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06944__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ _04943_ _05030_ _05031_ _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__or4_1
X_11087_ _05721_ net1021 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nor2_4
X_10038_ net702 _03909_ _04449_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__nand3_1
XANTENNA__11952__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11989_ datapath.mulitply_result\[2\] datapath.multiplication_module.multiplicand_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13728_ clknet_leaf_94_clk datapath.multiplication_module.multiplier_i_n\[13\] net1206
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10256__A2 _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07657__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12783__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13659_ clknet_leaf_67_clk _00597_ net1258 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07409__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07180_ datapath.rf.registers\[20\]\[25\] net902 net898 datapath.rf.registers\[6\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07188__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
XANTENNA__07042__D1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _04721_ _04747_ _04720_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a21o_1
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
Xfanout439 _06462_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_4
X_09752_ _01640_ _04678_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__nor2_1
X_06964_ datapath.rf.registers\[20\]\[30\] net902 net862 datapath.rf.registers\[28\]\[30\]
+ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ net393 _03629_ _03520_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__o21a_1
X_09683_ _03565_ _03566_ net838 vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a21o_1
X_06895_ datapath.rf.registers\[11\]\[31\] net971 _01807_ _01815_ _01821_ vssd1 vssd1
+ vccd1 vccd1 _01822_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12958__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__A1 datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08634_ _03504_ net634 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nor2_1
XANTENNA__07896__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07360__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _03482_ _03491_ net418 vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XANTENNA__09098__C1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08456__B net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07516_ datapath.rf.registers\[4\]\[17\] net809 net718 datapath.rf.registers\[28\]\[17\]
+ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a221o_1
XANTENNA__10247__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ _03371_ _03419_ _02348_ _03369_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08175__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07447_ datapath.rf.registers\[19\]\[19\] net944 net908 datapath.rf.registers\[30\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a22o_1
XANTENNA__12693__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07378_ datapath.rf.registers\[30\]\[20\] net772 net747 datapath.rf.registers\[21\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a22o_1
X_09117_ _03323_ net613 _04009_ _04043_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_118_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08073__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08612__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06704__B _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09048_ net616 _03959_ _03971_ _03973_ net492 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07820__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10941__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 datapath.rf.registers\[19\]\[14\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 datapath.rf.registers\[13\]\[20\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net244 net1767 net584 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
XANTENNA__07179__A2 _02104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 datapath.rf.registers\[12\]\[20\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 datapath.rf.registers\[6\]\[14\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout940 net943 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_4
Xfanout951 _01813_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_4
Xfanout962 _01806_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_4
Xfanout973 _01732_ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_2
Xfanout984 _01654_ vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_2
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_51_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ net169 net2240 net543 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12868__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 datapath.rf.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 screen.register.currentXbus\[6\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net1456 _05897_ net157 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
Xhold1182 datapath.rf.registers\[26\]\[22\] vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07887__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 datapath.rf.registers\[2\]\[21\] vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ net188 net2072 net551 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
XANTENNA__07551__A _02457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11843_ _06237_ _06238_ datapath.PC\[23\] net304 vssd1 vssd1 vccd1 vccd1 _00467_
+ sky130_fd_sc_hd__a2bb2o_1
X_14562_ screen.dcx vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
X_11774_ net698 _04336_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__nand2_1
XANTENNA__07103__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ clknet_leaf_66_clk _00463_ net1270 vssd1 vssd1 vccd1 vccd1 datapath.PC\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_10725_ net842 _03565_ _03566_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14493_ clknet_leaf_33_clk _01380_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13444_ clknet_leaf_82_clk _00400_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ datapath.mulitply_result\[21\] net427 net662 vssd1 vssd1 vccd1 vccd1 _05511_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__08382__A _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11199__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587_ net423 _05333_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[15\]
+ sky130_fd_sc_hd__nor2_1
X_13375_ clknet_leaf_91_clk keypad.decode.button_n\[3\] net1205 vssd1 vssd1 vccd1
+ vccd1 keypad.apps.button\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11012__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12326_ net2215 net219 net479 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11947__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ net217 net2573 net486 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__mux2_1
XANTENNA__10851__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09564__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ net1459 net144 net138 _05154_ vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__a22o_1
X_12188_ columns.count\[7\] _06434_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11910__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__inv_2
XANTENNA__07590__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12778__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ mmio.memload_or_instruction\[30\] net1063 net1008 datapath.ru.latched_instruction\[30\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a32o_1
XANTENNA__07878__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ datapath.rf.registers\[12\]\[0\] net734 net719 datapath.rf.registers\[28\]\[0\]
+ _03276_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_22_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ datapath.rf.registers\[21\]\[22\] net747 net728 datapath.rf.registers\[2\]\[22\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08281_ _01602_ net839 _01645_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08842__A2 _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07232_ datapath.rf.registers\[22\]\[24\] net954 net894 datapath.rf.registers\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06805__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08055__B1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ datapath.rf.registers\[5\]\[25\] net785 net764 datapath.rf.registers\[17\]\[25\]
+ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07802__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ datapath.rf.registers\[7\]\[27\] net958 net942 datapath.rf.registers\[26\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout203 net205 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
Xfanout214 _05526_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_130_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06540__A mmio.memload_or_instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _05512_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_1
Xfanout236 _05665_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06908__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ datapath.PC\[3\] _03088_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__or2_1
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
Xfanout258 net260 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_89_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout269 net272 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
X_07996_ datapath.rf.registers\[14\]\[7\] net799 net770 datapath.rf.registers\[30\]\[7\]
+ _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a221o_1
XANTENNA__09307__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _04627_ _04659_ _04660_ net674 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a31o_1
XANTENNA__12688__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06947_ datapath.rf.registers\[14\]\[30\] net800 net763 datapath.rf.registers\[17\]\[30\]
+ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout657_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _01904_ net534 net405 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__mux2_1
X_06878_ net1001 net983 net978 net976 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__and4_1
X_08617_ _01681_ _03532_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout824_A _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ _02060_ _02080_ net682 vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08548_ _03448_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10936__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08479_ _03401_ _03402_ _02791_ _03381_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__o211a_1
X_10510_ _05405_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__and2_1
X_11490_ _05745_ _05959_ _05680_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08046__A0 _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ screen.register.currentXbus\[1\] screen.register.currentXbus\[0\] screen.register.currentXbus\[3\]
+ screen.register.currentXbus\[2\] vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10372_ _05277_ screen.controlBus\[7\] screen.controlBus\[6\] _05293_ vssd1 vssd1
+ vccd1 vccd1 _05294_ sky130_fd_sc_hd__and4bb_2
X_13160_ clknet_leaf_13_clk _00152_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ datapath.mulitply_result\[22\] datapath.multiplication_module.multiplicand_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__nand2_1
X_13091_ clknet_leaf_103_clk _00083_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12042_ datapath.mulitply_result\[10\] net325 net321 _06319_ vssd1 vssd1 vccd1 vccd1
+ _00585_ sky130_fd_sc_hd__a22o_1
Xhold290 datapath.rf.registers\[18\]\[4\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout770 net773 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
Xfanout781 _01762_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_4
Xfanout792 _01759_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12598__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13993_ clknet_leaf_2_clk _00880_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12944_ net253 net2507 net541 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__mux2_1
XANTENNA__10055__A_N _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ net266 net2383 net549 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
XANTENNA__11007__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ net833 _04784_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14545_ net1356 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_11757_ screen.counter.ct\[22\] _06074_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__or2_1
XANTENNA__10846__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09482__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10708_ net185 net1797 net607 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ clknet_leaf_31_clk _01363_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11688_ screen.counter.currentCt\[17\] _06132_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08037__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ clknet_leaf_88_clk _00383_ net1216 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10639_ net244 net2185 net607 vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08588__A1 _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_95_clk _00343_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ net2378 net284 net476 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__mux2_1
X_13289_ clknet_leaf_110_clk _00279_ net1106 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10147__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07850_ datapath.rf.registers\[18\]\[10\] net789 net730 datapath.rf.registers\[16\]\[10\]
+ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a221o_1
XANTENNA__08760__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ _01614_ _01727_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nor2_2
X_07781_ datapath.rf.registers\[6\]\[11\] net813 net755 datapath.rf.registers\[24\]\[11\]
+ _02704_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a221o_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06771__B1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ _04420_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nand2_1
X_06732_ datapath.ru.latched_instruction\[5\] _01589_ vssd1 vssd1 vccd1 vccd1 _01659_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07315__A2 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06663_ _01477_ net1029 net1010 net1040 datapath.ru.latched_instruction\[4\] vssd1
+ vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a32oi_4
X_09451_ net624 _04363_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08402_ _02526_ _02568_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__or3_1
X_06594_ datapath.ru.latched_instruction\[5\] _01499_ _01500_ vssd1 vssd1 vccd1 vccd1
+ _01524_ sky130_fd_sc_hd__and3_1
X_09382_ _04306_ _04308_ net670 _04279_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ datapath.rf.registers\[27\]\[0\] net988 _01763_ vssd1 vssd1 vccd1 vccd1 _03260_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout140_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout238_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08264_ datapath.rf.registers\[31\]\[1\] net951 net919 datapath.rf.registers\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10622__A2 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07215_ datapath.rf.registers\[9\]\[24\] net780 net747 datapath.rf.registers\[21\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12971__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ net506 _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_99_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07146_ datapath.rf.registers\[10\]\[26\] net917 net881 datapath.rf.registers\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08750__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07077_ datapath.rf.registers\[23\]\[27\] net787 net746 datapath.rf.registers\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1009 _01581_ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_4
XANTENNA_fanout774_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ net847 _01726_ _01611_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _04613_ _03385_ _03383_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__and3b_1
XANTENNA__12211__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ net165 net2389 net587 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ net637 _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12660_ net195 net2148 net437 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_67_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11611_ net1281 screen.counter.ct\[21\] net1280 _06073_ vssd1 vssd1 vccd1 vccd1 _06074_
+ sky130_fd_sc_hd__and4_1
XANTENNA__06580__C_N mmio.memload_or_instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10666__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12591_ net2524 net213 net445 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14330_ clknet_leaf_23_clk _01217_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11542_ screen.register.currentYbus\[22\] _05775_ _05776_ screen.register.currentYbus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire423 _02545_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
XANTENNA__08019__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14261_ clknet_leaf_28_clk _01148_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11473_ screen.register.currentYbus\[10\] _05776_ _05940_ _05941_ _05943_ vssd1 vssd1
+ vccd1 vccd1 _05944_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12881__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ clknet_leaf_58_clk _00204_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10424_ keypad.debounce.debounce\[9\] keypad.debounce.debounce\[8\] keypad.debounce.debounce\[11\]
+ keypad.debounce.debounce\[10\] vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__and4_1
X_14192_ clknet_leaf_0_clk _01079_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13143_ clknet_leaf_45_clk _00135_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ screen.controlBus\[5\] screen.controlBus\[4\] vssd1 vssd1 vccd1 vccd1 _05277_
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_76_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10286_ net317 _03942_ _04618_ net682 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__o22a_1
X_13074_ clknet_leaf_34_clk _00066_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12025_ datapath.mulitply_result\[8\] datapath.multiplication_module.multiplicand_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__and2_1
XANTENNA__08742__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ clknet_leaf_40_clk _00863_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12927_ net1730 net172 net547 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11960__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12858_ net194 net2189 net554 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__mux2_1
XANTENNA__08258__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ net834 _06213_ _06214_ _05095_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_107_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12789_ net215 net2479 net563 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14528_ net1350 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_32_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08046__S net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14459_ clknet_leaf_52_clk _01346_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12791__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07000_ datapath.rf.registers\[18\]\[29\] net791 _01926_ net832 vssd1 vssd1 vccd1
+ vccd1 _01927_ sky130_fd_sc_hd__a211o_1
XANTENNA__08570__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07784__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ _02479_ _03494_ net680 _03873_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_94_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10324__B _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07902_ datapath.rf.registers\[15\]\[9\] net806 net738 datapath.rf.registers\[8\]\[9\]
+ _02817_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__a221o_1
X_08882_ net373 _03674_ _03675_ net381 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a31o_1
XANTENNA__07536__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ datapath.rf.registers\[23\]\[10\] net932 _02757_ _02758_ _02759_ vssd1 vssd1
+ vccd1 vccd1 _02760_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12817__A0 _05496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ datapath.rf.registers\[6\]\[12\] net896 net884 datapath.rf.registers\[9\]\[12\]
+ _02690_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ _03654_ _03656_ net408 vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
X_06715_ _01514_ net1027 net1006 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__and3_1
XANTENNA__12966__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ datapath.rf.registers\[9\]\[13\] net778 net717 datapath.rf.registers\[29\]\[13\]
+ _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a221o_1
X_09434_ _02886_ _03399_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__xnor2_1
X_06646_ _01530_ _01551_ _01575_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _03067_ _03313_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__xnor2_1
X_06577_ net1305 net1303 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ _01507_ sky130_fd_sc_hd__or3b_4
XANTENNA_fanout522_A _02476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08316_ _03232_ _03234_ _03238_ _03242_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _05350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ net640 _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08247_ _03170_ _03171_ _03172_ _03173_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__or4_1
XFILLER_0_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08178_ datapath.rf.registers\[12\]\[3\] net993 _01776_ vssd1 vssd1 vccd1 vccd1 _03105_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout989_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ datapath.rf.registers\[8\]\[26\] net738 net720 datapath.rf.registers\[28\]\[26\]
+ _02055_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a221o_1
XANTENNA__12206__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _04797_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__nand2_1
XANTENNA__11308__A0 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _04988_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__and2_1
XANTENNA__11859__B2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07527__A2 _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13830_ clknet_leaf_106_clk _00717_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10819__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ clknet_leaf_43_clk _00648_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12876__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10973_ net249 net1728 net587 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12712_ net257 net2534 net569 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__mux2_1
XANTENNA__10295__B1 _03496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13692_ clknet_leaf_68_clk datapath.multiplication_module.multiplicand_i_n\[9\] net1225
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07160__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ net272 net1832 net437 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12574_ net2313 net280 net444 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__mux2_1
XANTENNA__10598__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14313_ clknet_leaf_3_clk _01200_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11525_ screen.register.currentXbus\[29\] net1013 _05989_ _05992_ vssd1 vssd1 vccd1
+ vccd1 _05993_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14244_ clknet_leaf_17_clk _01131_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09486__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11456_ _05925_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11547__B1 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ net1012 _05326_ _05328_ _05322_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ clknet_leaf_36_clk _01062_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11387_ _02633_ net669 vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__and2_1
XANTENNA__11020__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07766__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ clknet_leaf_111_clk _00118_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ _01404_ _05256_ _05253_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06974__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__B _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ clknet_leaf_41_clk _00049_ net1162 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ net508 net353 _04217_ net388 vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a211o_1
XANTENNA__07518__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ datapath.mulitply_result\[5\] datapath.multiplication_module.multiplicand_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__nor2_1
X_13959_ clknet_leaf_24_clk _00846_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12786__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06500_ datapath.PC\[22\] vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ datapath.rf.registers\[18\]\[18\] net790 net731 datapath.rf.registers\[16\]\[18\]
+ _02392_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a221o_1
XANTENNA__10825__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08284__B _03210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ net708 _04049_ net624 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10589__A1 _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ datapath.rf.registers\[3\]\[4\] net965 net881 datapath.rf.registers\[17\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__a22o_1
X_09081_ _02702_ _03407_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09424__A2_N net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08032_ datapath.rf.registers\[26\]\[6\] net820 net717 datapath.rf.registers\[29\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07909__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06813__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold801 datapath.rf.registers\[13\]\[27\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 datapath.rf.registers\[18\]\[21\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold823 datapath.rf.registers\[20\]\[26\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 datapath.rf.registers\[8\]\[27\] vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold845 datapath.rf.registers\[27\]\[11\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A2 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold856 datapath.rf.registers\[9\]\[20\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold867 datapath.rf.registers\[19\]\[26\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08954__B2 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold878 datapath.rf.registers\[24\]\[22\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 datapath.rf.registers\[8\]\[12\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _01715_ _03747_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__nor2_1
XANTENNA__06965__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ net401 _03854_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__or2_1
X_08865_ net415 _03789_ _03791_ net317 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout472_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08459__B _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07816_ _02722_ net516 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__nor2_1
X_08796_ _01904_ net352 _03627_ net388 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07390__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08178__C _01776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12696__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ datapath.rf.registers\[9\]\[12\] net778 net734 datapath.rf.registers\[12\]\[12\]
+ _02670_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout737_A _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09131__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07678_ datapath.rf.registers\[23\]\[14\] net932 net888 datapath.rf.registers\[12\]\[14\]
+ _02604_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a221o_1
XANTENNA__07142__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12018__A1 datapath.mulitply_result\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ net377 _03718_ _03719_ net333 vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__o211a_1
X_06629_ datapath.ru.latched_instruction\[12\] datapath.ru.latched_instruction\[13\]
+ datapath.ru.latched_instruction\[14\] datapath.ru.latched_instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout904_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06707__B _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ _04236_ _04270_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_43_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11241__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _04200_ _04201_ net374 vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11310_ net123 _05400_ _05851_ vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA__07996__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ net2166 net224 net482 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09198__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11241_ net1491 net140 net136 _02971_ vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__a22o_1
XANTENNA__10245__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10201__B1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _05726_ _05763_ _05819_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__and4b_1
X_10123_ _01426_ _03572_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ net1056 _03579_ _04980_ _04979_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a31o_1
XANTENNA__09370__A1 _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A2 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ clknet_leaf_28_clk _00700_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13744_ clknet_leaf_99_clk _00631_ net1227 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10956_ net168 net2442 net592 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__mux2_1
XANTENNA__07133__B1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13675_ clknet_leaf_109_clk _00610_ net1107 vssd1 vssd1 vccd1 vccd1 columns.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10887_ net169 datapath.rf.registers\[26\]\[30\] net601 vssd1 vssd1 vccd1 vccd1 _00081_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11015__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12626_ net1711 net197 net442 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__mux2_1
XANTENNA__09425__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11768__B1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11232__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ net218 net2404 net450 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ screen.register.currentXbus\[20\] _05707_ _05709_ screen.register.currentXbus\[12\]
+ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__a221o_1
XANTENNA__07987__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06633__A mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ net227 net1912 net457 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__mux2_1
Xhold108 net78 vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09189__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold119 datapath.multiplication_module.multiplicand_i\[16\] vssd1 vssd1 vccd1 vccd1
+ net1485 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ clknet_leaf_48_clk _01114_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11439_ screen.register.currentXbus\[8\] _05709_ _05777_ screen.register.currentYbus\[24\]
+ _05773_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07739__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14158_ clknet_leaf_119_clk _01045_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06947__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ clknet_leaf_28_clk _00101_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10305__D net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14089_ clknet_leaf_2_clk _00976_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_06980_ _01885_ _01905_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__or2_1
XANTENNA__11299__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1170 net1171 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_2
X_08650_ net1276 datapath.PC\[13\] _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__or3_2
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_4
Xfanout1192 net1198 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07911__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ datapath.rf.registers\[6\]\[15\] net814 net779 datapath.rf.registers\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a22o_1
X_08581_ net657 net640 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nand2_1
XANTENNA__09113__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07532_ datapath.rf.registers\[2\]\[17\] net920 net900 datapath.rf.registers\[20\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06808__A _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07463_ _02369_ net523 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ net367 _03919_ _03920_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ datapath.rf.registers\[24\]\[20\] net757 _02320_ net832 vssd1 vssd1 vccd1
+ vccd1 _02321_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09133_ _04058_ _04059_ net392 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__a21o_1
XANTENNA__11223__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10764__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout220_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09064_ net390 _03951_ _03990_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08015_ datapath.rf.registers\[26\]\[6\] net940 net936 datapath.rf.registers\[21\]\[6\]
+ _02938_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a221o_1
Xhold620 datapath.rf.registers\[1\]\[27\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 datapath.rf.registers\[9\]\[9\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 datapath.rf.registers\[0\]\[19\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold653 datapath.rf.registers\[27\]\[5\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 datapath.rf.registers\[26\]\[25\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold675 datapath.rf.registers\[2\]\[7\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 datapath.rf.registers\[22\]\[21\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 datapath.rf.registers\[24\]\[7\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09966_ net836 _04890_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08917_ net371 _03710_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__o21a_1
X_09897_ _04680_ _04681_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_96_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08155__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ net657 _03754_ _03774_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__and3_1
XANTENNA__07363__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _03339_ _03704_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or2_1
X_10810_ net841 _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11790_ net204 _04803_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__nand2_1
XANTENNA__07115__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ net1492 net288 net605 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_40_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ clknet_leaf_77_clk _00416_ net1247 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10670__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672_ datapath.mulitply_result\[23\] _01636_ net711 vssd1 vssd1 vccd1 vccd1 _05525_
+ sky130_fd_sc_hd__o21a_1
X_12411_ net1840 net276 net466 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
X_13391_ clknet_leaf_92_clk net1374 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10674__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__B1 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07969__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ net2259 net283 net472 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__mux2_1
XANTENNA__08091__A1 _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12273_ net1541 net295 net480 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ clknet_leaf_53_clk _00899_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11224_ net1421 net145 net139 _04920_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09591__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _05750_ _05803_ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_8_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ _04946_ _04953_ _04988_ _04997_ _04944_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__a221o_1
X_11086_ _05719_ net1020 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__nor2_4
Xclkbuf_leaf_87_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08146__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ datapath.PC\[18\] net1251 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__nor2_1
XANTENNA__07354__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ net322 _06273_ _06274_ net326 net2623 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a32o_1
XANTENNA__07106__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ clknet_leaf_95_clk datapath.multiplication_module.multiplier_i_n\[12\] net1206
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[12\] sky130_fd_sc_hd__dfrtp_1
X_10939_ net255 net2150 net590 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08854__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13658_ clknet_leaf_67_clk _00596_ net1258 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12609_ net2266 net276 net443 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XANTENNA__08606__A0 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06880__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13589_ clknet_leaf_79_clk _00539_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _04724_ _04726_ _04745_ _04723_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__a31o_1
Xfanout407 _03459_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09582__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout418 _03451_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_2
XANTENNA__12304__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_2
X_09751_ _01597_ net844 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__nand2_2
X_06963_ datapath.rf.registers\[12\]\[30\] net889 net854 datapath.rf.registers\[5\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_78_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_08702_ _03522_ _03525_ _03628_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_107_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09682_ _03637_ _04585_ _04608_ net836 vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a31o_1
XANTENNA__07345__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06894_ datapath.rf.registers\[23\]\[31\] net933 net931 datapath.rf.registers\[4\]\[31\]
+ _01818_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08633_ _01607_ _03353_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout170_A _05569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_A _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07641__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14458__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _03487_ _03490_ net411 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07515_ datapath.rf.registers\[25\]\[17\] net796 net722 datapath.rf.registers\[27\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a22o_1
XANTENNA__12974__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08495_ _02346_ _03369_ _03370_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1177_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10652__B1 _05506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07446_ datapath.rf.registers\[16\]\[19\] net962 net941 datapath.rf.registers\[26\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout602_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ _02282_ net526 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__nor2_2
XANTENNA__06871__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ net656 _04038_ _04042_ net491 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09047_ net688 _03973_ _03972_ net624 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09584__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 datapath.rf.registers\[7\]\[9\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 datapath.rf.registers\[4\]\[23\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 datapath.mulitply_result\[9\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__B2 _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08376__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 datapath.rf.registers\[12\]\[14\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12214__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07816__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold494 datapath.rf.registers\[25\]\[15\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07584__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 _01820_ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
Xfanout952 net955 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_8
X_09949_ _04855_ _04860_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__xnor2_1
Xfanout963 _01806_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10242__B _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
Xfanout974 _01732_ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08128__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout985 net986 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_2
X_12960_ net173 net2611 net542 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__mux2_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_51_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07336__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1150 datapath.rf.registers\[29\]\[12\] vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 datapath.rf.registers\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ _05896_ _06263_ net149 net1436 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__a22o_1
Xhold1172 datapath.rf.registers\[17\]\[20\] vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 datapath.rf.registers\[30\]\[20\] vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ net192 net2231 net551 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
Xhold1194 datapath.rf.registers\[17\]\[0\] vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10891__A0 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__B net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11842_ net208 _04831_ _05522_ _04663_ net304 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a221o_1
X_14561_ screen.csx vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11073__B _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ datapath.PC\[4\] net302 _06185_ _06187_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a22o_1
XANTENNA__12884__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08300__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13512_ clknet_leaf_66_clk _00462_ net1269 vssd1 vssd1 vccd1 vccd1 datapath.PC\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09759__A _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10724_ net167 net2267 net607 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__mux2_1
X_14492_ clknet_leaf_52_clk _01379_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13443_ clknet_leaf_83_clk _00399_ net1237 vssd1 vssd1 vccd1 vccd1 screen.csx sky130_fd_sc_hd__dfstp_1
XFILLER_0_126_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10655_ _03785_ _05509_ net845 vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__mux2_2
XANTENNA__06862__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13374_ clknet_leaf_91_clk keypad.decode.button_n\[2\] net1205 vssd1 vssd1 vccd1
+ vccd1 keypad.apps.button\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ net1401 _02587_ net351 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[14\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12325_ net1895 net222 net478 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
XANTENNA__10715__A1_N _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ net224 net2559 net485 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08367__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ net1451 net144 net138 _05134_ vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09564__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ _05850_ _06426_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__and2_1
XANTENNA__07575__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ net1023 _05710_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08119__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11963__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _05698_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_0_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12794__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07300_ datapath.rf.registers\[10\]\[22\] net750 _01775_ datapath.rf.registers\[8\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08280_ _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08573__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07231_ datapath.rf.registers\[20\]\[24\] net902 net879 datapath.rf.registers\[29\]\[24\]
+ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06805__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ datapath.rf.registers\[31\]\[25\] net819 net732 datapath.rf.registers\[16\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07093_ datapath.rf.registers\[3\]\[27\] net966 net850 datapath.rf.registers\[1\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06821__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout204 net205 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_130_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout215 _05526_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_130_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout226 _05502_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07566__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout237 _05665_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
X_09803_ datapath.PC\[3\] _03088_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__and2_1
XANTENNA__07030__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 _05654_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_1
XANTENNA__12969__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ datapath.rf.registers\[28\]\[7\] net718 net717 datapath.rf.registers\[29\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a22o_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09307__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _04627_ _04659_ _04660_ net674 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a31oi_4
XPHY_EDGE_ROW_105_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06946_ datapath.rf.registers\[23\]\[30\] net787 net723 datapath.rf.registers\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
XANTENNA__07318__B1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ _03456_ _04569_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__or2_1
X_06877_ net984 net978 _01803_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout552_A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08467__B net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _01682_ net617 vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nor2_2
X_09596_ net420 _04392_ _04393_ _03448_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ _03466_ _03473_ net421 vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout817_A _01747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _03381_ _03382_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07429_ datapath.rf.registers\[14\]\[19\] net800 net793 datapath.rf.registers\[13\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_114_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12209__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ screen.register.currentXbus\[5\] screen.register.currentXbus\[4\] screen.register.currentXbus\[7\]
+ screen.register.currentXbus\[6\] vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10371_ _05285_ _05291_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nor3_1
XANTENNA__10952__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ net323 _06375_ _06376_ net327 net1721 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13090_ clknet_leaf_43_clk _00082_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12041_ _06317_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_53_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold280 datapath.rf.registers\[21\]\[1\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 datapath.rf.registers\[10\]\[17\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07557__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_123_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout760 net762 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
Xfanout771 net773 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout782 _01761_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_4
X_13992_ clknet_leaf_13_clk _00879_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout793 _01757_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_29_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ net258 net1729 net541 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ net270 net1732 net551 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11825_ _01430_ net306 _06224_ _06226_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11408__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ net1355 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
X_11756_ net2627 net664 _06173_ _06174_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10707_ _05554_ _05553_ net710 _01459_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14475_ clknet_leaf_18_clk _01362_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11687_ _06088_ _06131_ _06133_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__and3_1
XANTENNA__11023__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13426_ clknet_leaf_87_clk _00382_ net1231 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10638_ _05495_ _05494_ net710 _01495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_95_clk _00342_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10862__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ _05405_ _05413_ _05426_ _05460_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12308_ net2419 net294 net476 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__mux2_1
X_13288_ clknet_leaf_92_clk _00278_ net1204 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07260__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ net296 net2485 net485 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__mux2_1
XANTENNA__11344__A1 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__C1 _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07012__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12789__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ net847 _01726_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__nor2_4
X_07780_ datapath.rf.registers\[21\]\[11\] net744 net740 datapath.rf.registers\[1\]\[11\]
+ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a221o_1
XANTENNA__08568__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ _01630_ _01631_ datapath.ru.latched_instruction\[13\] vssd1 vssd1 vccd1 vccd1
+ _01658_ sky130_fd_sc_hd__mux2_1
XANTENNA__09170__C1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ net638 _04367_ _04375_ _04376_ net655 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_84_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06662_ _01586_ _01587_ _01591_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_84_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ _02614_ _02656_ _03325_ _02610_ _02567_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__o311a_1
X_09381_ net613 _04282_ _04307_ _04303_ net671 vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__o311a_1
X_06593_ _01499_ _01500_ datapath.ru.latched_instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ _01523_ sky130_fd_sc_hd__a21oi_1
X_08332_ datapath.rf.registers\[3\]\[0\] net974 _01738_ vssd1 vssd1 vccd1 vccd1 _03259_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07079__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06816__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08263_ datapath.rf.registers\[27\]\[1\] net869 net867 datapath.rf.registers\[13\]\[1\]
+ _03187_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_15_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout133_A _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06535__B _01464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ datapath.rf.registers\[10\]\[24\] net750 net732 datapath.rf.registers\[16\]\[24\]
+ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ net646 _03118_ _03119_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_99_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07145_ datapath.rf.registers\[3\]\[26\] net965 net926 datapath.rf.registers\[8\]\[26\]
+ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1042_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07787__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ datapath.rf.registers\[10\]\[27\] net750 net736 datapath.rf.registers\[12\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11259__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07539__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A1 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07003__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ datapath.rf.registers\[0\]\[7\] net690 _02890_ _02904_ vssd1 vssd1 vccd1
+ vccd1 _02905_ sky130_fd_sc_hd__o22a_4
X_09717_ _04617_ _04642_ _04643_ _04614_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a22o_1
X_06929_ net1001 net984 net980 _01803_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__B _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09648_ net333 net377 _03800_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_143_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07711__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10947__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _03875_ _04505_ net417 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11610_ net1284 net1286 net1282 _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12590_ net2168 net219 net446 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ screen.register.currentXbus\[6\] _05704_ _06007_ vssd1 vssd1 vccd1 vccd1
+ _06008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14260_ clknet_leaf_115_clk _01147_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11472_ screen.register.currentYbus\[18\] _05775_ _05942_ vssd1 vssd1 vccd1 vccd1
+ _05943_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07490__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ clknet_leaf_52_clk _00203_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10423_ keypad.debounce.debounce\[13\] keypad.debounce.debounce\[12\] keypad.debounce.debounce\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and3_1
X_14191_ clknet_leaf_5_clk _01078_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07778__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ clknet_leaf_25_clk _00134_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10354_ screen.controlBus\[9\] screen.controlBus\[8\] screen.controlBus\[11\] screen.controlBus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13073_ clknet_leaf_8_clk _00065_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10285_ datapath.PC\[0\] _03286_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__or2_1
X_12024_ net2647 net326 net322 _06304_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__a22o_1
XANTENNA__11807__A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__B _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_8
X_13975_ clknet_leaf_45_clk _00862_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11018__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ net1678 net185 net546 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10857__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12857_ net197 net2402 net555 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ _04665_ _05640_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__or2_1
XANTENNA__06636__A mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ net218 net2029 net564 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11262__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11739_ _06084_ _06164_ _06163_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__o21ai_1
X_14527_ net1349 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_44_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10158__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09207__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07481__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ clknet_leaf_23_clk _01345_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11014__A0 _05519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07218__C1 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_87_clk _00365_ net1221 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14389_ clknet_leaf_30_clk _01276_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08570__B _03496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07233__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10605__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ net416 _03874_ _03876_ net318 vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07901_ datapath.rf.registers\[6\]\[9\] net814 net810 datapath.rf.registers\[4\]\[9\]
+ _02823_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a221o_1
X_08881_ net371 _03682_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ datapath.rf.registers\[19\]\[10\] net944 net912 datapath.rf.registers\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a22o_1
XANTENNA__12312__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07941__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ datapath.rf.registers\[26\]\[12\] net940 net916 datapath.rf.registers\[10\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a22o_1
X_09502_ net333 _04426_ _04427_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__o31a_1
XFILLER_0_154_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06714_ mmio.memload_or_instruction\[19\] net1058 net1004 datapath.ru.latched_instruction\[19\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07694_ datapath.rf.registers\[7\]\[13\] net824 net786 datapath.rf.registers\[23\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ _04191_ _04310_ _04336_ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__and4_1
X_06645_ _01562_ net1028 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout250_A _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09364_ _04289_ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__or2_2
X_06576_ _01417_ _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09446__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08315_ datapath.rf.registers\[18\]\[1\] net789 _03239_ _03240_ _03241_ vssd1 vssd1
+ vccd1 vccd1 _03242_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11253__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09295_ net340 _03860_ _03861_ _04220_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__a32o_1
XANTENNA_20 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout515_A _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1257_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08246_ datapath.rf.registers\[6\]\[2\] net816 _01777_ datapath.rf.registers\[12\]\[2\]
+ _03153_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07472__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ datapath.rf.registers\[17\]\[3\] _01735_ net972 vssd1 vssd1 vccd1 vccd1 _03104_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ datapath.rf.registers\[13\]\[26\] net793 net749 datapath.rf.registers\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a22o_1
XANTENNA__07224__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A _01841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ datapath.rf.registers\[7\]\[28\] net957 net933 datapath.rf.registers\[23\]\[28\]
+ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10070_ net202 _04990_ _04994_ _04996_ net1312 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a311o_1
XANTENNA__11859__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12222__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07932__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__B1 _05645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ clknet_leaf_48_clk _00647_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10972_ net254 net2141 net586 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ net263 net1959 net569 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__mux2_1
X_13691_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[8\] net1225
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12642_ net273 net1923 net439 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10047__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11244__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12573_ net1998 net283 net444 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12892__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11524_ screen.register.currentYbus\[29\] _05742_ _05990_ _05991_ vssd1 vssd1 vccd1
+ vccd1 _05992_ sky130_fd_sc_hd__a211o_1
XANTENNA__09767__A _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14312_ clknet_leaf_14_clk _01199_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire221 _04541_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_1
XFILLER_0_124_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14243_ clknet_leaf_104_clk _01130_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11455_ _05741_ _05746_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nand2_1
XANTENNA__12193__A _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ screen.counter.ct\[1\] _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07215__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14174_ clknet_leaf_51_clk _01061_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11386_ screen.register.currentYbus\[12\] net132 _05878_ net161 vssd1 vssd1 vccd1
+ vccd1 _00370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ clknet_leaf_93_clk _00117_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10337_ _05037_ _05081_ _05244_ _05259_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__nor4b_1
X_13056_ clknet_leaf_46_clk _00048_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ net317 _03880_ _05193_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__o211a_1
X_12007_ _06286_ _06287_ _06285_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__o21ba_1
X_10199_ datapath.PC\[8\] _04384_ net537 vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__mux2_1
XANTENNA__07923__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11971__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ clknet_leaf_111_clk _00845_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09676__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10286__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ net1616 net261 net545 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
XANTENNA__10286__B2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13889_ clknet_leaf_42_clk _00776_ net1162 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11235__B1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07439__C1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08100__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ datapath.rf.registers\[2\]\[4\] net921 net865 datapath.rf.registers\[13\]\[4\]
+ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__a221o_1
XANTENNA__10319__C _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ _04000_ _04006_ net672 vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__mux2_2
XANTENNA__07454__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08031_ datapath.rf.registers\[3\]\[6\] net766 net718 datapath.rf.registers\[28\]\[6\]
+ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12307__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06813__B _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold802 datapath.rf.registers\[12\]\[22\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07206__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 datapath.rf.registers\[26\]\[24\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 datapath.rf.registers\[28\]\[28\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 datapath.multiplication_module.multiplicand_i\[21\] vssd1 vssd1 vccd1 vccd1
+ net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 datapath.rf.registers\[13\]\[31\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 datapath.rf.registers\[24\]\[13\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold868 datapath.rf.registers\[11\]\[19\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ datapath.PC\[27\] net1271 _04905_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_
+ sky130_fd_sc_hd__o22a_1
Xhold879 datapath.rf.registers\[10\]\[27\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ _03858_ _03859_ net400 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08864_ net415 _03790_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07914__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ datapath.rf.registers\[0\]\[11\] net690 _02730_ _02741_ vssd1 vssd1 vccd1
+ vccd1 _02742_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_127_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12977__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ net533 net352 _03721_ net384 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout465_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ datapath.rf.registers\[3\]\[12\] net766 net740 datapath.rf.registers\[1\]\[12\]
+ _02664_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07677_ datapath.rf.registers\[3\]\[14\] net964 net928 datapath.rf.registers\[4\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
X_09416_ net374 _04200_ _04201_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__and3_1
X_06628_ datapath.ru.latched_instruction\[4\] datapath.ru.latched_instruction\[0\]
+ datapath.ru.latched_instruction\[1\] datapath.ru.latched_instruction\[2\] vssd1
+ vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07693__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11226__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ net640 _04267_ _04273_ net625 net653 vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a221oi_1
X_06559_ net1305 net1303 mmio.memload_or_instruction\[31\] vssd1 vssd1 vccd1 vccd1
+ _01489_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_43_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07445__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09278_ net361 _04202_ _04204_ net370 vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__a211o_1
X_08229_ datapath.rf.registers\[17\]\[2\] _01735_ net972 vssd1 vssd1 vccd1 vccd1 _03156_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12217__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11240_ net1510 net141 net136 _03017_ vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09198__A2 _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _05721_ _05728_ _05731_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a31o_1
XANTENNA__10960__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ _01426_ _04359_ net536 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08158__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ datapath.PC\[16\] _03578_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__nand2_1
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ clknet_leaf_113_clk _00699_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10268__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ net173 net2136 net593 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__mux2_1
X_13743_ clknet_leaf_8_clk _00630_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07133__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ clknet_leaf_109_clk _00609_ net1106 vssd1 vssd1 vccd1 vccd1 columns.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10886_ net172 net2500 net601 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ net1568 net211 net442 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07436__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ net222 net2174 net449 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ screen.register.currentXbus\[28\] _05700_ _05973_ _05975_ vssd1 vssd1 vccd1
+ vccd1 _05976_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07729__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ net242 net2510 net457 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__mux2_1
XANTENNA__06633__B mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold109 screen.controlBus\[10\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11438_ _05302_ _05781_ _05909_ net1017 _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__a221o_1
X_14226_ clknet_leaf_35_clk _01113_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11966__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ clknet_leaf_0_clk _01044_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10870__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _03060_ net669 vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10743__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09436__S net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13108_ clknet_leaf_116_clk _00100_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14088_ clknet_leaf_13_clk _00975_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08149__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13039_ clknet_leaf_3_clk _00031_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07464__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1163 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_2
Xfanout1171 net1199 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_2
Xfanout1182 net1185 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12797__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1198 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_2
X_07600_ datapath.rf.registers\[5\]\[15\] net784 net771 datapath.rf.registers\[30\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a22o_1
X_08580_ net654 _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__nor2_2
XFILLER_0_135_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10259__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ datapath.rf.registers\[22\]\[17\] net952 net895 datapath.rf.registers\[14\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06808__B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__B net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07462_ datapath.rf.registers\[0\]\[19\] net692 _02377_ _02388_ vssd1 vssd1 vccd1
+ vccd1 _02389_ sky130_fd_sc_hd__o22a_4
XANTENNA__07675__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09201_ net363 _03803_ _03804_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__and3_1
XANTENNA__11208__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07393_ datapath.rf.registers\[20\]\[20\] net803 net785 datapath.rf.registers\[5\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09132_ _02608_ net355 _03989_ net390 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a211o_1
XANTENNA__07427__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09063_ net519 net355 _03989_ net386 vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout213_A _05526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ datapath.rf.registers\[16\]\[6\] net960 net860 datapath.rf.registers\[28\]\[6\]
+ _02939_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold610 datapath.rf.registers\[25\]\[17\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold621 datapath.rf.registers\[13\]\[5\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold632 datapath.rf.registers\[12\]\[5\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 datapath.rf.registers\[22\]\[30\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10780__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 datapath.rf.registers\[29\]\[16\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold665 datapath.rf.registers\[4\]\[31\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1122_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 datapath.rf.registers\[29\]\[9\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10734__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__S net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 datapath.rf.registers\[27\]\[24\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 datapath.rf.registers\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _03590_ _04891_ net1053 vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout582_A _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net362 _03546_ net371 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__o21ai_1
X_09896_ _04817_ _04819_ _04821_ _04784_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__or4b_1
X_08847_ net337 _03763_ net316 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout847_A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ _03425_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12500__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _02634_ net518 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__nor2_1
X_10740_ _01464_ net709 _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07666__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ net842 _05522_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__o21ai_2
X_12410_ net1574 net279 net464 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ clknet_leaf_92_clk net1381 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08615__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ net2177 net294 net473 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12272_ net1624 net293 net481 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14011_ clknet_leaf_22_clk _00898_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11223_ net1405 net144 _05842_ vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_56_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09256__S net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net1281 net1282 net1290 net1285 vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_8_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ _04909_ _04963_ _05009_ _04986_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__or4b_1
X_11085_ _05711_ net1020 vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__nor2_4
X_10036_ datapath.PC\[20\] net1269 _04960_ _04962_ vssd1 vssd1 vccd1 vccd1 _04963_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12410__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ datapath.mulitply_result\[0\] datapath.multiplication_module.multiplicand_i\[0\]
+ _06271_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__a21o_1
X_13726_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[11\] net1206
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10938_ net259 net1929 net590 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__mux2_1
XANTENNA__07657__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08854__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10869_ net259 net1980 net598 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__mux2_1
XANTENNA__10865__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13657_ clknet_leaf_67_clk _00595_ net1258 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07409__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12608_ net2202 net277 net440 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
X_13588_ clknet_leaf_88_clk _00538_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ _05596_ net2394 net449 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07290__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14209_ clknet_leaf_41_clk _01096_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout408 net410 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_4
X_14541__1328 vssd1 vssd1 vccd1 vccd1 _14541__1328/HI net1328 sky130_fd_sc_hd__conb_1
Xfanout419 net421 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_2
X_09750_ _01599_ _01723_ _01614_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__o21ba_1
X_06962_ datapath.rf.registers\[9\]\[30\] net886 net878 datapath.rf.registers\[29\]\[30\]
+ _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a221o_1
X_08701_ _01904_ net352 _03627_ net384 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a211o_1
X_09681_ _04587_ _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06893_ net1002 net986 net981 _01808_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__and4_4
X_08632_ _01607_ _03353_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__and2_1
XANTENNA__12320__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07896__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06819__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08563_ _03488_ _03489_ net341 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__D_N net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ datapath.rf.registers\[15\]\[17\] net808 net733 datapath.rf.registers\[16\]\[17\]
+ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07648__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ _02346_ _03371_ _03419_ _02348_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07445_ datapath.rf.registers\[12\]\[19\] net888 net868 datapath.rf.registers\[27\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XANTENNA__10652__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07376_ _02302_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__inv_2
X_09115_ net634 _04033_ _04039_ net612 vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__o22a_1
XANTENNA__08073__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ _03327_ _03947_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07281__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07820__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold440 datapath.rf.registers\[27\]\[28\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 datapath.rf.registers\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 datapath.rf.registers\[0\]\[12\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold473 datapath.rf.registers\[4\]\[19\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 datapath.rf.registers\[3\]\[27\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 datapath.rf.registers\[7\]\[6\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net923 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_8
Xfanout931 _01820_ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08781__B1 _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_4
X_09948_ _04609_ _04869_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__o21bai_1
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_4
Xfanout964 net967 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_8
Xfanout975 _05797_ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_2
Xfanout986 _01653_ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_2
Xfanout997 _01647_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _04711_ _04712_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08533__A0 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1140 datapath.rf.registers\[11\]\[10\] vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 datapath.rf.registers\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 datapath.rf.registers\[5\]\[2\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _05895_ _06263_ net149 net1457 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__a22o_1
XANTENNA__12230__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 datapath.rf.registers\[10\]\[8\] vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ net196 net1622 net552 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
XANTENNA__07887__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1184 datapath.rf.registers\[21\]\[19\] vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 datapath.rf.registers\[19\]\[3\] vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ net837 _03747_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nor2_1
XANTENNA__09089__A1 _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14560_ net1333 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
X_11772_ _05593_ net175 _06186_ net177 vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__a22o_1
XANTENNA__07639__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13511_ clknet_leaf_74_clk _00461_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_10723_ _01492_ net661 _05567_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_24_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ clknet_leaf_22_clk _01378_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13442_ clknet_leaf_85_clk _00398_ net1237 vssd1 vssd1 vccd1 vccd1 screen.dcx sky130_fd_sc_hd__dfstp_1
X_10654_ datapath.PC\[21\] _05503_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11199__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13373_ clknet_leaf_93_clk keypad.decode.button_n\[1\] net1205 vssd1 vssd1 vccd1
+ vccd1 keypad.apps.button\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10585_ net1507 _02633_ net351 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[13\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07272__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ net1906 net230 net479 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ net233 net2188 net486 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__mux2_1
XANTENNA__12405__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ net1913 net143 net137 _05058_ vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12186_ _06434_ _06435_ _06426_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_71_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ _05703_ _05713_ net1021 vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a21o_1
X_11068_ net1301 net1300 vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08524__A0 _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net200 _04829_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__or3b_1
XFILLER_0_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07878__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08827__A1 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ clknet_leaf_57_clk datapath.multiplication_module.multiplicand_i_n\[26\]
+ net1257 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07230_ datapath.rf.registers\[4\]\[24\] net931 net922 datapath.rf.registers\[2\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10608__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__C _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ datapath.rf.registers\[25\]\[25\] net798 net772 datapath.rf.registers\[30\]\[25\]
+ _02086_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a221o_1
XANTENNA__08055__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ _02018_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__inv_2
XANTENNA__07802__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07015__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _04665_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08763__A0 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout216 _05526_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_1
X_09802_ datapath.PC\[4\] _03040_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__and2_1
Xfanout227 _05502_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_1
Xfanout238 net241 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
X_07994_ datapath.rf.registers\[10\]\[7\] net748 _02919_ _02920_ net831 vssd1 vssd1
+ vccd1 vccd1 _02921_ sky130_fd_sc_hd__a2111o_1
Xfanout249 _05650_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09307__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ net681 net685 _04658_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__mux2_1
X_06945_ datapath.rf.registers\[25\]\[30\] net798 net756 datapath.rf.registers\[24\]\[30\]
+ _01869_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a221o_1
X_06876_ _01672_ _01674_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__nor4_1
X_09664_ _01906_ net686 net678 _01910_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__o221a_1
XANTENNA__07869__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06549__A mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ net651 _03285_ _03286_ _03532_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a211o_1
X_09595_ net642 _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout545_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08049__A_N _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ _03469_ _03472_ net413 vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ _02789_ _03403_ _02790_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_137_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07428_ datapath.rf.registers\[24\]\[19\] net756 net727 datapath.rf.registers\[2\]\[19\]
+ _02354_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07359_ datapath.rf.registers\[3\]\[21\] net965 net926 datapath.rf.registers\[8\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09243__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07254__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ screen.controlBus\[0\] screen.controlBus\[1\] vssd1 vssd1 vccd1 vccd1 _05292_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ net400 _03729_ _03955_ net340 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12225__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ _06310_ _06311_ _06312_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07006__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08349__A3 _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 datapath.rf.registers\[22\]\[15\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 datapath.rf.registers\[25\]\[13\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08004__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 datapath.rf.registers\[24\]\[25\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout750 _01772_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_2
Xfanout783 _01761_ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_2
X_13991_ clknet_leaf_25_clk _00878_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout794 _01757_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_4
XANTENNA__11365__A _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ net263 net2119 net541 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12895__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ net275 net2038 net550 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__mux2_1
X_11824_ _04664_ _05662_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14543_ net1354 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_11755_ _06074_ net1019 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__and2b_1
XANTENNA__09482__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540__1327 vssd1 vssd1 vccd1 vccd1 _14540__1327/HI net1327 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_64_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07493__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ datapath.mulitply_result\[28\] net427 net660 vssd1 vssd1 vccd1 vccd1 _05554_
+ sky130_fd_sc_hd__a21oi_1
X_14474_ clknet_leaf_9_clk _01361_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11686_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ clknet_leaf_79_clk _00381_ net1233 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08037__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10637_ datapath.mulitply_result\[18\] net428 net662 vssd1 vssd1 vccd1 vccd1 _05495_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__09234__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13356_ clknet_leaf_95_clk _00341_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_10568_ keypad.apps.button\[4\] net1032 _05419_ _05460_ vssd1 vssd1 vccd1 vccd1 _05475_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08613__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ net1595 net293 net477 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap343_A _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ clknet_leaf_91_clk _00277_ net1204 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
X_10499_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__inv_2
X_12238_ net291 net2519 net487 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__mux2_1
XANTENNA__11974__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ net2563 net327 net323 _06425_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a22o_1
XANTENNA__06771__A2 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ datapath.ru.latched_instruction\[23\] net1039 net1007 _01655_ vssd1 vssd1
+ vccd1 vccd1 _01657_ sky130_fd_sc_hd__a22o_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08287__C _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ datapath.ru.latched_instruction\[5\] net1042 _01501_ net1009 vssd1 vssd1
+ vccd1 vccd1 _01591_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_84_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08400_ _02614_ _02656_ _03325_ _02610_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__o31a_1
X_09380_ net634 _04291_ _04304_ net612 vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__o22a_1
X_06592_ _01409_ _01456_ _01464_ _01407_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o22ai_1
XANTENNA__08584__A _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ datapath.rf.registers\[14\]\[0\] net994 _01752_ vssd1 vssd1 vccd1 vccd1 _03258_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06816__B _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11823__B1_N net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ datapath.rf.registers\[16\]\[1\] net960 net891 datapath.rf.registers\[12\]\[1\]
+ _03188_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__a221o_1
XANTENNA__07484__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07213_ datapath.rf.registers\[7\]\[24\] net826 net739 datapath.rf.registers\[8\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08193_ net646 _03118_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_144_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout126_A _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07144_ datapath.rf.registers\[21\]\[26\] net938 net870 datapath.rf.registers\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
XANTENNA__07236__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06832__A _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08984__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ datapath.rf.registers\[11\]\[27\] net776 net732 datapath.rf.registers\[16\]\[27\]
+ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout495_A _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07977_ _02899_ _02901_ _02903_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout662_A datapath.MemRead vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _02930_ _02977_ _03396_ _04616_ _02931_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a221o_1
X_06928_ net1001 net984 net980 _01808_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__and4_1
XANTENNA__09161__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _03448_ _04035_ _04568_ _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a211o_1
X_06859_ datapath.rf.registers\[30\]\[31\] net771 net760 datapath.rf.registers\[19\]\[31\]
+ _01784_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout927_A _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _03611_ _03616_ net411 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08529_ net409 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ screen.register.currentXbus\[30\] _05700_ _05707_ screen.register.currentXbus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07475__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10248__B _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ screen.register.currentXbus\[2\] _05704_ _05772_ screen.register.currentYbus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a22o_1
XANTENNA__08019__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire425 _01971_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_4
XANTENNA__10963__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ keypad.debounce.debounce\[2\] _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_
+ sky130_fd_sc_hd__and3_1
X_13210_ clknet_leaf_23_clk _00202_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07227__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ clknet_leaf_116_clk _01077_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ screen.controlBus\[13\] screen.controlBus\[12\] screen.controlBus\[15\] screen.controlBus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13141_ clknet_leaf_29_clk _00133_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10782__B1 _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ clknet_leaf_3_clk _00064_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10284_ net200 _05210_ _05183_ net1309 vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a211o_1
XANTENNA__08727__A0 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ _06302_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__xnor2_1
Xfanout580 _06266_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_8
Xfanout591 _05673_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_4
X_13974_ clknet_leaf_26_clk _00861_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12925_ net1889 net190 net547 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ net211 net1886 net555 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08608__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net205 _04811_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__nand2_1
XANTENNA__08258__A2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12787_ net223 net2178 net563 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__mux2_1
XANTENNA__06636__B mmio.memload_or_instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14526_ net1317 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XANTENNA__07466__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ net1289 _06078_ _06098_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11262__B2 _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11969__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14457_ clknet_leaf_61_clk _01344_ net1265 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10873__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ net667 _06119_ _06121_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13408_ clknet_leaf_87_clk _00364_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06652__A _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388_ clknet_leaf_116_clk _01275_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13339_ clknet_leaf_97_clk _00324_ net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10174__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07900_ _02814_ _02816_ _02819_ _02822_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_110_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ net375 _03805_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__and3_1
XANTENNA__08579__A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08194__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ datapath.rf.registers\[6\]\[10\] net896 net856 datapath.rf.registers\[15\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a22o_1
X_07762_ datapath.rf.registers\[20\]\[12\] net900 net860 datapath.rf.registers\[28\]\[12\]
+ _02688_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ net333 _04425_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nand2_1
X_06713_ mmio.memload_or_instruction\[19\] net1058 net1004 datapath.ru.latched_instruction\[19\]
+ net1037 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a32oi_4
XPHY_EDGE_ROW_142_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07693_ datapath.rf.registers\[2\]\[13\] net726 net722 datapath.rf.registers\[27\]\[13\]
+ _02619_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06644_ _01568_ _01570_ _01572_ _01573_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__or4_1
X_09432_ _04355_ _04358_ net670 _04340_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_154_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06827__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06575_ mmio.memload_or_instruction\[20\] net1058 vssd1 vssd1 vccd1 vccd1 _01505_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09363_ net376 _03808_ _03809_ net332 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__o211a_1
XANTENNA__09446__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_A _05496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ datapath.rf.registers\[13\]\[1\] net995 _01756_ vssd1 vssd1 vccd1 vccd1 _03241_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07457__B1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11253__B2 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _04214_ _04219_ net335 vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__o21a_1
XANTENNA_10 _03774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_21 net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ datapath.rf.registers\[7\]\[2\] net824 _03156_ _03157_ _03159_ vssd1 vssd1
+ vccd1 vccd1 _03172_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10783__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1152_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout508_A _03039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06680__A1 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ datapath.rf.registers\[26\]\[3\] net987 _01743_ vssd1 vssd1 vccd1 vccd1 _03103_
+ sky130_fd_sc_hd__and3_1
X_07127_ datapath.rf.registers\[22\]\[26\] net752 net746 datapath.rf.registers\[21\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a22o_1
XANTENNA__07377__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07058_ datapath.rf.registers\[18\]\[28\] net914 net858 datapath.rf.registers\[15\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout877_A _01844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12503__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09382__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10023__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__B2 _05648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net257 net2516 net586 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12710_ net268 net2335 net569 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__mux2_1
XANTENNA__07696__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13690_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[7\] net1224
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07160__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ net277 net2100 net436 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10047__A2 _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__B2 _02831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ net1602 net296 net446 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ clknet_leaf_20_clk _01198_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11523_ screen.register.currentXbus\[13\] net1016 _05736_ screen.register.currentYbus\[13\]
+ _05734_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14242_ clknet_leaf_33_clk _01129_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11454_ _05745_ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__nor2_1
XANTENNA__06472__A datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11547__A2 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net1295 _05299_ _01437_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a21o_1
X_11385_ _02677_ net669 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__and2_1
X_14173_ clknet_leaf_32_clk _01060_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07287__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13124_ clknet_leaf_102_clk _00116_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09783__A _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10336_ _05037_ _05168_ _05179_ _05257_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__and4bb_1
XANTENNA__06974__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12413__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _03248_ _03494_ net684 _03249_ _01633_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a221oi_1
X_13055_ clknet_leaf_37_clk _00047_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12006_ net322 _06288_ _06289_ net326 net1781 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__a32o_1
X_10198_ _04360_ _04383_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__nor2_1
XANTENNA__10868__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13957_ clknet_leaf_108_clk _00844_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09676__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ net1743 net266 net545 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13888_ clknet_leaf_50_clk _00775_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11272__B net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12839_ net278 net1648 net553 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11235__B2 _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ clknet_leaf_0_clk _01396_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08581__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08030_ datapath.rf.registers\[20\]\[6\] net804 net744 datapath.rf.registers\[21\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold803 datapath.rf.registers\[10\]\[12\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 datapath.rf.registers\[26\]\[14\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 datapath.rf.registers\[26\]\[23\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 datapath.rf.registers\[13\]\[7\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 datapath.rf.registers\[21\]\[11\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 datapath.rf.registers\[22\]\[13\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ net206 _04907_ net1313 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a21o_1
Xhold869 datapath.rf.registers\[8\]\[22\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06965__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _03727_ _03728_ net394 vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a21o_1
XANTENNA__12323__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A2 _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _03642_ _03658_ net412 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout193_A _05544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_150_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07814_ _02725_ _02726_ _02738_ _02740_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__or4_1
X_08794_ net501 net622 net490 net532 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__o211a_1
XANTENNA__09116__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07390__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ datapath.rf.registers\[4\]\[12\] net809 net737 datapath.rf.registers\[8\]\[12\]
+ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout458_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07678__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07676_ datapath.rf.registers\[22\]\[14\] net952 _02602_ vssd1 vssd1 vccd1 vccd1
+ _02603_ sky130_fd_sc_hd__a21o_1
XANTENNA__07142__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ net641 _04339_ _04341_ net625 vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o211a_1
X_06627_ datapath.ru.latched_instruction\[3\] datapath.ru.latched_instruction\[5\]
+ datapath.ru.latched_instruction\[6\] datapath.ru.latched_instruction\[7\] vssd1
+ vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout625_A _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06558_ mmio.memload_or_instruction\[31\] _01455_ vssd1 vssd1 vccd1 vccd1 _01488_
+ sky130_fd_sc_hd__and2_2
X_09346_ _04271_ _04272_ net641 vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11777__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06489_ datapath.ru.latched_instruction\[28\] vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
X_09277_ net507 net360 _04203_ net365 vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__o211a_1
XANTENNA__08642__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08228_ datapath.rf.registers\[4\]\[2\] net994 _01734_ vssd1 vssd1 vccd1 vccd1 _03155_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07850__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout994_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08159_ _03072_ _03084_ _03085_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11170_ _05731_ _05770_ _05802_ _05728_ _05810_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__o221a_1
XANTENNA__07602__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net1243 _05040_ _05047_ _05038_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a31o_1
XANTENNA__12233__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _01715_ _03946_ _04978_ net1051 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__o211a_1
XANTENNA__07381__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ clknet_leaf_49_clk _00698_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11373__A _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13742_ clknet_leaf_115_clk _00629_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07669__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ net186 net2190 net592 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__mux2_1
XANTENNA__07133__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ clknet_leaf_109_clk _00608_ net1106 vssd1 vssd1 vccd1 vccd1 columns.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ net187 net2012 net600 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09778__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ net1601 net214 net441 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11768__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08094__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12555_ net230 net2088 net450 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__mux2_1
XANTENNA__12408__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ screen.register.currentXbus\[4\] _05704_ _05974_ vssd1 vssd1 vccd1 vccd1
+ _05975_ sky130_fd_sc_hd__a21o_1
XANTENNA__07841__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ net235 net2341 net456 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14225_ clknet_leaf_7_clk _01112_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11437_ _05294_ _05767_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ clknet_leaf_30_clk _01043_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11368_ screen.register.currentYbus\[3\] net130 _05869_ net159 vssd1 vssd1 vccd1
+ vccd1 _00361_ sky130_fd_sc_hd__a22o_1
XANTENNA__06947__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_49_clk _00099_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ _05081_ _05166_ _05167_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__or4_1
XANTENNA__10452__A _02831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ clknet_leaf_21_clk _00974_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11299_ net20 net1047 net1036 mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1
+ vccd1 _00313_ sky130_fd_sc_hd__a22o_1
X_13038_ clknet_leaf_118_clk _00030_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_4
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_4
Xfanout1172 net1175 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_4
Xfanout1183 net1185 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
X_07530_ net650 _02456_ net627 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a21o_1
XANTENNA__08857__C1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08321__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08295__C _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07461_ _02372_ _02373_ _02385_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09200_ _02978_ net680 _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a21boi_1
X_07392_ datapath.rf.registers\[31\]\[20\] net819 net811 datapath.rf.registers\[4\]\[20\]
+ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ net517 net355 _04057_ net386 vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__a211o_1
XANTENNA__08085__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06824__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09062_ net499 net620 net488 net518 vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o211a_1
XANTENNA__07832__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ datapath.rf.registers\[24\]\[6\] net904 net872 datapath.rf.registers\[25\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold600 datapath.multiplication_module.multiplicand_i\[7\] vssd1 vssd1 vccd1 vccd1
+ net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 datapath.rf.registers\[14\]\[12\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 datapath.rf.registers\[17\]\[8\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold633 datapath.rf.registers\[5\]\[12\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 datapath.rf.registers\[11\]\[25\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06840__A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__A1 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold655 datapath.rf.registers\[12\]\[8\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 datapath.rf.registers\[31\]\[16\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 datapath.rf.registers\[6\]\[27\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 datapath.rf.registers\[25\]\[26\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 datapath.rf.registers\[24\]\[11\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ datapath.PC\[28\] _03589_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1115_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _03448_ _03841_ _03839_ _03837_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a211o_1
X_09895_ _04817_ _04819_ _04821_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout575_A _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08846_ net329 _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__and2_1
XANTENNA__07363__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout742_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _03366_ _03367_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ net518 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07115__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ _02577_ _02578_ _02582_ _02585_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or4_1
XFILLER_0_138_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ net842 _03747_ net429 vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08076__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ net391 _04178_ _04255_ net399 vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__a211o_1
XANTENNA__12228__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08615__A2 _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ net2253 net292 net475 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__A1_N net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12271_ net1555 net298 net481 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__mux2_1
XANTENNA__10971__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14010_ clknet_leaf_23_clk _00897_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09576__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11222_ _01404_ _05256_ _05838_ _04931_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_56_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ net1291 screen.counter.ct\[17\] _05749_ _05751_ vssd1 vssd1 vccd1 vccd1 _05803_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_56_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ _04964_ _04975_ _05018_ net1311 _05010_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__o221ai_1
X_11084_ _05724_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__or2_2
XANTENNA__12898__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ net208 _04961_ net1312 vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a21o_1
XANTENNA__07354__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__inv_2
XANTENNA__07106__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13725_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[10\] net1206
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[10\] sky130_fd_sc_hd__dfrtp_1
X_10937_ net262 net2269 net590 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ clknet_leaf_67_clk _00594_ net1262 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10868_ net263 net2424 net598 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__mux2_1
XANTENNA__08067__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ net1947 net282 net440 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XANTENNA__09301__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10447__A _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ clknet_leaf_89_clk _00537_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ _04081_ _05631_ net844 vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ net291 net2351 net451 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__mux2_1
XANTENNA__11977__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10881__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12469_ net181 net1726 net456 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XANTENNA__09955__B _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14208_ clknet_leaf_48_clk _01095_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ clknet_leaf_52_clk _01026_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06603__A2_N _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ datapath.rf.registers\[6\]\[30\] net897 _01887_ net695 vssd1 vssd1 vccd1
+ vccd1 _01888_ sky130_fd_sc_hd__a211o_1
X_08700_ net501 net622 net490 net534 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__o211a_1
XANTENNA__12601__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _04589_ _04602_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_107_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06892_ net1000 net984 net979 _01808_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__and4_1
XANTENNA__07345__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08631_ _01584_ net847 vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__nand2_2
X_14556__1329 vssd1 vssd1 vccd1 vccd1 _14556__1329/HI net1329 sky130_fd_sc_hd__conb_1
XANTENNA__06819__B _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ _01860_ _01904_ net405 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07513_ datapath.rf.registers\[26\]\[17\] net823 net786 datapath.rf.registers\[23\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ _03371_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout156_A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10652__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07444_ datapath.rf.registers\[4\]\[19\] net930 net865 datapath.rf.registers\[13\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06835__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08058__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07375_ _02282_ net526 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout323_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1065_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ net624 _04010_ _04011_ net301 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__o31a_1
XANTENNA__07805__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09045_ net642 _03970_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and2_1
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold430 datapath.rf.registers\[21\]\[4\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 datapath.rf.registers\[28\]\[18\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 datapath.rf.registers\[18\]\[2\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 datapath.rf.registers\[25\]\[27\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 datapath.rf.registers\[7\]\[8\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 datapath.rf.registers\[19\]\[7\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 datapath.rf.registers\[17\]\[28\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 _01831_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_4
XANTENNA__07584__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout921 net923 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_4
Xfanout932 net935 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_8
X_09947_ net836 _04871_ _04873_ net206 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a31o_1
Xfanout943 _01816_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_4
XANTENNA_fanout957_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net967 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_4
XANTENNA__12865__A0 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout987 net988 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_2
X_09878_ _04787_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 datapath.rf.registers\[20\]\[18\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07336__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1141 datapath.rf.registers\[23\]\[13\] vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 datapath.rf.registers\[14\]\[13\] vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ net533 net352 _03721_ net388 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a211o_1
Xhold1163 datapath.rf.registers\[30\]\[28\] vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06544__B1 _01473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 datapath.rf.registers\[12\]\[31\] vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 datapath.rf.registers\[10\]\[11\] vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 datapath.rf.registers\[29\]\[27\] vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ datapath.PC\[22\] net304 _06236_ _04922_ vssd1 vssd1 vccd1 vccd1 _00466_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13349__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06583__C_N mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10966__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ net835 _04791_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__nand2_1
X_13510_ clknet_leaf_74_clk _00460_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ datapath.mulitply_result\[30\] net427 net661 vssd1 vssd1 vccd1 vccd1 _05568_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_24_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14490_ clknet_leaf_23_clk _01377_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ clknet_leaf_89_clk _00397_ net1214 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
X_10653_ net231 net2437 net608 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__mux2_1
X_13372_ clknet_leaf_91_clk keypad.decode.button_n\[0\] net1204 vssd1 vssd1 vccd1
+ vccd1 keypad.apps.button\[0\] sky130_fd_sc_hd__dfrtp_1
X_10584_ net1402 _02677_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[12\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net1839 net228 net478 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
X_12254_ net228 net2309 net485 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__mux2_1
XANTENNA__10159__A1 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ net2014 net143 net137 _05069_ vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12185_ columns.count\[6\] _06433_ _05850_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08772__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ _05723_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__nand2_1
XANTENNA__06783__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11826__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ net1300 net1301 _05701_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__or3_2
XANTENNA__12421__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__A1 _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _04783_ _04784_ _04822_ _04825_ _04828_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a41o_1
XANTENNA__06639__B mmio.memload_or_instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ net218 net2592 net581 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
X_13708_ clknet_leaf_56_clk datapath.multiplication_module.multiplicand_i_n\[25\]
+ net1257 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__B2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13639_ clknet_leaf_70_clk _00577_ net1228 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07160_ datapath.rf.registers\[13\]\[25\] net794 net767 datapath.rf.registers\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07091_ net648 _02016_ net626 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06821__C _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10116__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09801_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__inv_2
XANTENNA__07566__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08763__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_2
Xfanout228 _05502_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
X_07993_ datapath.rf.registers\[4\]\[7\] net809 net755 datapath.rf.registers\[24\]\[7\]
+ _02908_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a221o_1
Xfanout239 net241 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_1
XANTENNA__10455__D_N net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ _03445_ _01634_ _04628_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__mux2_1
XANTENNA__12331__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06944_ datapath.rf.registers\[9\]\[30\] net779 net735 datapath.rf.registers\[12\]\[30\]
+ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a221o_1
XANTENNA__07318__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _01885_ _01904_ _03497_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__o21ai_1
X_06875_ net1002 net984 net979 _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__and4_2
XANTENNA__08110__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _01646_ _03246_ net617 vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09594_ _02085_ _03430_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08545_ _03470_ _03471_ net408 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout440_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout538_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _03401_ _03402_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__nor2_1
XANTENNA__06565__A mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ datapath.rf.registers\[17\]\[19\] net763 net738 datapath.rf.registers\[8\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout705_A _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07358_ datapath.rf.registers\[6\]\[21\] net897 net853 datapath.rf.registers\[5\]\[21\]
+ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10815__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12506__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ datapath.rf.registers\[5\]\[22\] net785 net716 datapath.rf.registers\[29\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09028_ net400 _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08203__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 datapath.rf.registers\[26\]\[7\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 datapath.rf.registers\[21\]\[2\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 datapath.rf.registers\[20\]\[7\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07557__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 datapath.rf.registers\[25\]\[19\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 net743 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
XANTENNA__07962__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout751 net754 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_4
Xfanout762 _01769_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
XANTENNA__12241__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13990_ clknet_leaf_106_clk _00877_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout773 _01765_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout784 _01761_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
Xfanout795 _01757_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_4
XANTENNA__11365__B _03175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ net267 net2334 net541 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ net279 net2301 net549 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__mux2_1
XANTENNA__08955__A _03877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07190__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ net833 _03909_ net303 vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_119_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_139_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09467__C1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__A _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ net1353 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11754_ net1279 _06086_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__A2 _04408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _04584_ _05551_ net845 vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14473_ clknet_leaf_2_clk _01360_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ screen.counter.currentCt\[15\] screen.counter.currentCt\[16\] _06128_ vssd1
+ vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ clknet_leaf_81_clk _00380_ net1235 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ _04471_ _05492_ net845 vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13355_ clknet_leaf_95_clk _00340_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_140_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12416__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ _05470_ _05472_ _05474_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[3\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ net1619 net299 net477 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ clknet_leaf_109_clk _00276_ net1106 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
X_10498_ net35 net36 _05344_ _05346_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__and4b_1
X_12237_ net297 net2428 net484 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ _06423_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__xnor2_1
X_11119_ net1016 _05762_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__or3_1
XANTENNA__10460__A _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ datapath.mulitply_result\[20\] datapath.multiplication_module.multiplicand_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__nand2_1
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06660_ _01501_ net1009 datapath.ru.latched_instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ _01590_ sky130_fd_sc_hd__a21o_1
XANTENNA__07181__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06591_ datapath.ru.latched_instruction\[9\] _01515_ _01468_ datapath.ru.latched_instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ datapath.rf.registers\[17\]\[0\] _01735_ net972 vssd1 vssd1 vccd1 vccd1 _03257_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06816__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08261_ datapath.rf.registers\[21\]\[1\] net937 net857 datapath.rf.registers\[15\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__a22o_1
XANTENNA__07484__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07212_ datapath.rf.registers\[18\]\[24\] net791 net768 datapath.rf.registers\[3\]\[24\]
+ _02138_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08192_ net650 _03088_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07143_ datapath.rf.registers\[7\]\[26\] net957 net853 datapath.rf.registers\[5\]\[26\]
+ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__a221o_1
XANTENNA__12326__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06832__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07787__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__A1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ datapath.rf.registers\[5\]\[27\] net785 net757 datapath.rf.registers\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06995__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1028_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ datapath.rf.registers\[8\]\[7\] net924 net876 datapath.rf.registers\[29\]\[7\]
+ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__a221o_1
X_09715_ _03125_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__nand2_1
XANTENNA__11185__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06927_ datapath.rf.registers\[8\]\[31\] net926 net858 datapath.rf.registers\[15\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout655_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ net422 _04571_ _04572_ net318 vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__o211a_1
X_06858_ datapath.rf.registers\[31\]\[31\] net818 net720 datapath.rf.registers\[28\]\[31\]
+ _01745_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a221o_1
XANTENNA__07172__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07711__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09577_ net689 _04501_ _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a21oi_1
X_06789_ _01606_ _01607_ _01618_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ _03246_ _01646_ _03446_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08459_ _03287_ _03307_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__nor2_1
XANTENNA__08672__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10248__C _04277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11470_ screen.register.currentXbus\[18\] _05707_ _05709_ screen.register.currentXbus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__a22o_1
XANTENNA__14411__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10421_ keypad.debounce.debounce\[1\] keypad.debounce.debounce\[0\] keypad.debounce.debounce\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__and3_1
XANTENNA__12236__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ clknet_leaf_113_clk _00132_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10231__B1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ _05265_ _05266_ _05269_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06986__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13071_ clknet_leaf_12_clk _00063_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ datapath.PC\[1\] _05209_ _05184_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__mux2_1
XANTENNA__08727__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _06297_ _06298_ _06295_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13364__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _06464_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
Xfanout581 _06266_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09137__D1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout592 _05673_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_8
X_13973_ clknet_leaf_32_clk _00860_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09152__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ net2104 net193 net546 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__mux2_1
XANTENNA__10837__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07702__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ net215 net2468 net554 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__mux2_1
XANTENNA__06910__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11806_ net1487 net303 _06210_ _06212_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ net230 net2372 net564 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__mux2_1
X_14525_ net1316 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_11737_ net1289 net665 vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__nand2_1
XANTENNA__11262__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14456_ clknet_leaf_39_clk _01343_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13407_ clknet_leaf_86_clk _00363_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619_ net1509 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[31\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10455__A _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ clknet_leaf_59_clk _01274_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06652__B net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11599_ net1012 _05763_ _06062_ _06061_ _05798_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__a311o_1
XANTENNA__08966__A1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ clknet_leaf_96_clk _00323_ net1218 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ clknet_leaf_90_clk _00259_ net1209 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08194__A2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ datapath.rf.registers\[31\]\[10\] net948 net872 datapath.rf.registers\[25\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a22o_1
XANTENNA__08298__C _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07941__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ datapath.rf.registers\[17\]\[12\] net880 net868 datapath.rf.registers\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a22o_1
X_09500_ net376 _04132_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nor2_1
X_06712_ datapath.ru.latched_instruction\[22\] net1039 net1006 _01637_ vssd1 vssd1
+ vccd1 vccd1 _01639_ sky130_fd_sc_hd__a22o_2
X_07692_ datapath.rf.registers\[13\]\[13\] net795 net748 datapath.rf.registers\[10\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ net491 _04339_ _04356_ _04357_ net670 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__o221a_1
X_06643_ _01460_ _01563_ _01569_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06827__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ net380 _04030_ _04287_ _04288_ net331 vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__o221a_1
X_06574_ datapath.ru.latched_instruction\[19\] _01494_ vssd1 vssd1 vccd1 vccd1 _01504_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08313_ datapath.rf.registers\[10\]\[1\] net995 _01743_ vssd1 vssd1 vccd1 vccd1 _03240_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11253__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _04060_ _04061_ net401 vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_11 _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ datapath.rf.registers\[2\]\[2\] net729 net722 datapath.rf.registers\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a22o_1
XANTENNA_33 _01848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08175_ datapath.rf.registers\[23\]\[3\] net987 _01739_ vssd1 vssd1 vccd1 vccd1 _03102_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ datapath.rf.registers\[19\]\[26\] net760 net715 datapath.rf.registers\[29\]\[26\]
+ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06968__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07057_ datapath.rf.registers\[25\]\[28\] net873 net849 datapath.rf.registers\[1\]\[28\]
+ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07932__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__inv_2
X_10970_ net261 net2239 net586 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__mux2_1
XANTENNA__10819__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07145__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ net635 _04553_ _04554_ net611 vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12640_ net282 net2637 net439 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ net2455 net293 net447 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__mux2_1
XANTENNA__11244__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_50_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
X_14310_ clknet_leaf_106_clk _01197_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11522_ screen.register.currentXbus\[21\] net1015 _05737_ screen.register.currentYbus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__a22o_1
XANTENNA__07999__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ clknet_leaf_41_clk _01128_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11453_ screen.register.currentYbus\[9\] _05736_ _05921_ _05924_ vssd1 vssd1 vccd1
+ vccd1 _05925_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10404_ net1299 net1292 net1285 _05325_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__and4b_1
X_14172_ clknet_leaf_57_clk _01059_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11384_ screen.register.currentYbus\[11\] net131 _05877_ net160 vssd1 vssd1 vccd1
+ vccd1 _00369_ sky130_fd_sc_hd__a22o_1
XANTENNA__06959__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13123_ clknet_leaf_104_clk _00115_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10335_ _05037_ _05257_ _05259_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__and3b_1
XANTENNA__09783__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07081__C1 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ clknet_leaf_52_clk _00046_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11818__B _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10266_ _01632_ _03248_ _03249_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or3b_1
Xfanout1310 net1311 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlymetal6s2s_1
X_12005_ _06285_ _06286_ _06287_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__o21ai_1
X_10197_ net703 _04385_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nand2_1
XANTENNA__07384__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ clknet_leaf_14_clk _00843_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07136__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12907_ net1645 net270 net547 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13887_ clknet_leaf_38_clk _00774_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12838_ net282 net2183 net553 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11235__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12769_ net293 net1584 net561 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__mux2_1
XANTENNA__10884__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08100__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14508_ clknet_leaf_30_clk _01395_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ clknet_leaf_24_clk _01326_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold804 datapath.rf.registers\[8\]\[14\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 datapath.rf.registers\[24\]\[19\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 datapath.rf.registers\[19\]\[11\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11943__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold837 datapath.rf.registers\[11\]\[5\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 datapath.rf.registers\[8\]\[26\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12604__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ _04841_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nand2_1
Xhold859 datapath.rf.registers\[25\]\[9\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
X_08931_ _03856_ _03857_ net392 vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ net412 _03655_ _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09903__A3 _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ datapath.rf.registers\[7\]\[11\] net956 net920 datapath.rf.registers\[2\]\[11\]
+ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__a221o_1
XANTENNA__07914__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08793_ net377 _03718_ _03719_ net329 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout186_A _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ datapath.rf.registers\[13\]\[12\] net795 net748 datapath.rf.registers\[10\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
XANTENNA__07127__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__C1 _03202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11474__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ datapath.rf.registers\[9\]\[14\] net884 net876 datapath.rf.registers\[29\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a22o_1
XANTENNA__08875__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09414_ net641 _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__nand2_1
X_06626_ _01552_ _01553_ _01554_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14074__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09345_ _03182_ _03387_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__xnor2_2
X_06557_ net1305 net1304 mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ _01487_ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout520_A _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1262_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_43_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ net498 net495 net506 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__a21o_1
X_06488_ datapath.ru.latched_instruction\[27\] vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08227_ datapath.rf.registers\[13\]\[2\] net994 _01756_ vssd1 vssd1 vccd1 vccd1 _03154_
+ sky130_fd_sc_hd__and3_1
X_08158_ datapath.rf.registers\[16\]\[3\] net961 net880 datapath.rf.registers\[17\]\[3\]
+ _03070_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__a221o_1
XANTENNA__11934__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ _02029_ _02031_ _02033_ _02035_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__or4_1
X_08089_ net832 _03013_ _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__or4_1
XANTENNA__12514__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10120_ net698 _05042_ _05046_ net203 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a211o_1
XANTENNA__08158__A2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10051_ _01429_ net537 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__or2_1
XANTENNA__07366__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ clknet_leaf_36_clk _00697_ net1149 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07118__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ clknet_leaf_1_clk _00628_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10953_ net189 net2508 net593 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__mux2_1
XANTENNA__08866__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10673__B1 _05524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ clknet_leaf_109_clk _00607_ net1107 vssd1 vssd1 vccd1 vccd1 columns.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ net190 net2205 net601 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__mux2_1
XANTENNA__08963__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12623_ net2416 net219 net442 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12554_ net228 net2234 net449 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ screen.register.currentYbus\[4\] _05772_ _05776_ screen.register.currentYbus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12485_ net240 net1989 net458 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14224_ clknet_leaf_4_clk _01111_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11436_ screen.register.currentYbus\[0\] _05737_ _05905_ _05907_ _05908_ vssd1 vssd1
+ vccd1 vccd1 _05909_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14155_ clknet_leaf_68_clk _01042_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12424__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ _03118_ net668 vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ clknet_leaf_35_clk _00098_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ _05179_ _05244_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__or2_1
X_14086_ clknet_leaf_114_clk _00973_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ net19 net1045 net1034 mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1
+ vccd1 _00312_ sky130_fd_sc_hd__o22a_1
XANTENNA__10452__B _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08149__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ clknet_leaf_119_clk _00029_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ net203 _05173_ _05174_ _05175_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or4_1
XANTENNA__07357__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1140 net1143 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_4
Xfanout1151 net1164 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_4
Xfanout1162 net1163 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_2
XANTENNA__10879__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1173 net1175 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1198 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_2
XFILLER_0_135_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13939_ clknet_leaf_59_clk _00826_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08321__A2 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07460_ datapath.rf.registers\[17\]\[19\] net881 net878 datapath.rf.registers\[29\]\[19\]
+ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a221o_1
XANTENNA__10664__B1 _05513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08609__A0 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11208__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ datapath.rf.registers\[9\]\[20\] net780 net742 datapath.rf.registers\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ net499 net620 net488 net516 vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09061_ net335 _03631_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08012_ datapath.rf.registers\[23\]\[6\] net932 net928 datapath.rf.registers\[4\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 datapath.mulitply_result\[18\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold612 datapath.rf.registers\[19\]\[0\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold623 datapath.rf.registers\[9\]\[16\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12334__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 datapath.rf.registers\[7\]\[28\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold645 datapath.rf.registers\[4\]\[1\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 datapath.rf.registers\[23\]\[6\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06840__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 datapath.rf.registers\[22\]\[1\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ net539 _04584_ _04889_ net1057 vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a211o_1
Xhold678 datapath.rf.registers\[20\]\[9\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 datapath.rf.registers\[27\]\[19\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ net419 _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nor2_1
X_09894_ _04763_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1108_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ net381 _03771_ _03764_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A _06465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1216_A mmio.memload_or_instruction\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net673 _03638_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ datapath.rf.registers\[0\]\[13\] _02653_ net691 vssd1 vssd1 vccd1 vccd1 _02654_
+ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_A _01777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10655__A0 _03785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07658_ _02572_ _02573_ _02583_ _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07520__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06609_ datapath.ru.latched_instruction\[15\] _01462_ _01494_ datapath.ru.latched_instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12509__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ datapath.rf.registers\[26\]\[16\] net942 net911 datapath.rf.registers\[30\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a22o_1
XANTENNA__10818__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ net389 _03816_ _04158_ net396 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__A2 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09259_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10029__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ net2513 net289 net481 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__mux2_1
X_11221_ net1462 net145 net139 _04954_ vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12244__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07587__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ _05028_ _05029_ datapath.PC\[24\] net1268 vssd1 vssd1 vccd1 vccd1 _05030_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11257__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083_ _05708_ net1020 vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07339__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _04783_ _04826_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11985_ datapath.mulitply_result\[0\] datapath.multiplication_module.multiplicand_i\[0\]
+ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__and3_1
X_13724_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[9\] net1206
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[9\] sky130_fd_sc_hd__dfrtp_1
X_10936_ net265 net2535 net590 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__mux2_1
XANTENNA__07511__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10867_ net268 net1941 net598 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__mux2_1
X_13655_ clknet_leaf_67_clk _00593_ net1258 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12419__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12606_ net1987 net285 net440 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13586_ clknet_leaf_88_clk _00536_ net1216 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__inv_2
XANTENNA__10447__B _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12537_ net297 net1866 net451 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _05479_ _05575_ net577 vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__or3_1
XANTENNA__09016__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07290__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11419_ net535 net714 vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__nor2_1
X_14207_ clknet_leaf_36_clk _01094_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12399_ net171 net2162 net470 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
XANTENNA__10177__A2 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07578__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ clknet_leaf_23_clk _01025_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07042__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ clknet_leaf_28_clk _00956_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_06960_ datapath.rf.registers\[8\]\[30\] net927 net865 datapath.rf.registers\[13\]\[30\]
+ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_3_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_06891_ datapath.rf.registers\[26\]\[31\] net941 net939 datapath.rf.registers\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a22o_1
X_08630_ _01584_ net847 vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06819__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ net534 net533 net405 vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
X_07512_ datapath.rf.registers\[6\]\[17\] net813 net759 datapath.rf.registers\[19\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
X_08492_ _02436_ _03415_ _03416_ _03372_ _02434_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__o311a_1
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07443_ _02369_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__inv_2
XANTENNA__12329__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06835__B _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07374_ datapath.rf.registers\[0\]\[21\] net692 _02288_ _02300_ vssd1 vssd1 vccd1
+ vccd1 _02301_ sky130_fd_sc_hd__o22a_4
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09113_ net639 _04033_ _04038_ _04039_ net653 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06608__A2 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ net611 _03968_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07281__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__A1 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 datapath.rf.registers\[15\]\[13\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 datapath.rf.registers\[24\]\[28\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1225_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 datapath.rf.registers\[25\]\[18\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 datapath.rf.registers\[11\]\[17\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold464 datapath.rf.registers\[15\]\[15\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 datapath.rf.registers\[6\]\[13\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 datapath.rf.registers\[8\]\[9\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net903 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__buf_4
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold497 datapath.rf.registers\[31\]\[17\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 _01831_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_4
X_09946_ _03592_ _04872_ net1052 vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a21o_1
Xfanout933 net935 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_4
Xfanout944 net947 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout955 _01810_ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07682__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
Xfanout977 _01681_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__buf_4
XANTENNA_fanout852_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1120 datapath.rf.registers\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ _04801_ _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__nand2_1
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_2
Xfanout999 _01641_ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_51_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 datapath.rf.registers\[1\]\[31\] vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 datapath.rf.registers\[28\]\[27\] vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 datapath.rf.registers\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _02079_ net352 _03725_ net384 vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a211o_1
Xhold1164 datapath.rf.registers\[8\]\[6\] vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 datapath.rf.registers\[30\]\[29\] vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 datapath.rf.registers\[27\]\[22\] vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 datapath.mulitply_result\[31\] vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ _01904_ _01860_ net353 vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__mux2_1
X_11770_ net698 _04309_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09402__A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ _04608_ _05565_ net846 vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__mux2_2
XFILLER_0_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12239__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ clknet_leaf_89_clk _00396_ net1213 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
X_10652_ _01505_ net710 _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__o22a_2
XFILLER_0_76_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13371_ clknet_leaf_90_clk _00356_ net1211 vssd1 vssd1 vccd1 vccd1 keypad.apps.app_c\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10982__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ net1444 _02721_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[11\]
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12322_ net2062 net242 net478 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XANTENNA__07272__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11379__A _02831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net243 net2612 net485 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__mux2_1
X_11204_ net1701 net143 net137 _05079_ vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ columns.count\[6\] _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11135_ _05779_ _05783_ _05784_ _05712_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__and4b_1
XANTENNA__12702__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ net1300 net1301 _05701_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__nor3_1
X_10017_ _01431_ net1269 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07732__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06639__C mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11968_ net224 net1968 net580 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13707_ clknet_leaf_56_clk datapath.multiplication_module.multiplicand_i_n\[24\]
+ net1257 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10919_ net186 net1806 net596 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__mux2_1
X_11899_ net1453 _05884_ net156 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10458__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09237__A0 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13638_ clknet_leaf_70_clk _00576_ net1229 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10892__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ clknet_leaf_88_clk _00519_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07799__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ net343 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__inv_2
XANTENNA__07263__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11347__A1 mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07015__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ datapath.PC\[5\] _02998_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__and2_1
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_130_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout218 _05519_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12612__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07992_ datapath.rf.registers\[22\]\[7\] net751 net744 datapath.rf.registers\[21\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a22o_1
Xfanout229 _05502_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__S net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _03440_ _04586_ _04625_ _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a31o_1
X_06943_ datapath.rf.registers\[6\]\[30\] net815 net810 datapath.rf.registers\[4\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
XANTENNA__08515__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10132__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _03350_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__nand2_1
X_06874_ _01677_ _01678_ _01673_ _01675_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__o211a_1
XANTENNA__07723__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _01645_ _03247_ net617 vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__mux2_1
X_09593_ _03344_ _04519_ net642 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout266_A _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ _03207_ _03307_ net404 vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _02931_ _03398_ _03383_ _02884_ _02930_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout433_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07426_ datapath.rf.registers\[11\]\[19\] net775 net741 datapath.rf.registers\[1\]\[19\]
+ _02352_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07357_ datapath.rf.registers\[31\]\[21\] net949 net914 datapath.rf.registers\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout600_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07254__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06581__A mmio.memload_or_instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ datapath.rf.registers\[6\]\[22\] net815 net811 datapath.rf.registers\[4\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
X_09027_ net396 _03952_ _03953_ _03949_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 datapath.rf.registers\[22\]\[11\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07006__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 datapath.multiplication_module.multiplicand_i\[29\] vssd1 vssd1 vccd1 vccd1
+ net1627 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold272 datapath.rf.registers\[7\]\[4\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 datapath.rf.registers\[12\]\[7\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 datapath.rf.registers\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12522__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net733 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 net743 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_4
Xfanout752 net753 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_4
X_09929_ datapath.PC\[30\] _01728_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06550__C_N mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 _01767_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout774 net777 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
Xfanout785 _01761_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_4
Xfanout796 _01755_ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
X_12940_ net269 net1676 net543 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__mux2_1
XANTENNA__07714__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ net282 net2293 net549 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
XANTENNA__10977__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ net205 _04821_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11381__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _06086_ _06172_ net664 net1502 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a2bb2o_1
X_14541_ net1328 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__11274__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11813__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10704_ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11684_ screen.counter.currentCt\[15\] screen.counter.currentCt\[14\] _06126_ screen.counter.currentCt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__a31o_1
X_14472_ clknet_leaf_13_clk _01359_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07493__A2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ clknet_leaf_80_clk _00379_ net1235 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10635_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__inv_2
Xmax_cap1003 _01624_ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_2
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13354_ clknet_leaf_95_clk _00339_ net1206 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10566_ _05402_ _05434_ _05473_ net1026 _01444_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12305_ net2011 net287 net477 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__mux2_1
X_13285_ clknet_leaf_64_clk _00275_ net1272 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
X_10497_ net36 _05344_ _05346_ net35 vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__and4b_1
XANTENNA__11329__A1 mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12236_ net287 net1716 net484 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08745__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12432__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ datapath.mulitply_result\[31\] datapath.multiplication_module.multiplicand_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_112_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ _05728_ _05766_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nor2_1
X_12098_ net324 _06365_ _06366_ net328 net1857 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__a32o_1
XANTENNA__10460__B _02812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ _05264_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__or2_2
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XANTENNA__10887__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06590_ datapath.ru.latched_instruction\[10\] _01481_ _01480_ datapath.ru.latched_instruction\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11265__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08130__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ datapath.rf.registers\[9\]\[1\] net885 net848 datapath.rf.registers\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a22o_1
XANTENNA__06816__D net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07484__A2 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07211_ datapath.rf.registers\[30\]\[24\] net771 net721 datapath.rf.registers\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a22o_1
X_08191_ _03109_ _03114_ _03117_ _03089_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o31a_4
XFILLER_0_43_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12607__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07142_ datapath.rf.registers\[23\]\[26\] net933 net921 datapath.rf.registers\[2\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__a22o_1
XANTENNA__07236__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08984__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ datapath.rf.registers\[7\]\[27\] net826 net798 datapath.rf.registers\[25\]\[27\]
+ _01997_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12342__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ datapath.rf.registers\[4\]\[7\] net928 net892 datapath.rf.registers\[14\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a22o_1
X_06926_ net1002 net984 net978 _01812_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__and4_4
X_09714_ _03123_ _03181_ _04615_ _04640_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__o22a_1
X_09645_ net422 _03789_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06857_ datapath.rf.registers\[25\]\[31\] net797 net790 datapath.rf.registers\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout550_A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09576_ net707 _04502_ net623 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a21o_1
X_06788_ net537 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__inv_2
X_08527_ net504 _03446_ _03452_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11256__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ _02881_ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07475__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11008__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ datapath.rf.registers\[3\]\[20\] net966 net859 datapath.rf.registers\[15\]\[20\]
+ _02335_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a221o_1
X_08389_ _03019_ _03315_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__nand2_1
XANTENNA__12517__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ keypad.debounce.debounce\[5\] keypad.debounce.debounce\[4\] keypad.debounce.debounce\[7\]
+ keypad.debounce.debounce\[6\] vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__and4_1
XANTENNA__07227__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10351_ net1287 net1288 _05270_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13070_ clknet_leaf_2_clk _00062_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10282_ _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08188__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ _06300_ _06301_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12252__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _06467_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_4
Xfanout571 _06464_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_6
Xfanout582 _05675_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_8
X_13972_ clknet_leaf_113_clk _00859_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout593 _05673_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10298__A1 _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ net2273 net196 net547 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__mux2_1
XANTENNA__08360__B1 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ net218 net1984 net555 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11247__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11805_ _05635_ net175 _06211_ net178 vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12785_ net229 net1883 net563 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__mux2_1
XANTENNA__08112__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14524_ net1315 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11736_ net1290 net665 _06162_ net713 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a22o_1
XANTENNA__07466__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ clknet_leaf_45_clk _01342_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11667_ screen.counter.currentCt\[9\] screen.counter.currentCt\[10\] _06116_ vssd1
+ vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_12_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12427__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13406_ clknet_leaf_80_clk _00362_ net1234 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ net1627 net346 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[30\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07218__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _05679_ _05747_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nor2_1
X_14386_ clknet_leaf_35_clk _01273_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07110__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13337_ clknet_leaf_94_clk _00322_ net1205 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_4
X_10549_ _05403_ _05406_ _05416_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13268_ clknet_leaf_90_clk _00258_ net1209 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08179__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11567__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12219_ net234 net2515 net573 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13199_ clknet_leaf_6_clk _00191_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07926__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ datapath.rf.registers\[11\]\[12\] net968 net924 datapath.rf.registers\[8\]\[12\]
+ _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a221o_1
X_06711_ datapath.ru.latched_instruction\[22\] net1043 net1006 _01637_ vssd1 vssd1
+ vccd1 vccd1 _01638_ sky130_fd_sc_hd__a22oi_4
XANTENNA__11486__B1 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07691_ datapath.rf.registers\[30\]\[13\] net770 net759 datapath.rf.registers\[19\]\[13\]
+ _02615_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a221o_1
X_09430_ net634 _04347_ _04353_ net612 vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__o22a_1
XFILLER_0_149_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06642_ mmio.memload_or_instruction\[17\] mmio.memload_or_instruction\[18\] _01566_
+ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__or4b_1
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11238__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06827__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ net373 _04283_ _04284_ net376 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06573_ _01502_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__inv_2
XANTENNA__08103__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ datapath.rf.registers\[20\]\[1\] net990 _01734_ vssd1 vssd1 vccd1 vccd1 _03239_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07457__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ net394 _04216_ _04218_ net400 vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ datapath.rf.registers\[25\]\[2\] _01755_ net762 datapath.rf.registers\[19\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a22o_1
XANTENNA_23 _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12337__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout229_A _05502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ datapath.rf.registers\[10\]\[3\] net993 _01743_ vssd1 vssd1 vccd1 vccd1 _03101_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07209__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ datapath.rf.registers\[31\]\[26\] net818 net810 datapath.rf.registers\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a22o_1
X_07056_ datapath.rf.registers\[22\]\[28\] net953 net905 datapath.rf.registers\[24\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_A _05668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout765_A _01767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12800__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _02881_ _02883_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__or2_2
XANTENNA__08786__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__B1 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ net1001 net986 net979 _01808_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout932_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ datapath.rf.registers\[25\]\[9\] net797 net771 datapath.rf.registers\[30\]\[9\]
+ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ net637 _04553_ _04554_ _04552_ net657 vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__o2111a_1
XANTENNA__07696__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11229__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ net334 _04155_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__nor2_1
X_12570_ net1868 net299 net447 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__mux2_1
XANTENNA__07448__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ screen.register.currentXbus\[5\] _05720_ _05735_ screen.register.currentYbus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a22o_1
X_14569__1339 vssd1 vssd1 vccd1 vccd1 _14569__1339/HI net1339 sky130_fd_sc_hd__conb_1
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12247__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11452_ screen.register.currentYbus\[1\] _05737_ _05922_ _05923_ vssd1 vssd1 vccd1
+ vccd1 _05924_ sky130_fd_sc_hd__a211o_1
X_14240_ clknet_leaf_46_clk _01127_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10403_ net1282 net1279 _05323_ _05324_ _05300_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a41o_1
X_14171_ clknet_leaf_54_clk _01058_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11383_ _02721_ net668 vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__and2_1
XANTENNA__10990__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10755__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _05037_ _05257_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__and3b_1
XANTENNA__07865__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ clknet_leaf_33_clk _00114_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11387__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ clknet_leaf_32_clk _00045_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _01621_ _05191_ _03916_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__o21ba_1
Xfanout1300 screen.counter.ct\[1\] vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__clkbuf_2
X_12004_ _06285_ _06286_ _06287_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__or3_1
Xfanout1311 _01451_ vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__clkbuf_2
X_10196_ net1276 net1250 _05119_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__o22a_1
XANTENNA__12710__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 _03522_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
X_13955_ clknet_leaf_104_clk _00842_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12906_ net2005 net275 net548 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13886_ clknet_leaf_50_clk _00773_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ net286 net2093 net556 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07439__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12768_ net298 net1818 net561 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14507_ clknet_leaf_18_clk _01394_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11719_ net1294 net665 _06152_ net712 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10466__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ _05478_ net630 _06443_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__or3_4
XFILLER_0_142_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14438_ clknet_leaf_108_clk _01325_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold805 datapath.rf.registers\[17\]\[27\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ clknet_leaf_44_clk _01256_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold816 datapath.rf.registers\[27\]\[31\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold827 datapath.rf.registers\[27\]\[17\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold838 datapath.rf.registers\[2\]\[31\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07611__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 datapath.rf.registers\[4\]\[22\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ net527 net354 _03758_ net390 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ net414 _03662_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__or2_1
X_07812_ datapath.rf.registers\[23\]\[11\] net932 net904 datapath.rf.registers\[24\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a22o_1
XANTENNA__12620__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ net377 _03547_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07743_ datapath.rf.registers\[7\]\[12\] net824 net805 datapath.rf.registers\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
XANTENNA__06838__B _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ datapath.rf.registers\[11\]\[14\] net968 net908 datapath.rf.registers\[30\]\[14\]
+ _02599_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a221o_1
XANTENNA__07678__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06625_ datapath.ru.latched_instruction\[24\] datapath.ru.latched_instruction\[25\]
+ datapath.ru.latched_instruction\[26\] datapath.ru.latched_instruction\[27\] vssd1
+ vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__or4_1
X_09413_ _02932_ _03398_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout346_A _05333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06556_ net1305 net1303 mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1 vccd1
+ _01486_ sky130_fd_sc_hd__or3b_1
X_09344_ _03182_ _03311_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_43_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09230__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09275_ net511 _02997_ net360 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06487_ datapath.ru.latched_instruction\[23\] vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout513_A _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ datapath.rf.registers\[26\]\[2\] net989 _01743_ vssd1 vssd1 vccd1 vccd1 _03153_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_145_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07850__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10095__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _03077_ _03079_ _03081_ _03083_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07108_ datapath.rf.registers\[20\]\[27\] net902 net866 datapath.rf.registers\[13\]\[27\]
+ _02034_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a221o_1
X_08088_ datapath.rf.registers\[9\]\[5\] net781 net748 datapath.rf.registers\[10\]\[5\]
+ _02999_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07602__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ datapath.rf.registers\[13\]\[28\] net793 net787 datapath.rf.registers\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
X_10050_ _04817_ _04819_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__xor2_1
XANTENNA__09355__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13740_ clknet_leaf_32_clk _00627_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07669__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ net192 net2363 net592 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__mux2_1
XANTENNA__10673__A1 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ clknet_leaf_97_clk net426 net1220 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.mul_prev
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10985__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ net193 net2347 net600 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__mux2_1
XANTENNA__08963__B _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12622_ net1720 net222 net441 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12553_ net242 net2399 net449 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__mux2_1
XANTENNA__08094__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09291__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11504_ screen.register.currentYbus\[20\] _05775_ _05777_ screen.register.currentYbus\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a22o_1
XANTENNA__07841__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ net248 net2173 net457 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14223_ clknet_leaf_5_clk _01110_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11435_ screen.register.currentYbus\[16\] _05735_ _05736_ screen.register.currentYbus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__a22o_1
XANTENNA__09794__B _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12705__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ net2650 net130 _05868_ net159 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__a22o_1
X_14154_ clknet_leaf_9_clk _01041_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10317_ _05181_ _05211_ _05236_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a211o_1
X_13105_ clknet_leaf_7_clk _00097_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14085_ clknet_leaf_108_clk _00972_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11297_ net18 net1046 net1035 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1
+ vccd1 _00311_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10452__C _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ net699 _04232_ _04277_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__and3_1
X_13036_ clknet_leaf_34_clk _00028_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1130 net1200 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_2
Xfanout1141 net1143 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
X_10179_ datapath.PC\[9\] _03574_ datapath.PC\[10\] vssd1 vssd1 vccd1 vccd1 _05106_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__12440__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1152 net1164 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__clkbuf_4
Xfanout1163 net1164 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1174 net1175 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1185 net1199 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_2
Xfanout1196 net1198 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ clknet_leaf_33_clk _00825_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06868__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B2 _05517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ clknet_leaf_119_clk _00756_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08609__A1 _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07390_ datapath.rf.registers\[22\]\[20\] net753 net728 datapath.rf.registers\[2\]\[20\]
+ _02316_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08085__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ net638 _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__nor2_1
XANTENNA__07293__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08011_ datapath.rf.registers\[20\]\[6\] net900 net892 datapath.rf.registers\[14\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__a22o_1
XANTENNA__12615__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold602 datapath.rf.registers\[31\]\[21\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 datapath.rf.registers\[10\]\[18\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold624 datapath.rf.registers\[23\]\[17\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap343 _02016_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_4
Xhold635 datapath.rf.registers\[29\]\[29\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold646 datapath.rf.registers\[26\]\[28\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 datapath.rf.registers\[6\]\[20\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 datapath.rf.registers\[11\]\[29\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ datapath.PC\[28\] net539 vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__nor2_1
Xhold679 datapath.rf.registers\[24\]\[16\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
X_08913_ net412 _03472_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_139_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09893_ _04687_ _04689_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout296_A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12350__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _03766_ _03770_ net375 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
X_14568__1338 vssd1 vssd1 vccd1 vccd1 _14568__1338/HI net1338 sky130_fd_sc_hd__conb_1
XANTENNA__07899__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06849__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ _03639_ _03696_ _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _02644_ _02646_ _02652_ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__or3_2
XANTENNA_hold1209_A mmio.memload_or_instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06859__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07657_ datapath.rf.registers\[6\]\[14\] net813 net805 datapath.rf.registers\[15\]\[14\]
+ _02579_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout728_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ datapath.ru.latched_instruction\[29\] _01487_ _01508_ _01521_ vssd1 vssd1
+ vccd1 vccd1 _01538_ sky130_fd_sc_hd__a211o_1
XANTENNA__06584__A mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07588_ datapath.rf.registers\[8\]\[16\] net927 net871 datapath.rf.registers\[27\]\[16\]
+ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06539_ datapath.ru.latched_instruction\[14\] _01468_ vssd1 vssd1 vccd1 vccd1 _01469_
+ sky130_fd_sc_hd__nor2_1
X_09327_ net384 _03686_ _03524_ net393 vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__o211a_1
XANTENNA__08076__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ net492 _04182_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__nand2_1
XANTENNA__07823__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ datapath.rf.registers\[21\]\[2\] net937 net912 datapath.rf.registers\[18\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_153_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09189_ net670 _04084_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12525__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11220_ net1450 net145 net139 _04963_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__a22o_1
XANTENNA__07036__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14529__1351 vssd1 vssd1 vccd1 vccd1 net1351 _14529__1351/LO sky130_fd_sc_hd__conb_1
X_11151_ _05757_ _05759_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_56_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ net208 _05021_ net1312 vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a21oi_1
X_11082_ net1295 _05271_ _05677_ net1296 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_8_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__A0 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _04474_ _04955_ _04959_ net201 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__o211a_1
XANTENNA__12260__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__A2 _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ datapath.mulitply_result\[1\] datapath.multiplication_module.multiplicand_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13723_ clknet_leaf_94_clk datapath.multiplication_module.multiplier_i_n\[8\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[8\] sky130_fd_sc_hd__dfrtp_1
X_10935_ net269 net1914 net592 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ clknet_leaf_68_clk _00592_ net1224 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10866_ net271 net1667 net600 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ net1575 net296 net442 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XANTENNA__08067__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09264__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ clknet_leaf_87_clk _00535_ net1231 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10797_ _05487_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__or2_1
XANTENNA__10447__C _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07275__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12536_ net289 net1604 net448 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12467_ net164 net2384 net461 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07027__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ clknet_leaf_51_clk _01093_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11418_ screen.register.currentYbus\[28\] net133 _05894_ net162 vssd1 vssd1 vccd1
+ vccd1 _00386_ sky130_fd_sc_hd__a22o_1
X_12398_ net184 net1661 net469 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
XANTENNA__11374__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14137_ clknet_leaf_60_clk _01024_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11349_ _01459_ net1029 net309 net313 datapath.ru.latched_instruction\[28\] vssd1
+ vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ clknet_leaf_115_clk _00955_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07772__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ clknet_leaf_19_clk _00011_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ net1000 net983 net981 _01808_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__and4_4
XANTENNA__07264__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06819__D _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ _03485_ _03486_ net410 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__mux2_1
XANTENNA__08884__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ datapath.rf.registers\[7\]\[17\] _01740_ net778 datapath.rf.registers\[9\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11834__B1 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08491_ _02436_ _03417_ _02434_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07442_ net651 _02368_ net627 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07373_ net694 _02290_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__or3_1
XANTENNA__08058__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ _03506_ _04022_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__nor2_1
XANTENNA__07805__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09043_ _03412_ _03947_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12345__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout309_A _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07018__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 datapath.rf.registers\[12\]\[25\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold421 datapath.rf.registers\[19\]\[9\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 datapath.rf.registers\[29\]\[24\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 datapath.rf.registers\[13\]\[29\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold454 datapath.mulitply_result\[24\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1159_A mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 datapath.rf.registers\[9\]\[4\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 datapath.rf.registers\[12\]\[27\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1218_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 datapath.mulitply_result\[17\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 datapath.rf.registers\[18\]\[14\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 net902 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
Xfanout912 _01830_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_4
X_09945_ datapath.PC\[30\] _03591_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout923 _01826_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_4
XANTENNA_fanout580_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout945 net947 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__B _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net959 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_4
Xfanout967 _01805_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_4
X_09876_ _04751_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__xnor2_1
Xfanout978 _01663_ vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06579__A mmio.memload_or_instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1110 datapath.mulitply_result\[12\] vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net992 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_2
Xhold1121 datapath.rf.registers\[24\]\[9\] vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 datapath.rf.registers\[31\]\[28\] vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _03449_ _03753_ _03752_ _03750_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__o211a_1
Xhold1143 screen.register.currentXbus\[0\] vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 datapath.rf.registers\[21\]\[18\] vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 columns.count\[0\] vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 datapath.rf.registers\[27\]\[10\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 datapath.rf.registers\[18\]\[28\] vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net637 net334 _03684_ net656 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__o31a_1
Xhold1198 datapath.rf.registers\[30\]\[27\] vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07709_ datapath.rf.registers\[26\]\[13\] net940 _02635_ vssd1 vssd1 vccd1 vccd1
+ _02636_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08689_ _03476_ _03486_ _03456_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10720_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ datapath.mulitply_result\[20\] net427 net660 vssd1 vssd1 vccd1 vccd1 _05507_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07257__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ net1417 _02783_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[10\]
+ sky130_fd_sc_hd__mux2_1
X_13370_ clknet_leaf_90_clk _00355_ net1211 vssd1 vssd1 vccd1 vccd1 keypad.apps.app_c\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ net1821 net236 net476 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XANTENNA__07857__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12255__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07009__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net234 net2122 net487 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__mux2_1
X_11203_ net1476 net144 net137 _05048_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__a22o_1
X_12183_ columns.count\[5\] columns.count\[4\] _05849_ vssd1 vssd1 vccd1 vccd1 _06433_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ _05678_ _05713_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__or2_1
XANTENNA__11395__A _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ _05264_ _05701_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__or2_2
XANTENNA__10316__B1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09182__B1 _04107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ datapath.PC\[25\] net1312 _04941_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06639__D mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ net232 net2574 net581 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
XANTENNA__08288__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__B2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06936__B _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ clknet_leaf_56_clk datapath.multiplication_module.multiplicand_i_n\[23\]
+ net1256 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07496__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ net189 net2297 net596 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__mux2_1
XANTENNA__11292__B2 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net1477 _05883_ net156 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10458__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13637_ clknet_leaf_69_clk _00575_ net1228 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09237__A1 _02812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10849_ net1829 net190 net604 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07248__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ clknet_leaf_80_clk _00518_ net1234 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14567__1337 vssd1 vssd1 vccd1 vccd1 _14567__1337/HI net1337 sky130_fd_sc_hd__conb_1
XFILLER_0_143_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12519_ net1657 net236 net452 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__mux2_1
X_13499_ clknet_leaf_72_clk _00449_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.PC\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08460__A2 _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout208 _04665_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout219 _05519_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
X_07991_ datapath.rf.registers\[18\]\[7\] net789 net730 datapath.rf.registers\[16\]\[7\]
+ _02915_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ _04632_ _04655_ _04656_ _04654_ _04629_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a2111oi_1
X_06942_ datapath.rf.registers\[5\]\[30\] net784 net715 datapath.rf.registers\[29\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
X_09661_ _01952_ _03349_ _01910_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__o21ai_1
X_06873_ net652 _01799_ _01729_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a21o_1
XANTENNA__08920__A0 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ _03178_ net617 _03537_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ _02127_ _03343_ _02085_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o21ai_1
X_08543_ net506 net505 net404 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout161_A _05261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14528__1350 vssd1 vssd1 vccd1 vccd1 net1350 _14528__1350/LO sky130_fd_sc_hd__conb_1
XANTENNA__07487__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__B2 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _03383_ _03385_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07425_ datapath.rf.registers\[7\]\[19\] net825 net818 datapath.rf.registers\[31\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1070_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11256__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ datapath.rf.registers\[9\]\[21\] net886 net865 datapath.rf.registers\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a22o_1
X_07287_ _02192_ net528 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_150_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10794__B1 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _02431_ net354 _03892_ net390 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout795_A _01757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold240 datapath.rf.registers\[15\]\[24\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08203__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 datapath.rf.registers\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 datapath.rf.registers\[31\]\[24\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold273 datapath.rf.registers\[25\]\[7\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07411__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 datapath.PC\[9\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 datapath.rf.registers\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout962_A _01806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__A2 _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _01782_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_4
Xfanout731 net733 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
Xfanout742 net743 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_4
X_09928_ _04849_ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__nand2_1
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_4
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
Xfanout786 _01760_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_4
X_09859_ _04756_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nor2_1
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_29_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08911__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ net285 net2111 net549 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
XANTENNA__07190__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ datapath.PC\[16\] net303 _06221_ _06223_ vssd1 vssd1 vccd1 vccd1 _00460_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ net1327 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07478__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11752_ net1280 _06080_ net1019 vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11274__B2 mmio.memload_or_instruction\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10703_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__or2_1
XANTENNA__10993__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14471_ clknet_leaf_21_clk _01358_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11683_ net1623 _06128_ _06130_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_81_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ clknet_leaf_80_clk _00378_ net1233 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ net1275 _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08978__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13353_ clknet_leaf_95_clk _00338_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_10565_ _05413_ _05469_ _05423_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10785__A0 _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap1048 _05400_ vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_1
XFILLER_0_107_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12304_ net1550 net182 net477 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XANTENNA__07650__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13284_ clknet_leaf_60_clk _00274_ net1266 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10496_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ net182 net1565 net484 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__mux2_1
XANTENNA__12713__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__D1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _06418_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ _05717_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__nor2_1
XANTENNA__12014__A datapath.mulitply_result\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _06363_ _06364_ _06362_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10460__C _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ net1297 net1298 vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__nand2b_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07181__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12999_ net1479 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07469__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07210_ _02130_ _02132_ _02134_ _02136_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__or4_1
X_08190_ datapath.rf.registers\[6\]\[3\] net813 _03115_ _03116_ net831 vssd1 vssd1
+ vccd1 vccd1 _03117_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07141_ datapath.rf.registers\[26\]\[26\] net941 net897 datapath.rf.registers\[6\]\[26\]
+ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07072_ datapath.rf.registers\[30\]\[27\] net772 net761 datapath.rf.registers\[19\]\[27\]
+ _01998_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a221o_1
XANTENNA__08984__A3 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06995__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12623__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ datapath.rf.registers\[11\]\[7\] net968 net920 datapath.rf.registers\[2\]\[7\]
+ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a221o_1
X_09713_ _03250_ _03288_ _03308_ _03251_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__o31ai_1
X_06925_ datapath.rf.registers\[13\]\[31\] net865 net862 datapath.rf.registers\[28\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a22o_1
X_09644_ _03666_ _04570_ net411 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__mux2_1
X_06856_ net989 _01756_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__and2_2
XFILLER_0_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07172__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ _03427_ _04500_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_143_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ _01695_ _01713_ _01601_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_78_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__B _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ net504 _03446_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08457_ net514 _02833_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07408_ datapath.rf.registers\[23\]\[20\] net934 net894 datapath.rf.registers\[14\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a22o_1
XANTENNA__07880__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ net509 _03018_ _03067_ _03313_ _03063_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a221o_1
XANTENNA__10216__C1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07339_ datapath.rf.registers\[13\]\[21\] net793 net727 datapath.rf.registers\[2\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22o_1
XANTENNA__07200__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ net1292 screen.counter.ct\[8\] _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10231__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07632__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06986__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09009_ net337 _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__nor2_1
X_10281_ net670 _05185_ _05204_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__o22a_2
XANTENNA__12533__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12020_ datapath.mulitply_result\[7\] datapath.multiplication_module.multiplicand_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__nor2_1
Xfanout550 _06469_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
Xfanout561 _06466_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_8
Xfanout572 _06464_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
Xfanout583 _05675_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
X_13971_ clknet_leaf_59_clk _00858_ net1267 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10988__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 _05670_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_8
X_14566__1336 vssd1 vssd1 vccd1 vccd1 _14566__1336/HI net1336 sky130_fd_sc_hd__conb_1
X_12922_ net1918 net212 net547 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
XANTENNA__07699__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08360__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ net224 net1961 net554 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06910__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ net700 _04786_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__or2_1
XANTENNA__11247__B2 _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12784_ net243 net2492 net563 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14523_ net1314 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
X_11735_ screen.counter.ct\[13\] _06083_ _06078_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12708__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14454_ clknet_leaf_26_clk _01341_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11666_ screen.counter.currentCt\[9\] screen.counter.currentCt\[8\] _06114_ screen.counter.currentCt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a31o_1
XANTENNA__07871__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ clknet_leaf_89_clk _00361_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net1536 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[29\]
+ sky130_fd_sc_hd__and2_1
X_14385_ clknet_leaf_7_clk _01272_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11597_ net1017 _05723_ _05792_ _06060_ _05712_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__a32o_1
XANTENNA__12009__A datapath.mulitply_result\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13336_ clknet_leaf_94_clk _00321_ net1206 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_114_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07623__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ _05409_ _05456_ net1025 vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06977__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ clknet_leaf_91_clk _00257_ net1204 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12443__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ screen.register.currentYbus\[25\] screen.register.currentYbus\[24\] screen.register.currentYbus\[27\]
+ screen.register.currentYbus\[26\] vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_94_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12218_ net238 net1812 net576 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ clknet_leaf_1_clk _00190_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_102_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12149_ _06407_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__nand2_1
XANTENNA__09128__B1 _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10898__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ datapath.ru.latched_instruction\[22\] _01485_ net1027 vssd1 vssd1 vccd1 vccd1
+ _01637_ sky130_fd_sc_hd__mux2_1
X_07690_ datapath.rf.registers\[24\]\[13\] net755 net718 datapath.rf.registers\[28\]\[13\]
+ _02616_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a221o_1
XANTENNA__08887__C1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ _01564_ _01565_ _01567_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06827__D _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _04285_ _04286_ net370 vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21a_1
XANTENNA__11238__B2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06572_ net1305 net1303 mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01502_ sky130_fd_sc_hd__or3b_1
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11789__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ datapath.rf.registers\[22\]\[1\] net754 _03235_ _03236_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _03238_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09300__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09291_ net507 net353 _04217_ net384 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__a211o_1
XANTENNA__12618__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _03165_ _03166_ _03167_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_24 _01841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08173_ datapath.rf.registers\[31\]\[3\] net987 _01746_ vssd1 vssd1 vccd1 vccd1 _03100_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_144_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09603__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07124_ _02046_ _02048_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__or3_1
XANTENNA__06968__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07055_ datapath.rf.registers\[26\]\[28\] net941 net921 datapath.rf.registers\[2\]\[28\]
+ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a221o_1
XANTENNA__12353__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1033_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1200_A _00004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__inv_2
X_06908_ datapath.rf.registers\[24\]\[31\] net905 net901 datapath.rf.registers\[20\]\[31\]
+ _01832_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a221o_1
X_07888_ datapath.rf.registers\[5\]\[9\] net784 net752 datapath.rf.registers\[22\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a22o_1
XANTENNA__07145__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13884__RESET_B net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09627_ net335 _04056_ net315 vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a21o_1
X_06839_ net973 _01738_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout925_A _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09558_ _03449_ _04124_ _04482_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ _03361_ _03432_ _01995_ _03358_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09489_ net670 _04387_ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__o21ba_2
XANTENNA__12528__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ net1412 _05902_ _05988_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_61_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07853__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09410__B _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ screen.register.currentXbus\[1\] _05720_ _05735_ screen.register.currentYbus\[17\]
+ _05724_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a221o_1
X_10402_ net1290 net1288 vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__and2_1
XANTENNA__07605__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ clknet_leaf_22_clk _01057_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11382_ screen.register.currentYbus\[10\] net130 _05876_ net159 vssd1 vssd1 vccd1
+ vccd1 _00368_ sky130_fd_sc_hd__a22o_1
XANTENNA__09070__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06959__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ clknet_leaf_41_clk _00113_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10333_ _05168_ _05179_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__nor2_1
XANTENNA__12263__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ clknet_leaf_58_clk _00044_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10264_ _03888_ _05190_ net331 vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__mux2_1
X_12003_ _06281_ _06283_ _06280_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__o21ba_1
Xfanout1301 screen.counter.ct\[0\] vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08030__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _04665_ _05121_ net1310 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__a21o_1
Xfanout1312 _01451_ vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__buf_2
XANTENNA__07384__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06592__B1 _01464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_2
X_13954_ clknet_leaf_33_clk _00841_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07136__A2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ net1810 net279 net545 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
X_13885_ clknet_leaf_32_clk _00772_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ net295 net2264 net554 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12438__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ net288 net2449 net562 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__mux2_1
XANTENNA__08636__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ clknet_leaf_9_clk _01393_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07844__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ net1294 _06068_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12698_ net2085 net163 net433 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__mux2_1
XANTENNA__10466__B _03087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14437_ clknet_leaf_94_clk _01324_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11649_ screen.counter.currentCt\[3\] screen.counter.currentCt\[4\] _06104_ vssd1
+ vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__and3_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09597__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14368_ clknet_leaf_46_clk _01255_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold806 datapath.rf.registers\[28\]\[0\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 datapath.rf.registers\[20\]\[6\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold828 datapath.rf.registers\[5\]\[10\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_112_clk _00309_ net1098 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold839 datapath.rf.registers\[26\]\[27\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14299_ clknet_leaf_54_clk _01186_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08021__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _02349_ _03335_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12901__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _02732_ _02733_ _02735_ _02737_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__or4_1
X_08791_ net371 _03710_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_127_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07742_ _02667_ _02668_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__or2_1
XANTENNA__08324__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ _02591_ _02593_ _02598_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_140_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ _02932_ _03317_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_140_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06624_ datapath.ru.latched_instruction\[28\] datapath.ru.latched_instruction\[29\]
+ datapath.ru.latched_instruction\[30\] datapath.ru.latched_instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__or4_1
XANTENNA__08088__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ net639 _04252_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand2_1
X_06555_ mmio.memload_or_instruction\[22\] net1061 vssd1 vssd1 vccd1 vccd1 _01485_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12348__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ _04087_ _04088_ net365 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__a21o_1
X_06486_ datapath.ru.latched_instruction\[22\] vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ datapath.rf.registers\[29\]\[2\] net989 _01756_ vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_105_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1189_A mmio.memload_or_instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout506_A _03087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ datapath.rf.registers\[8\]\[3\] net925 net913 datapath.rf.registers\[18\]\[3\]
+ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__a221o_1
X_14565__1335 vssd1 vssd1 vccd1 vccd1 _14565__1335/HI net1335 sky130_fd_sc_hd__conb_1
XFILLER_0_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07107_ datapath.rf.registers\[16\]\[27\] net963 net874 datapath.rf.registers\[25\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a22o_1
XANTENNA__08260__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ datapath.rf.registers\[24\]\[5\] net755 net751 datapath.rf.registers\[22\]\[5\]
+ _03001_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__a221o_1
X_07038_ _01958_ _01960_ _01962_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__or4_1
XANTENNA__08012__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12811__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net656 net637 _03552_ net610 vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07118__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06586__C_N mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ net197 net2395 net593 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10122__A1 _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ clknet_leaf_78_clk net1394 net1233 vssd1 vssd1 vccd1 vccd1 datapath.pc_module.i_ack2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11870__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10882_ net197 net2030 net601 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__mux2_1
X_12621_ net1837 net230 net442 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__mux2_1
XANTENNA__08079__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12258__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12552_ net236 net1819 net448 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
XANTENNA__07826__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ net1440 _05902_ _05972_ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__a21o_1
X_12483_ net252 net1875 net457 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ clknet_leaf_118_clk _01109_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11434_ screen.register.currentXbus\[8\] net1016 _05906_ vssd1 vssd1 vccd1 vccd1
+ _05907_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_78_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14153_ clknet_leaf_13_clk _01040_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07595__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11365_ _03148_ _03175_ net669 vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_100_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13104_ clknet_leaf_0_clk _00096_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10316_ _05169_ _05238_ _05241_ net1309 net1278 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a32o_1
X_14084_ clknet_leaf_16_clk _00971_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11296_ net17 net1044 net1033 mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1
+ vccd1 _00310_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_91_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ clknet_leaf_55_clk _00027_ net1175 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12721__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10247_ datapath.PC\[3\] net1055 _04935_ _05171_ vssd1 vssd1 vccd1 vccd1 _05174_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07357__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_4
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_4
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_2
X_10178_ _01427_ _04416_ net537 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__mux2_1
Xfanout1153 net1164 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_2
Xfanout1164 net1200 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1175 net1180 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1186 net1187 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_4
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_2
XANTENNA__11310__A0 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13937_ clknet_leaf_8_clk _00824_ net1084 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13868_ clknet_leaf_30_clk _00755_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12819_ net230 net2049 net558 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__mux2_1
X_13799_ clknet_leaf_18_clk _00686_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ datapath.rf.registers\[29\]\[6\] net876 net864 datapath.rf.registers\[13\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11916__A2 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 datapath.rf.registers\[29\]\[1\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold614 datapath.rf.registers\[26\]\[12\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 datapath.mulitply_result\[22\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold636 datapath.rf.registers\[19\]\[5\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 datapath.rf.registers\[8\]\[19\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 datapath.rf.registers\[4\]\[10\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _04886_ _04887_ datapath.PC\[29\] net1313 vssd1 vssd1 vccd1 vccd1 _04888_
+ sky130_fd_sc_hd__a2bb2o_1
Xhold669 datapath.rf.registers\[15\]\[19\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ _03499_ _03832_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a21bo_1
X_09892_ _04762_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__nor2_1
XANTENNA__12631__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ net367 _03768_ _03769_ _03767_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout191_A _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06849__B net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ _03695_ _03697_ _03700_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07725_ _02636_ _02647_ _02649_ _02651_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11771__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1198_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ datapath.rf.registers\[5\]\[14\] net782 net778 datapath.rf.registers\[9\]\[14\]
+ _02575_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a221o_1
XANTENNA__07520__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06607_ datapath.ru.latched_instruction\[28\] _01460_ _01509_ _01413_ _01536_ vssd1
+ vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ datapath.rf.registers\[20\]\[16\] net902 net879 datapath.rf.registers\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a22o_1
X_09326_ net634 _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__nor2_1
XANTENNA__07808__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06538_ net1307 net1304 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ _01468_ sky130_fd_sc_hd__or3b_2
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ net639 _04156_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12806__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08208_ datapath.rf.registers\[31\]\[2\] net951 net920 datapath.rf.registers\[2\]\[2\]
+ _03134_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_153_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09188_ _04086_ _04112_ _04114_ net675 vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08233__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ net507 _03062_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08304__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07587__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ net1279 screen.counter.ct\[22\] _05760_ net1280 vssd1 vssd1 vccd1 vccd1 _05800_
+ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_56_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10591__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10101_ net704 _04499_ _05027_ _05026_ net208 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a311o_1
XANTENNA__12541__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ net1297 net1299 _05718_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_8_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07339__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09733__A0 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ net1052 _04956_ _04958_ net704 vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a211o_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ datapath.multiplication_module.multiplier_i\[0\] net346 vssd1 vssd1 vccd1
+ vccd1 _06270_ sky130_fd_sc_hd__and2_1
XANTENNA__10996__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[7\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ net274 net2456 net591 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07511__A2 _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09151__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ clknet_leaf_68_clk _00591_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10865_ net275 net2027 net599 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__mux2_1
XANTENNA__10297__A _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12604_ net1696 net292 net443 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
X_13584_ clknet_leaf_79_clk _00534_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10796_ datapath.PC\[11\] _05486_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10447__D _02721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12535_ net182 net1523 net448 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12716__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ net170 net2289 net462 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__mux2_1
X_14205_ clknet_leaf_31_clk _01092_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11417_ net425 net714 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12397_ net190 net2043 net470 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__mux2_1
XANTENNA__07578__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output85_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ clknet_leaf_40_clk _01023_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11348_ _01512_ net1027 net308 net312 datapath.ru.latched_instruction\[27\] vssd1
+ vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__a32o_1
XANTENNA__10582__A1 _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ clknet_leaf_49_clk _00954_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12451__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ net30 net1045 net1034 mmio.memload_or_instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _00293_ sky130_fd_sc_hd__o22a_1
XANTENNA__08527__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__D1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ clknet_leaf_23_clk _00010_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14564__1334 vssd1 vssd1 vccd1 vccd1 _14564__1334/HI net1334 sky130_fd_sc_hd__conb_1
XFILLER_0_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _02435_ _02436_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__nor2_2
XANTENNA__10637__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08490_ _03415_ _03416_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__or2_1
XANTENNA__07502__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ datapath.rf.registers\[0\]\[19\] net828 _02358_ _02367_ vssd1 vssd1 vccd1
+ vccd1 _02368_ sky130_fd_sc_hd__o22a_4
XFILLER_0_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ _02292_ _02294_ _02296_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09111_ net319 _04035_ _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12626__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10270__A0 _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ net638 _03968_ _03959_ net655 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08215__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 datapath.rf.registers\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 datapath.rf.registers\[11\]\[8\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 datapath.rf.registers\[5\]\[14\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 datapath.rf.registers\[5\]\[31\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 datapath.rf.registers\[22\]\[7\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 datapath.rf.registers\[4\]\[17\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A1 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 datapath.rf.registers\[14\]\[9\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 datapath.mulitply_result\[16\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11766__A _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_4
X_09944_ net538 _04587_ _04607_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a31o_1
Xhold488 datapath.rf.registers\[21\]\[15\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 datapath.rf.registers\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 _01830_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_2
XANTENNA__12361__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 _01825_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 _01819_ vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _04716_ _04718_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__nor2_1
Xfanout957 net959 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_4
Xfanout968 _01802_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_4
Xhold1100 datapath.rf.registers\[14\]\[16\] vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__B1 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 _01663_ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1111 datapath.rf.registers\[2\]\[27\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 datapath.rf.registers\[17\]\[23\] vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net416 _03606_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__nand2_1
Xhold1133 datapath.rf.registers\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 datapath.rf.registers\[9\]\[18\] vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 datapath.rf.registers\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 datapath.rf.registers\[13\]\[16\] vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net369 _03676_ _03683_ net376 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__a211o_1
Xhold1177 datapath.rf.registers\[1\]\[28\] vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 datapath.rf.registers\[20\]\[31\] vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 datapath.rf.registers\[15\]\[10\] vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
X_07708_ datapath.rf.registers\[16\]\[13\] net960 net924 datapath.rf.registers\[8\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22o_1
X_08688_ _03485_ _03488_ net341 vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07639_ datapath.rf.registers\[0\]\[15\] net692 _02553_ _02565_ vssd1 vssd1 vccd1
+ vccd1 _02566_ sky130_fd_sc_hd__o22a_4
XFILLER_0_137_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _03831_ _05505_ net845 vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09309_ _04233_ _04234_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__and3_1
X_10581_ net1410 _02831_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[9\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12536__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ net1682 net240 net479 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XANTENNA__10800__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net238 net2061 net486 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__mux2_1
X_11202_ net1573 net143 net138 _05180_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__a22o_1
XANTENNA__09954__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net1442 _06432_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11133_ _05780_ _05781_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__nor2_1
XANTENNA__12271__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ _05264_ _05701_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
XANTENNA__11395__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__B1 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09182__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09182__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net201 _04836_ _04933_ net1268 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__o31a_1
XANTENNA__07193__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06940__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output123_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11966_ net228 net1845 net580 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13705_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[22\]
+ net1256 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10917_ net193 net2195 net596 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__mux2_1
X_11897_ net1478 _05882_ net156 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__mux2_1
XANTENNA__10458__C net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13636_ clknet_leaf_51_clk _00574_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07113__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10848_ net2054 net194 net603 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12446__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ clknet_leaf_86_clk _00517_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10779_ _05485_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nor2_1
XANTENNA__07799__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12518_ net1605 net238 net453 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13498_ clknet_leaf_73_clk _00448_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.PC\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08460__A3 _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ net255 net2069 net460 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14119_ clknet_leaf_21_clk _01006_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10490__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ datapath.rf.registers\[3\]\[7\] net766 net740 datapath.rf.registers\[1\]\[7\]
+ _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a221o_1
Xfanout209 _05531_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_130_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07971__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__A_N net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ datapath.rf.registers\[18\]\[30\] net790 net753 datapath.rf.registers\[22\]\[30\]
+ _01866_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a221o_1
XANTENNA__10307__A1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ _03558_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__or2_1
X_06872_ datapath.rf.registers\[0\]\[31\] _01798_ net828 vssd1 vssd1 vccd1 vccd1 _01799_
+ sky130_fd_sc_hd__mux2_8
XANTENNA__07184__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ net504 net618 _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08920__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ net676 _04513_ _04516_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__o31a_1
X_08542_ _03467_ _03468_ net408 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__mux2_1
XANTENNA__06846__C _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ _02882_ _03399_ _02883_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__a21o_1
X_07424_ datapath.rf.registers\[25\]\[19\] net797 net715 datapath.rf.registers\[29\]\[19\]
+ _02350_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07355_ net648 net342 _01730_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12356__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1063_A _01455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07286_ _02192_ net528 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06998__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09025_ _02520_ net354 _03950_ net386 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1230_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 datapath.rf.registers\[3\]\[25\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 datapath.rf.registers\[17\]\[2\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 datapath.rf.registers\[13\]\[28\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 datapath.rf.registers\[13\]\[15\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold274 datapath.rf.registers\[12\]\[28\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 datapath.rf.registers\[7\]\[5\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold296 datapath.rf.registers\[3\]\[30\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_4
Xfanout721 _01782_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
X_09927_ _04850_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__xnor2_1
Xfanout743 _01774_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_2
Xfanout754 _01771_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout765 _01767_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_4
X_09858_ _04712_ _04755_ _04708_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a21oi_1
Xfanout787 _01760_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_4
Xfanout798 _01755_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_4
XANTENNA__07714__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ net416 _03473_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__and2_1
X_09789_ net1277 _02832_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__nor2_1
XANTENNA__06922__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ _05657_ net176 _06222_ net178 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ net1764 net664 _06171_ net713 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__a22o_1
XANTENNA__11274__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_80_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10702_ datapath.PC\[27\] _05538_ datapath.PC\[28\] vssd1 vssd1 vccd1 vccd1 _05550_
+ sky130_fd_sc_hd__a21oi_1
X_14470_ clknet_leaf_114_clk _01357_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11682_ screen.counter.currentCt\[15\] _06128_ _06088_ vssd1 vssd1 vccd1 vccd1 _06130_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13421_ clknet_leaf_89_clk _00377_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ datapath.PC\[17\] _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12266__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08978__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ clknet_leaf_71_clk _00337_ net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ _05460_ _05469_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap1049 _05398_ vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06989__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ net577 _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__nor2_4
XFILLER_0_122_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13283_ clknet_leaf_60_clk _00273_ net1266 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
X_10495_ net122 net123 net124 net121 vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__or4b_2
X_12234_ _05666_ _06443_ net577 vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__or3_1
XANTENNA__07884__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12165_ net323 _06421_ _06422_ net327 net1939 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_112_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ _05269_ _05270_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__or3_1
X_12096_ _06362_ _06363_ _06364_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__or3_1
XANTENNA__10460__D _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ net1296 net1295 _05271_ _05677_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__or4_1
XANTENNA__07166__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06913__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12998_ net2345 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11949_ net298 net1553 net579 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08130__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13619_ clknet_leaf_8_clk _00557_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ datapath.rf.registers\[15\]\[26\] net858 net849 datapath.rf.registers\[1\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07071_ datapath.rf.registers\[26\]\[27\] net822 net791 datapath.rf.registers\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_33_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12904__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07944__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ datapath.rf.registers\[20\]\[7\] net900 net888 datapath.rf.registers\[12\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a22o_1
X_09712_ _02436_ _03372_ _03415_ _04638_ _03371_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a221o_1
X_06924_ net999 net985 net980 _01812_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and4_4
X_09643_ _04526_ _04569_ _03456_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__mux2_1
X_06855_ net988 _01776_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__and2_2
X_09574_ _03342_ _04500_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__xnor2_1
X_06786_ datapath.ru.latched_instruction\[8\] _01668_ _01697_ _01700_ _01712_ vssd1
+ vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_143_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _01638_ _03446_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08456_ _02833_ net514 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__nand2b_1
X_07407_ datapath.rf.registers\[31\]\[20\] net950 net906 datapath.rf.registers\[24\]\[20\]
+ _02333_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ _03067_ _03313_ _03063_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout703_A _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07338_ datapath.rf.registers\[26\]\[21\] net821 net797 datapath.rf.registers\[25\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ datapath.rf.registers\[2\]\[23\] net922 net862 datapath.rf.registers\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a22o_1
XANTENNA__12814__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ _03692_ _03934_ net402 vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__mux2_1
X_10280_ net655 _01633_ net641 _05185_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__a41o_1
XFILLER_0_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08188__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _01714_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
Xfanout551 _06469_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_8
Xfanout562 _06466_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
Xfanout573 _06446_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_6
X_13970_ clknet_leaf_35_clk _00857_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07148__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout584 _05675_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_8
Xfanout595 _05670_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_4
X_12921_ net2047 net215 net546 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
XANTENNA__08360__A2 _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ net230 net2298 net555 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11803_ net701 _04046_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12783_ net237 net2067 net561 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__mux2_1
XANTENNA__11247__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_53_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
X_11734_ net1291 net664 _06161_ net713 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__a22o_1
X_14522_ net1348 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11665_ net1489 _06116_ _06118_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a21oi_1
X_14453_ clknet_leaf_27_clk _01340_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ clknet_leaf_89_clk _00360_ net1231 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10616_ net1554 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[28\]
+ sky130_fd_sc_hd__and2_1
X_14384_ clknet_leaf_4_clk _01271_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ _05323_ _06053_ _06059_ _05294_ _06052_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13335_ clknet_leaf_93_clk _00320_ net1205 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_4
X_10547_ _05413_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12724__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ clknet_leaf_109_clk _00256_ net1107 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10478_ screen.register.currentYbus\[29\] screen.register.currentYbus\[28\] screen.register.currentYbus\[31\]
+ screen.register.currentYbus\[30\] vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__or4_1
XANTENNA__08179__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ net245 net2501 net575 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13197_ clknet_leaf_119_clk _00189_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11567__C _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07387__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ datapath.mulitply_result\[28\] datapath.multiplication_module.multiplicand_i\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__or2_1
XANTENNA__09128__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11255__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ _06342_ _06349_ _06348_ _06347_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__o211ai_1
XANTENNA__11486__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08351__A2 _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ _01457_ _01458_ _01477_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10694__B1 _05542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06571_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nand2_2
XANTENNA__11238__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_08310_ datapath.rf.registers\[2\]\[1\] net974 _01741_ vssd1 vssd1 vccd1 vccd1 _03237_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08103__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ net499 net622 net490 net506 vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07311__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ datapath.rf.registers\[9\]\[2\] net778 net773 datapath.rf.registers\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_14 mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_25 _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_36 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08172_ datapath.rf.registers\[4\]\[3\] net993 _01734_ vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10749__A1 _01456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ datapath.rf.registers\[3\]\[26\] net767 net723 datapath.rf.registers\[27\]\[26\]
+ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12634__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ datapath.rf.registers\[31\]\[28\] net949 net930 datapath.rf.registers\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a22o_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XFILLER_0_88_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_3_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07378__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _02879_ net513 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_145_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06907_ net1000 net985 net980 _01808_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__and4_1
X_07887_ datapath.rf.registers\[7\]\[9\] net825 net741 datapath.rf.registers\[1\]\[9\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout653_A _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06838_ net987 _01752_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__and2_1
X_09626_ net332 net377 _03844_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_39_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ _02256_ net686 net678 _02260_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__o221a_1
XANTENNA__11229__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06769_ datapath.ru.latched_instruction\[0\] _01586_ _01612_ datapath.ru.latched_instruction\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__a22o_1
XANTENNA__12809__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
X_08508_ _01994_ _03358_ _03360_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__a21o_1
X_09488_ net670 _04410_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__and3_1
XANTENNA__07302__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ _02193_ _02212_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11450_ screen.register.currentXbus\[25\] net1013 _05742_ screen.register.currentYbus\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11937__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10401_ screen.controlBus\[6\] _05277_ _05293_ screen.controlBus\[7\] vssd1 vssd1
+ vccd1 vccd1 _05323_ sky130_fd_sc_hd__and4bb_2
X_11381_ _02783_ net668 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__and2_1
XANTENNA__12544__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13120_ clknet_leaf_46_clk _00112_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10332_ _05168_ _05180_ _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__or3b_1
XANTENNA__07081__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ clknet_leaf_19_clk _00043_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09138__B _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ net382 _04092_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07369__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12002_ datapath.mulitply_result\[4\] datapath.multiplication_module.multiplicand_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nor2_1
Xfanout1302 net1304 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__buf_2
XANTENNA__10999__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _04809_ _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__nand2_1
Xfanout1313 _01451_ vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout370 _03539_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_2
Xfanout381 net383 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_2
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_2
XANTENNA__10125__C1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13953_ clknet_leaf_42_clk _00840_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12904_ net2127 _05607_ net545 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
X_13884_ clknet_leaf_57_clk _00771_ net1261 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08993__A _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ net292 net1823 net556 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
XANTENNA__06895__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12719__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12766_ net180 net1833 net562 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14505_ clknet_leaf_13_clk _01392_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11717_ net1422 net663 _06151_ net712 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__a22o_1
X_12697_ net1762 net168 net433 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10466__C _03146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ _06106_ _06107_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__nor2_1
X_14436_ clknet_leaf_14_clk _01323_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11928__B1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11579_ net1017 _05723_ _05790_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__a31o_1
XANTENNA__12454__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ clknet_leaf_39_clk _01254_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold807 datapath.rf.registers\[9\]\[15\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_110_clk _00308_ net1104 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold818 datapath.rf.registers\[5\]\[18\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold829 datapath.rf.registers\[27\]\[26\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_23_clk _01185_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09349__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13249_ clknet_leaf_65_clk _00239_ net1269 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ datapath.rf.registers\[3\]\[11\] net964 net944 datapath.rf.registers\[19\]\[11\]
+ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a221o_1
XANTENNA__11594__A _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ net375 _03715_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__and3_1
XANTENNA__14311__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07780__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ datapath.rf.registers\[5\]\[12\] net782 net765 datapath.rf.registers\[17\]\[12\]
+ _02665_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a221o_1
XANTENNA__08324__A2 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07672_ datapath.rf.registers\[20\]\[14\] net900 net880 datapath.rf.registers\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
XANTENNA__07532__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ _04192_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_140_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06623_ datapath.ru.latched_instruction\[16\] datapath.ru.latched_instruction\[17\]
+ datapath.ru.latched_instruction\[18\] datapath.ru.latched_instruction\[19\] vssd1
+ vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12629__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ _04253_ _04268_ net616 _04236_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__o211ai_2
X_06554_ net1307 net1304 mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ _01484_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ _04198_ _04199_ net361 vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__a21o_1
X_06485_ datapath.ru.latched_instruction\[20\] vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08224_ datapath.rf.registers\[3\]\[2\] net973 _01738_ vssd1 vssd1 vccd1 vccd1 _03151_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11919__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ datapath.rf.registers\[31\]\[3\] net951 net875 datapath.rf.registers\[25\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__a22o_1
XANTENNA__12364__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ datapath.rf.registers\[27\]\[27\] net870 net862 datapath.rf.registers\[28\]\[27\]
+ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a221o_1
X_08086_ datapath.rf.registers\[8\]\[5\] net737 _03010_ _03011_ _03012_ vssd1 vssd1
+ vccd1 vccd1 _03013_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_12_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07037_ datapath.rf.registers\[4\]\[28\] net810 net763 datapath.rf.registers\[17\]\[28\]
+ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_58_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout770_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A _01848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ _03329_ _03914_ _03912_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a21oi_1
X_07939_ datapath.rf.registers\[19\]\[8\] net762 net716 datapath.rf.registers\[29\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a22o_1
XANTENNA__08315__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10950_ net209 net2375 net593 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09609_ _03344_ _04519_ _03556_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__a21o_1
X_10881_ net210 net2179 net601 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__mux2_1
XANTENNA__12539__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ net1770 net228 net441 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__mux2_1
XANTENNA__09276__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ net239 net2333 net450 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net975 _05808_ _05815_ _05901_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__o311a_1
XFILLER_0_109_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12482_ net254 net2385 net456 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11433_ screen.register.currentXbus\[16\] net1015 _05742_ screen.register.currentYbus\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a22o_1
X_14221_ clknet_leaf_119_clk _01108_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12274__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11386__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ clknet_leaf_13_clk _01039_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07054__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ screen.register.currentYbus\[1\] net130 _05867_ net159 vssd1 vssd1 vccd1
+ vccd1 _00359_ sky130_fd_sc_hd__a22o_1
X_13103_ clknet_leaf_5_clk _00095_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10315_ _05169_ _05238_ _05241_ net1309 datapath.PC\[2\] vssd1 vssd1 vccd1 vccd1
+ _05242_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_132_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14083_ clknet_leaf_103_clk _00970_ net1121 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11295_ net16 net1045 net1034 mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1
+ vccd1 _00309_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ clknet_leaf_9_clk _00026_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ _05169_ _05172_ _04232_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a21oi_1
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_2
Xfanout1121 net1124 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_2
Xfanout1132 net1135 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_4
X_10177_ _04386_ _04416_ net700 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__o21a_1
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07762__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1154 net1163 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_4
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1176 net1180 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1187 net1199 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_2
Xfanout1198 net1199 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_2
X_13936_ clknet_leaf_4_clk _00823_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07514__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12449__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ clknet_leaf_101_clk _00754_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12818_ net227 net1768 net558 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ clknet_leaf_111_clk _00685_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12749_ net238 net1937 net568 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07293__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14419_ clknet_leaf_49_clk _01306_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold604 datapath.rf.registers\[26\]\[18\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 datapath.rf.registers\[8\]\[8\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 datapath.rf.registers\[15\]\[3\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 datapath.rf.registers\[13\]\[2\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold648 net68 vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12912__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09960_ net207 _04855_ _04883_ net1313 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a31o_1
Xhold659 datapath.rf.registers\[7\]\[30\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_08911_ _02391_ net685 net681 _02390_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o22a_1
X_09891_ _04696_ _04761_ _04693_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a21oi_1
X_08842_ _03542_ _03544_ net526 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a21o_1
XANTENNA__07753__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06849__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ net615 _03669_ _03699_ net676 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a31o_1
X_07724_ datapath.rf.registers\[19\]\[13\] net944 net904 datapath.rf.registers\[24\]\[13\]
+ _02650_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11301__B2 mmio.memload_or_instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ datapath.rf.registers\[11\]\[14\] net774 _02574_ _02581_ vssd1 vssd1 vccd1
+ vccd1 _02582_ sky130_fd_sc_hd__a211o_1
XANTENNA__06859__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ datapath.ru.latched_instruction\[26\] _01466_ _01489_ datapath.ru.latched_instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout449_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ datapath.rf.registers\[17\]\[16\] net882 net854 datapath.rf.registers\[5\]\[16\]
+ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a221o_1
XANTENNA__08138__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ _04241_ _04245_ _04251_ net332 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__a22o_1
X_06537_ datapath.ru.latched_instruction\[26\] _01466_ vssd1 vssd1 vccd1 vccd1 _01467_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1260_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _04117_ _04182_ net688 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XANTENNA__07284__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08207_ datapath.rf.registers\[20\]\[2\] net900 net892 datapath.rf.registers\[14\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ net616 _04110_ _04113_ net492 _04083_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_153_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ net507 _03062_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__nand2_1
XANTENNA__07036__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__B1 _04353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _02991_ _02993_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12822__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _03703_ _04498_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_73_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ net1013 vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _03583_ _04957_ net1052 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07744__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ datapath.multiplication_module.multiplier_i\[0\] net350 vssd1 vssd1 vccd1
+ vccd1 _06269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13721_ clknet_leaf_88_clk datapath.multiplication_module.multiplier_i_n\[6\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[6\] sky130_fd_sc_hd__dfrtp_1
X_10933_ net277 net2133 net590 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__mux2_1
XANTENNA__12269__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09151__B _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net277 net1626 net598 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__mux2_1
X_13652_ clknet_leaf_68_clk _00590_ net1223 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08048__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ net2003 net299 net443 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13583_ clknet_leaf_80_clk _00533_ net1233 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10795_ net2369 net265 net602 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ _05479_ _05669_ net577 vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__or3_1
XANTENNA__07275__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ net171 net2299 net463 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14204_ clknet_leaf_53_clk _01091_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07027__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ screen.register.currentYbus\[27\] net131 _05893_ net160 vssd1 vssd1 vccd1
+ vccd1 _00385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12396_ net195 net2098 net469 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
X_11347_ mmio.memload_or_instruction\[26\] net1063 net310 net314 datapath.ru.latched_instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a32o_1
X_14135_ clknet_leaf_44_clk _01022_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07983__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ net29 net1046 net1035 mmio.memload_or_instruction\[5\] vssd1 vssd1 vccd1
+ vccd1 _00292_ sky130_fd_sc_hd__a22o_1
X_14066_ clknet_leaf_35_clk _00953_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09185__C1 _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _04814_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__nand2_1
X_13017_ clknet_leaf_60_clk _00009_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09326__B _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 mmio.WEN1 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11295__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13919_ clknet_leaf_37_clk _00806_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10488__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07440_ _02360_ _02362_ _02364_ _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07371_ datapath.rf.registers\[21\]\[21\] net938 net893 datapath.rf.registers\[14\]\[21\]
+ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12907__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ _02699_ net687 net679 _02702_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ net329 net377 _03547_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__o31a_1
XANTENNA__10270__A1 _03146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07018__A2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 datapath.rf.registers\[30\]\[18\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 datapath.rf.registers\[17\]\[24\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 net75 vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 datapath.rf.registers\[25\]\[5\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 datapath.rf.registers\[8\]\[17\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12642__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold456 datapath.rf.registers\[7\]\[11\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06777__A1 datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold467 datapath.rf.registers\[18\]\[0\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 datapath.rf.registers\[27\]\[2\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 datapath.rf.registers\[30\]\[11\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ datapath.PC\[30\] net538 net1053 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout903 _01834_ vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 _01830_ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_4
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout925 _01825_ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout936 _01817_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_4
Xfanout947 _01814_ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nor2_1
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
Xhold1101 datapath.rf.registers\[7\]\[13\] vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 _01802_ vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
Xhold1112 datapath.rf.registers\[2\]\[28\] vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 datapath.rf.registers\[1\]\[10\] vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _02302_ net685 net681 _02304_ _03751_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__o221a_1
Xhold1134 datapath.rf.registers\[26\]\[29\] vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 datapath.rf.registers\[20\]\[28\] vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _06465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 datapath.rf.registers\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 datapath.rf.registers\[18\]\[13\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 datapath.rf.registers\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ net371 _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__nor2_1
Xhold1189 mmio.memload_or_instruction\[20\] vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
X_07707_ net650 _02633_ net627 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a21o_1
XANTENNA__11825__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ net411 _03612_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08151__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ net694 _02555_ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout900_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ datapath.rf.registers\[4\]\[16\] net811 net742 datapath.rf.registers\[1\]\[16\]
+ _02495_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__a221o_1
XANTENNA__12817__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11589__A1 _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _03179_ _03494_ net680 _03182_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__a22oi_1
X_10580_ net1506 _02876_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[8\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07257__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ net512 net357 _04165_ net385 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ net245 net2087 net485 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__mux2_1
XANTENNA__07009__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ net1494 net144 net138 _05243_ vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__a22o_1
XANTENNA__11210__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__A1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _05851_ _06431_ _06432_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__and3b_1
XFILLER_0_102_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12552__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07965__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ _05715_ net1021 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__or2_1
Xhold990 datapath.rf.registers\[8\]\[2\] vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11063_ net1297 net1298 _05702_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__or3_1
XANTENNA__09146__B _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08050__B _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07717__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _04499_ _04940_ _04939_ _04934_ net206 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08390__B1 _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ net244 net1982 net580 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08142__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09485__A3 _04408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13704_ clknet_leaf_68_clk datapath.multiplication_module.multiplicand_i_n\[21\]
+ net1258 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10916_ net198 net2278 net597 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__mux2_1
XANTENNA__07496__A2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net1429 _05881_ net158 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10458__D _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13635_ clknet_leaf_44_clk _00573_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net1597 net199 net604 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__mux2_1
XANTENNA__12727__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07248__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09642__A0 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ clknet_leaf_86_clk _00516_ net1234 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10778_ datapath.PC\[8\] _05484_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12517_ net2429 net245 net454 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__mux2_1
X_13497_ clknet_leaf_73_clk _00447_ net1243 vssd1 vssd1 vccd1 vccd1 datapath.PC\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12448_ net258 net2255 net460 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11201__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12462__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12379_ net271 net1738 net469 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
X_14118_ clknet_leaf_105_clk _01005_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10490__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06940_ datapath.rf.registers\[11\]\[30\] net775 net720 datapath.rf.registers\[28\]\[30\]
+ _01865_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a221o_1
X_14049_ clknet_leaf_42_clk _00936_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07708__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06871_ datapath.rf.registers\[11\]\[31\] net775 _01795_ _01796_ _01797_ vssd1 vssd1
+ vccd1 vccd1 _01798_ sky130_fd_sc_hd__a2111o_1
XANTENNA_max_cap998_A _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _01638_ net617 vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__nor2_1
X_09590_ net677 _04502_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09072__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11268__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ _02997_ net508 net404 vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__mux2_1
X_08472_ _02931_ _03398_ _02930_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07487__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07423_ datapath.rf.registers\[4\]\[19\] net810 net802 datapath.rf.registers\[20\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12637__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07354_ net648 net342 net626 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07285_ datapath.rf.registers\[0\]\[23\] net692 _02199_ _02211_ vssd1 vssd1 vccd1
+ vccd1 _02212_ sky130_fd_sc_hd__o22a_2
XFILLER_0_143_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout314_A _05859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1056_A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ _02520_ net354 _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_150_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold220 datapath.rf.registers\[19\]\[1\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12372__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 datapath.rf.registers\[25\]\[25\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1223_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 datapath.rf.registers\[25\]\[28\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 datapath.rf.registers\[4\]\[2\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 datapath.rf.registers\[15\]\[8\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07411__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 datapath.rf.registers\[27\]\[16\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 net703 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_2
Xhold286 datapath.rf.registers\[12\]\[15\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 datapath.rf.registers\[16\]\[2\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout711 _01603_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_2
Xfanout722 net725 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
X_09926_ _04851_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__nand2b_1
Xfanout733 _01778_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 _01773_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_4
Xfanout755 net758 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_4
Xfanout766 net769 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_8
Xfanout777 _01764_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_4
X_09857_ _04685_ _04765_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 _01760_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_4
Xfanout799 _01753_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout948_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _02213_ net686 net682 _02214_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__o22ai_2
X_09788_ _04713_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11259__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ _03664_ _03665_ net409 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__mux2_1
XANTENNA__08124__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _06080_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__nor2_1
XANTENNA__07478__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ datapath.PC\[27\] datapath.PC\[28\] _05538_ vssd1 vssd1 vccd1 vccd1 _05549_
+ sky130_fd_sc_hd__and3_1
X_11681_ _06128_ _06129_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__nor2_1
XANTENNA__12547__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13420_ clknet_leaf_89_clk _00376_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ datapath.PC\[15\] datapath.PC\[16\] _05489_ vssd1 vssd1 vccd1 vccd1 _05490_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_63_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10563_ keypad.alpha net1050 _05418_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__or3_1
X_13351_ clknet_4_9_0_clk _00336_ net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08045__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ _05478_ _06450_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ clknet_leaf_112_clk _00272_ net1094 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
X_10494_ net1048 _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__nor2_1
XANTENNA__07650__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12282__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ net165 net2497 net575 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12164_ _06414_ _06420_ _06419_ _06418_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07402__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ _05748_ net1295 net1288 _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_112_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ datapath.mulitply_result\[19\] datapath.multiplication_module.multiplicand_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__nor2_1
X_11046_ net1397 _05696_ mmio.WEN vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__a21o_1
XANTENNA__08363__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08115__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ net1503 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11948_ net287 net1916 net579 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XANTENNA__07469__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12457__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ _05180_ _05251_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_119_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ clknet_leaf_2_clk _00556_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13549_ clknet_leaf_79_clk _00499_ net1243 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10776__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07070_ datapath.rf.registers\[31\]\[27\] net819 net720 datapath.rf.registers\[28\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10705__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07929__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ _02892_ _02894_ _02896_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__or4_1
XANTENNA__12920__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__inv_2
X_06923_ net1001 net983 net980 _01812_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__and4_1
X_09642_ net533 net532 net405 vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__mux2_1
X_06854_ datapath.rf.registers\[2\]\[31\] net727 net723 datapath.rf.registers\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a22o_1
X_06785_ datapath.ru.latched_instruction\[31\] _01614_ _01701_ _01703_ _01711_ vssd1
+ vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a2111o_1
X_09573_ _02126_ _02128_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__nand2_2
XANTENNA__08106__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_A _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09303__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ _03120_ _01656_ _03446_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ _02723_ net516 _02789_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12367__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14077__RESET_B net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ datapath.rf.registers\[16\]\[20\] net963 net931 datapath.rf.registers\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ _03127_ _03312_ _03122_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_34_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07880__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1281_A datapath.mulitply_result\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07337_ datapath.rf.registers\[5\]\[21\] net784 net715 datapath.rf.registers\[29\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07093__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ datapath.rf.registers\[6\]\[23\] net897 net889 datapath.rf.registers\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
XANTENNA__07632__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ net391 _03817_ _03818_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__a31o_1
X_07199_ _02106_ net531 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08312__C _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout541 net544 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_8
X_09909_ _04780_ _04832_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__and3_1
Xfanout552 _06469_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_4
Xfanout563 _06466_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_8
Xfanout574 _06446_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_4
Xfanout585 _05675_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
Xfanout596 _05670_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_8
X_12920_ net1670 net217 net547 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XANTENNA__07699__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ net229 net1993 net554 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _06209_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ net239 net1934 net564 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__mux2_1
X_14521_ net1308 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
X_11733_ _01439_ _06082_ _06071_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12277__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14452_ clknet_leaf_113_clk _01339_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11664_ screen.counter.currentCt\[9\] _06116_ net667 vssd1 vssd1 vccd1 vccd1 _06118_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07871__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ clknet_leaf_89_clk _00359_ net1214 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10615_ net1564 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[27\]
+ sky130_fd_sc_hd__and2_1
X_14383_ clknet_leaf_5_clk _01270_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11595_ _05267_ _06054_ _06058_ _05763_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__o31a_1
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ clknet_leaf_92_clk _00319_ net1203 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfstp_1
XANTENNA__07084__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ keypad.apps.button\[2\] net1032 vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_114_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07623__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13265_ clknet_leaf_90_clk _00255_ net1204 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
X_10477_ _05385_ _05386_ _05387_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__or4_1
X_12216_ net249 net2324 net573 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13196_ clknet_leaf_32_clk _00188_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08222__C _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ datapath.mulitply_result\[28\] datapath.multiplication_module.multiplicand_i\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__nand2_1
X_12078_ _06347_ _06348_ _06349_ _06342_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a211o_1
X_11029_ _01441_ _05279_ _05285_ _05349_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or4_2
XANTENNA__11583__C _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06570_ net1306 net1302 mmio.key_data\[5\] vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08240_ datapath.rf.registers\[5\]\[2\] net783 net719 datapath.rf.registers\[28\]\[2\]
+ _03152_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a221o_1
XANTENNA_15 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_37 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ datapath.rf.registers\[29\]\[3\] net987 _01756_ vssd1 vssd1 vccd1 vccd1 _03098_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_133_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12915__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ datapath.rf.registers\[9\]\[26\] net779 net735 datapath.rf.registers\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07075__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08811__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07614__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ datapath.rf.registers\[30\]\[28\] net910 net886 datapath.rf.registers\[9\]\[28\]
+ _01979_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a221o_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08575__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12650__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _02881_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout479_A _06452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ net1000 net986 net981 _01801_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__and4_1
XANTENNA__10170__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ datapath.rf.registers\[20\]\[9\] net802 net746 datapath.rf.registers\[21\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a22o_1
X_09625_ _02039_ net685 _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__o211a_1
X_06837_ net996 _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout646_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09556_ _02235_ _02255_ _03497_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__o21ai_1
X_06768_ datapath.ru.latched_instruction\[17\] _01676_ _01689_ _01692_ _01694_ vssd1
+ vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ _01994_ _03361_ _03432_ _01995_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout813_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ datapath.ru.latched_instruction\[12\] net1040 net1008 _01626_ vssd1 vssd1
+ vccd1 vccd1 _01627_ sky130_fd_sc_hd__a22oi_4
X_09487_ net655 _04411_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08438_ _02105_ _02125_ _02170_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__o21a_1
XANTENNA__07853__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08369_ datapath.rf.registers\[3\]\[0\] net967 net937 datapath.rf.registers\[21\]\[0\]
+ _03295_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a221o_1
XANTENNA__12825__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _01437_ net1011 screen.counter.ct\[1\] vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a21o_1
X_11380_ screen.register.currentYbus\[9\] net130 _05875_ net159 vssd1 vssd1 vccd1
+ vccd1 _00367_ sky130_fd_sc_hd__a22o_1
XANTENNA__07605__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08604__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__C1 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ _05081_ _05237_ _05242_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__nor3_1
X_13050_ clknet_leaf_22_clk _00042_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ net373 _04317_ _05188_ net382 vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__o211ai_1
X_12001_ datapath.mulitply_result\[4\] datapath.multiplication_module.multiplicand_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08030__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ _04756_ _04785_ _04808_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__or3_1
XANTENNA__12560__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1303 net1304 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_2
Xfanout360 _03545_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_2
XANTENNA__06592__A2 _01456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout371 _03539_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_2
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_2
Xfanout393 _03519_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_2
X_13952_ clknet_leaf_48_clk _00839_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12903_ net1752 net285 net545 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
XANTENNA__11873__B1 _05234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ clknet_leaf_55_clk _00770_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ net297 net1633 net553 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12765_ net630 _05666_ _06443_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__or3_4
XANTENNA__08097__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14504_ clknet_leaf_12_clk _01391_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11716_ _06068_ _06150_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__nor2_1
XANTENNA__07844__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12696_ net2139 net172 net434 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ clknet_leaf_103_clk _01322_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10466__D _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11647_ net2603 _06104_ net666 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12735__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11928__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07057__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput35 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_96_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14366_ clknet_leaf_51_clk _01253_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11578_ _06036_ _06042_ _06031_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13317_ clknet_leaf_112_clk _00307_ net1098 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10600__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold808 datapath.rf.registers\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ keypad.apps.button\[1\] net1032 vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__and2_1
Xhold819 datapath.rf.registers\[24\]\[18\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
X_14297_ clknet_leaf_47_clk _01184_ net1197 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13248_ clknet_leaf_76_clk _00238_ net1248 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ clknet_leaf_55_clk _00171_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07740_ datapath.rf.registers\[6\]\[12\] net813 net755 datapath.rf.registers\[24\]\[12\]
+ _02666_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ datapath.rf.registers\[7\]\[14\] net956 net920 datapath.rf.registers\[2\]\[14\]
+ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08190__D1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09410_ _04310_ _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06622_ datapath.ru.latched_instruction\[20\] datapath.ru.latched_instruction\[21\]
+ datapath.ru.latched_instruction\[22\] datapath.ru.latched_instruction\[23\] vssd1
+ vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_140_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06553_ mmio.memload_or_instruction\[25\] net1063 vssd1 vssd1 vccd1 vccd1 _01483_
+ sky130_fd_sc_hd__and2_1
X_09341_ net640 _04267_ net612 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08088__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09285__A1 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07296__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06484_ datapath.ru.latched_instruction\[17\] vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
X_09272_ net498 net495 net512 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08223_ datapath.rf.registers\[14\]\[2\] net994 _01752_ vssd1 vssd1 vccd1 vccd1 _03150_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12645__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_A _05502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__B1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ datapath.rf.registers\[3\]\[3\] net964 net929 datapath.rf.registers\[4\]\[3\]
+ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10052__C1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ datapath.rf.registers\[2\]\[27\] net922 net894 datapath.rf.registers\[14\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
X_08085_ datapath.rf.registers\[25\]\[5\] net796 net740 datapath.rf.registers\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a22o_1
XANTENNA__08260__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07036_ datapath.rf.registers\[1\]\[28\] net741 net715 datapath.rf.registers\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout596_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10679__A1_N _01473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _02568_ _03328_ _02526_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout763_A _01767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07938_ datapath.rf.registers\[26\]\[8\] net820 _02863_ _02864_ net831 vssd1 vssd1
+ vccd1 vccd1 _02865_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__09512__A2 _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__B1 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ datapath.rf.registers\[31\]\[9\] net949 net889 datapath.rf.registers\[12\]\[9\]
+ _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout930_A _01820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ net625 _04520_ _04522_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a31o_1
X_10880_ net215 net2191 net600 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ net707 _04450_ net623 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08079__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08318__B _03210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ net246 net2359 net449 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__mux2_1
XANTENNA__07826__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _05930_ _05960_ _05961_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__or4b_1
XFILLER_0_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12481_ net257 net2323 net456 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__mux2_1
XANTENNA__12555__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07039__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ clknet_leaf_31_clk _01107_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11432_ screen.register.currentXbus\[0\] _05720_ net1013 screen.register.currentXbus\[24\]
+ _05724_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11386__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ clknet_leaf_19_clk _01038_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11363_ _03244_ net668 vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08251__A2 _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ clknet_leaf_1_clk _00094_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10314_ net844 _04661_ _05240_ net1245 vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_60_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14082_ clknet_leaf_43_clk _00969_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294_ net15 net1046 net1035 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1
+ vccd1 _00308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ clknet_leaf_3_clk _00025_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12290__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net536 _05171_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__nand2_1
Xfanout1100 net1102 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
Xfanout1111 net1125 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07211__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1122 net1124 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_4
X_10176_ datapath.PC\[13\] net1310 _05101_ _05102_ vssd1 vssd1 vccd1 vccd1 _05103_
+ sky130_fd_sc_hd__a22o_1
Xfanout1133 net1135 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
Xfanout1144 net1200 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_2
Xfanout1155 net1163 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_2
Xfanout1166 net1171 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1177 net1180 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
Xfanout1188 net1189 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_4
Xfanout1199 net1200 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_2
XANTENNA__08306__A3 _01776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13935_ clknet_leaf_3_clk _00822_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13866_ clknet_leaf_11_clk _00753_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10758__B _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12817_ _05496_ net2004 net558 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13797_ clknet_leaf_108_clk _00684_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07278__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ net247 net1700 net567 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13744__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12465__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ net2340 net258 net431 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14418_ clknet_leaf_35_clk _01305_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14349_ clknet_leaf_1_clk _01236_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold605 datapath.rf.registers\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 datapath.rf.registers\[31\]\[18\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 datapath.rf.registers\[20\]\[19\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 datapath.rf.registers\[19\]\[18\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold649 datapath.rf.registers\[8\]\[20\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ net415 _03836_ _03835_ net318 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__o211a_1
X_09890_ _04814_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09075__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07202__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08841_ net527 net359 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__or2_1
XANTENNA__06849__D net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ net611 _03694_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a21o_1
XANTENNA__06961__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ datapath.rf.registers\[22\]\[13\] net952 net920 datapath.rf.registers\[2\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_108_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ datapath.rf.registers\[4\]\[14\] net809 net740 datapath.rf.registers\[1\]\[14\]
+ _02580_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06605_ _01491_ _01498_ _01527_ _01534_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__or4_1
X_07585_ datapath.rf.registers\[4\]\[16\] net931 net863 datapath.rf.registers\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a22o_1
XANTENNA__08138__B _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07269__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ net383 _04249_ _04250_ _04248_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__a31o_1
X_06536_ net1307 net1304 mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ _01466_ sky130_fd_sc_hd__or3b_2
XANTENNA__07808__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09255_ _02978_ _03316_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__xor2_1
XANTENNA__12375__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_A _02951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1253_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ datapath.rf.registers\[11\]\[2\] net969 _03128_ _03130_ _03132_ vssd1 vssd1
+ vccd1 vccd1 _03133_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_117_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09186_ net636 _04096_ _04111_ net611 vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08137_ net507 _03062_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__and2_1
XANTENNA__08233__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09430__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ datapath.rf.registers\[25\]\[5\] net872 net864 datapath.rf.registers\[13\]\[5\]
+ _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout880_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ datapath.rf.registers\[10\]\[29\] net918 net866 datapath.rf.registers\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ datapath.PC\[20\] _03582_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_126_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11981_ _06267_ _06268_ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__nor2_1
X_13720_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[5\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[5\] sky130_fd_sc_hd__dfrtp_1
X_10932_ net281 net2126 net590 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13651_ clknet_leaf_68_clk _00589_ net1225 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10863_ _05607_ net2216 net598 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08048__B _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12602_ net2330 net289 net443 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
X_13582_ clknet_leaf_80_clk _00532_ net1234 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10794_ _01481_ net659 _05626_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_155_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ net2145 net164 net454 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__mux2_1
XANTENNA__12285__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12464_ net184 net2164 net461 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14203_ clknet_leaf_52_clk _01090_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11415_ net343 net714 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12395_ net196 net1871 net470 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ clknet_leaf_26_clk _01021_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07432__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _01483_ net1030 net310 net314 net2646 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14065_ clknet_leaf_7_clk _00952_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06634__A_N mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ net28 net1044 net1033 net2582 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__o22a_1
X_13016_ clknet_leaf_34_clk _00008_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10228_ _04812_ _04813_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08230__C _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2 keypad.debounce.debounce\[5\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ datapath.PC\[11\] _04081_ net536 vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07499__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11295__B2 mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ clknet_leaf_49_clk _00805_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10488__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13849_ clknet_leaf_61_clk _00736_ net1265 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07370_ datapath.rf.registers\[10\]\[21\] net917 net849 datapath.rf.registers\[1\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10708__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ net329 _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__nand2_1
XANTENNA__07671__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08215__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold402 datapath.rf.registers\[19\]\[19\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold413 datapath.rf.registers\[25\]\[21\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 datapath.rf.registers\[10\]\[26\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 datapath.rf.registers\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 datapath.rf.registers\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 datapath.rf.registers\[20\]\[3\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 datapath.rf.registers\[5\]\[11\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _03637_ _04585_ _04608_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a21oi_1
Xhold479 datapath.rf.registers\[31\]\[19\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout904 net907 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_55_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout915 _01830_ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
Xfanout926 net927 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 _01817_ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_2
X_09873_ _04748_ _04750_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__xnor2_1
Xfanout948 net951 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout294_A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 _01809_ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ _03499_ _03748_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__nand2_1
Xhold1102 datapath.rf.registers\[20\]\[23\] vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 datapath.rf.registers\[18\]\[23\] vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 datapath.rf.registers\[9\]\[3\] vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 datapath.rf.registers\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 datapath.rf.registers\[21\]\[13\] vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11782__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1157 datapath.rf.registers\[16\]\[3\] vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net362 _03677_ _03678_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a31o_1
Xhold1168 datapath.rf.registers\[16\]\[12\] vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1179 datapath.rf.registers\[8\]\[7\] vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ datapath.rf.registers\[0\]\[13\] _02632_ net830 vssd1 vssd1 vccd1 vccd1 _02633_
+ sky130_fd_sc_hd__mux2_4
XANTENNA__11286__B2 mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ net414 _03611_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__or2_1
X_07637_ _02557_ _02559_ _02561_ _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout726_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ datapath.rf.registers\[3\]\[16\] net768 net750 datapath.rf.registers\[10\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ net505 net504 net684 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__o21ai_1
X_06519_ keypad.decode.push net1448 net1032 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky_n\[4\]
+ sky130_fd_sc_hd__mux2_1
X_07499_ datapath.rf.registers\[8\]\[18\] net926 net858 datapath.rf.registers\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07662__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ net500 net621 net489 net511 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08206__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12833__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ net329 _04093_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o21a_1
X_11200_ _05181_ _05211_ net137 net144 net1524 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__a32o_1
X_12180_ columns.count\[4\] _01447_ _05849_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__nand3_1
XANTENNA__06768__A2 _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _05715_ net1020 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08331__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold980 datapath.rf.registers\[2\]\[24\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold991 datapath.rf.registers\[23\]\[31\] vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net1022 _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__or2_2
X_10013_ net705 _04518_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__and2_1
XANTENNA__07193__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06940__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ net236 net1863 net578 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13703_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[20\]
+ net1262 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ net211 net2053 net597 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__mux2_1
X_11895_ _05880_ _06263_ net149 net1434 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13634_ clknet_leaf_45_clk _00572_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10846_ net1609 net211 net604 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13565_ clknet_leaf_80_clk _00515_ net1234 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ net1639 _05613_ net602 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09642__A1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ net1706 net249 net452 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__mux2_1
XANTENNA__10252__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07653__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13496_ clknet_leaf_73_clk _00446_ net1245 vssd1 vssd1 vccd1 vccd1 datapath.PC\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08225__C _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12447_ net262 net1953 net460 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12743__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10004__A2 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12378_ net275 net2413 net470 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__mux2_1
XANTENNA__10771__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ clknet_leaf_93_clk _01004_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11329_ mmio.memload_or_instruction\[8\] net1062 net307 net311 datapath.ru.latched_instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10490__C net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09158__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14048_ clknet_leaf_48_clk _00935_ net1195 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_06870_ _01785_ _01786_ _01792_ _01794_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__or4_1
XANTENNA__07184__A2 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07572__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ net512 net510 net407 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08471_ _02977_ _03395_ _03396_ _02976_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__o31a_1
XANTENNA__12918__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07422_ _02346_ _02347_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__nor2_2
XANTENNA__07892__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06543__C_N mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07353_ net832 _02279_ _02261_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11123__A _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07644__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07284_ datapath.rf.registers\[7\]\[23\] net958 _02206_ _02207_ _02210_ vssd1 vssd1
+ vccd1 vccd1 _02211_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06998__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09023_ net499 net620 net488 net520 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12653__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_A _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 datapath.rf.registers\[22\]\[17\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 datapath.multiplication_module.multiplicand_i\[10\] vssd1 vssd1 vccd1 vccd1
+ net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 datapath.rf.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 datapath.rf.registers\[25\]\[24\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 datapath.rf.registers\[16\]\[7\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 datapath.rf.registers\[16\]\[1\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold276 datapath.rf.registers\[17\]\[4\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 datapath.rf.registers\[31\]\[25\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 net703 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout712 _06097_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_2
Xhold298 datapath.rf.registers\[10\]\[25\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ datapath.PC\[29\] net628 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nand2_1
Xfanout723 net725 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
Xfanout734 _01777_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
Xfanout745 _01773_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net758 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
XANTENNA__10901__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ _04676_ _04767_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__xor2_2
Xfanout767 net769 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_8
Xfanout778 net781 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
Xfanout789 net792 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_4
XANTENNA__07175__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ net417 _03466_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_29_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ datapath.PC\[10\] _02784_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout843_A _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ datapath.rf.registers\[20\]\[29\] net803 net724 datapath.rf.registers\[27\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XANTENNA__06922__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ net527 net526 net405 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12828__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ net189 net2303 net608 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__mux2_1
XANTENNA__06686__A1 _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ screen.counter.currentCt\[14\] _06126_ net667 vssd1 vssd1 vccd1 vccd1 _06129_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10631_ datapath.PC\[14\] _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_81_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08326__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13350_ clknet_leaf_69_clk _00335_ net1224 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07635__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10562_ _05410_ _05413_ _05469_ _05468_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a31oi_1
Xmax_cap1018 _01530_ vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_1
X_12301_ _01643_ _01667_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__or2_2
XANTENNA__06989__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ clknet_leaf_112_clk _00271_ net1096 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10493_ net1050 _05399_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12232_ net168 net2422 net575 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__mux2_1
XANTENNA__08060__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _06418_ _06419_ _06420_ _06414_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a211o_1
XANTENNA__10942__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11114_ net1296 net1292 screen.counter.ct\[8\] net1287 vssd1 vssd1 vccd1 vccd1 _05764_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_112_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ datapath.mulitply_result\[19\] datapath.multiplication_module.multiplicand_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__and2_1
X_11045_ _01435_ screen.register.xFill3 _01436_ screen.register.cFill3 _05695_ vssd1
+ vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__o221a_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07166__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06913__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ net2320 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09312__A0 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06566__C_N mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11947_ net182 net1561 net579 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__mux2_1
XANTENNA__12738__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ net1383 _01443_ _06262_ net1499 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a22o_1
XANTENNA__08517__A _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13617_ clknet_leaf_3_clk _00555_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ _05490_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13548_ clknet_leaf_88_clk _00498_ net1211 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11422__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08823__C1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13479_ clknet_leaf_83_clk _00432_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12473__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08252__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ datapath.rf.registers\[25\]\[7\] net872 net868 datapath.rf.registers\[27\]\[7\]
+ _02897_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a221o_1
X_09710_ _02435_ _02436_ _03832_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__or3_1
X_06922_ datapath.rf.registers\[25\]\[31\] net873 net870 datapath.rf.registers\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a22o_1
XANTENNA__10721__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09641_ _01996_ net678 _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__o21ai_1
X_06853_ net988 _01763_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__and2_1
XANTENNA__10161__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09572_ _03703_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__nand2_1
X_06784_ _01658_ _01660_ _01670_ _01710_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__or4_1
X_08523_ _03121_ _01657_ _03446_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12648__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _02723_ net516 vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07405_ datapath.rf.registers\[22\]\[20\] net954 net874 datapath.rf.registers\[25\]\[20\]
+ _02331_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ _03182_ _03311_ _03179_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_63_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1166_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ datapath.rf.registers\[11\]\[21\] net775 net746 datapath.rf.registers\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12383__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ datapath.rf.registers\[4\]\[23\] net930 net910 datapath.rf.registers\[30\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09006_ net396 _03931_ _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__and3_1
XANTENNA__09258__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07198_ datapath.rf.registers\[0\]\[25\] net693 _02111_ _02124_ vssd1 vssd1 vccd1
+ vccd1 _02125_ sky130_fd_sc_hd__o22a_2
XANTENNA_fanout793_A _01757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08253__A_N net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout960_A _01806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _02566_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_4
Xfanout531 _02125_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_8
X_09908_ _04774_ _04834_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__xnor2_2
Xfanout553 net556 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_6
Xfanout564 _06466_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_4
Xfanout575 _06446_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07148__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 net589 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_6
XANTENNA__06589__C_N mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _04685_ _04687_ _04764_ _04683_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a31o_1
Xfanout597 _05670_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_4
X_12850_ net242 net2496 net554 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11801_ datapath.PC\[11\] net302 _06206_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_83_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12558__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12781_ net245 net2430 net563 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__mux2_1
X_14520_ net1308 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
X_11732_ net2644 net663 _06160_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07856__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07320__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14451_ clknet_leaf_59_clk _01338_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11663_ _06116_ _06117_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13402_ clknet_leaf_86_clk _00358_ net1231 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10614_ net2624 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[26\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07608__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ clknet_leaf_116_clk _01269_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ _05705_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ clknet_leaf_78_clk mmio.ack_center.key_en net1243 vssd1 vssd1 vccd1 vccd1
+ mmio.key_en1 sky130_fd_sc_hd__dfrtp_1
X_10545_ keypad.alpha _05453_ _05454_ _05448_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[1\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08281__B1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12293__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13264_ clknet_leaf_109_clk _00254_ net1107 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10476_ screen.register.currentYbus\[13\] screen.register.currentYbus\[12\] screen.register.currentYbus\[15\]
+ screen.register.currentYbus\[14\] vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__or4_1
XANTENNA__12904__A1 _05607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net254 net2218 net573 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__mux2_1
XANTENNA__08033__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ clknet_leaf_68_clk _00187_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07387__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net323 _06405_ _06406_ net327 net2146 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a32o_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07792__C1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _06335_ _06340_ _06343_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07139__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ _05265_ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13351__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09631__A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12979_ net241 net2045 net608 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07847__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07151__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07311__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09049__C1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_27 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__A2 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08170_ datapath.rf.registers\[1\]\[3\] net740 net719 datapath.rf.registers\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a22o_1
XANTENNA_38 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07121_ datapath.rf.registers\[20\]\[26\] net802 net787 datapath.rf.registers\[23\]\[26\]
+ _02047_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a221o_1
XANTENNA__08272__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11401__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07052_ datapath.rf.registers\[11\]\[28\] net970 net870 datapath.rf.registers\[27\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__10707__A2_N _05553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__12931__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07954_ net513 _02879_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_145_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06905_ datapath.rf.registers\[18\]\[31\] net914 net910 datapath.rf.registers\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a22o_1
X_07885_ datapath.rf.registers\[0\]\[9\] net692 _02799_ _02811_ vssd1 vssd1 vccd1
+ vccd1 _02812_ sky130_fd_sc_hd__o22a_4
XANTENNA__07535__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _02040_ net681 net678 _04542_ _04547_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__o221a_1
X_06836_ _01638_ _01646_ net982 _01682_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__and4_2
XANTENNA__10685__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13021__RESET_B net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09555_ net416 _04431_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__o21ai_1
X_06767_ datapath.ru.latched_instruction\[6\] _01583_ net997 datapath.ru.latched_instruction\[24\]
+ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12378__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09288__C1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ _03361_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__nor2_1
XANTENNA__07838__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ net613 _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06698_ datapath.ru.latched_instruction\[12\] _01509_ net1029 vssd1 vssd1 vccd1 vccd1
+ _01626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07302__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08437_ _03363_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout806_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ datapath.rf.registers\[22\]\[0\] net952 net935 datapath.rf.registers\[23\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07319_ datapath.rf.registers\[24\]\[22\] net906 net898 datapath.rf.registers\[6\]\[22\]
+ _02245_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a221o_1
XANTENNA__08263__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08299_ datapath.rf.registers\[31\]\[1\] net991 _01746_ vssd1 vssd1 vccd1 vccd1 _03226_
+ sky130_fd_sc_hd__and3_1
X_10330_ mmio.wishbone.curr_state\[0\] _05248_ _05251_ _05254_ vssd1 vssd1 vccd1 vccd1
+ _05256_ sky130_fd_sc_hd__and4_4
XANTENNA__08015__B1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ net365 _05187_ _05186_ net369 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a211o_1
XANTENNA__12841__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07369__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ datapath.mulitply_result\[3\] net326 net322 _06284_ vssd1 vssd1 vccd1 vccd1
+ _00578_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10192_ net701 _05118_ _05115_ net200 vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1304 mmio.key_en2 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__clkbuf_2
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xfanout361 net364 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_2
Xfanout372 _03539_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_1
XANTENNA__10125__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout383 _03535_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_1
X_13951_ clknet_leaf_36_clk _00838_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout394 net397 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_2
X_12902_ net1744 net295 net546 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
XANTENNA__11873__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13882_ clknet_leaf_22_clk _00769_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07541__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ net288 net1674 net553 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12288__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ net166 net2591 net568 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11715_ net1296 _05714_ net1295 vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__a21oi_1
X_14503_ clknet_leaf_25_clk _01390_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12695_ net2071 net186 net433 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11646_ screen.counter.currentCt\[3\] _06104_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__and2_1
X_14434_ clknet_leaf_43_clk _01321_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ clknet_leaf_32_clk _01252_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput36 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_11577_ _05721_ _05806_ _05810_ _05711_ _05323_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_103_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_96_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13316_ clknet_leaf_110_clk _00306_ net1106 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_10528_ _05430_ _05438_ _05428_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[0\]
+ sky130_fd_sc_hd__a21oi_1
X_14296_ clknet_leaf_40_clk _01183_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold809 datapath.rf.registers\[18\]\[26\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08006__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13247_ clknet_leaf_75_clk _00237_ net1251 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12751__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ net519 _02654_ _02698_ _02742_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13178_ clknet_leaf_22_clk _00170_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08530__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _06387_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__nand2_1
XANTENNA_wire342_A _02280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07780__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11313__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ datapath.rf.registers\[14\]\[14\] net892 net872 datapath.rf.registers\[25\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
XANTENNA__07532__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ _01532_ _01535_ _01543_ _01550_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__nor4_1
XFILLER_0_149_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ net339 _04256_ _04257_ _04265_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a32o_1
X_06552_ datapath.ru.latched_instruction\[10\] _01481_ _01416_ _01479_ vssd1 vssd1
+ vccd1 vccd1 _01482_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ net502 net617 net496 net513 vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__a211o_1
XANTENNA__12926__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06483_ datapath.ru.latched_instruction\[16\] vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
X_08222_ datapath.rf.registers\[20\]\[2\] net989 _01734_ vssd1 vssd1 vccd1 vccd1 _03149_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08153_ datapath.rf.registers\[21\]\[3\] net937 net867 datapath.rf.registers\[13\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07104_ datapath.rf.registers\[10\]\[27\] net918 net906 datapath.rf.registers\[24\]\[27\]
+ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a221o_1
XANTENNA__08796__A1 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ datapath.rf.registers\[26\]\[5\] net820 net782 datapath.rf.registers\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__a22o_1
X_07035_ datapath.rf.registers\[14\]\[28\] net800 net797 datapath.rf.registers\[25\]\[28\]
+ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a221o_1
XANTENNA__12661__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout491_A _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__inv_2
XANTENNA__07771__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ datapath.rf.registers\[4\]\[8\] net809 net781 datapath.rf.registers\[9\]\[8\]
+ _02857_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__a221o_1
XANTENNA__11304__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ datapath.rf.registers\[19\]\[9\] net945 net858 datapath.rf.registers\[15\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__a22o_1
XANTENNA__07523__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06819_ _01639_ _01646_ net982 _01682_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__and4_2
X_09607_ net654 _04533_ _04530_ _04532_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__or4b_1
X_07799_ datapath.rf.registers\[13\]\[11\] net864 net852 datapath.rf.registers\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a22o_1
X_09538_ net707 _04464_ _03556_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__o21a_1
XANTENNA__07503__B net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _02787_ net687 _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12836__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ net975 _05917_ _05967_ _05969_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and4_1
X_12480_ net261 net2499 net456 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ net975 _05816_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150_ clknet_leaf_114_clk _01037_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09984__B1 _03567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ net2613 net130 _05866_ net159 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__a22o_1
XANTENNA__08251__A3 _03175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10594__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ clknet_leaf_119_clk _00093_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ _01423_ _05239_ net1051 vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__mux2_1
XANTENNA__12571__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ clknet_leaf_43_clk _00968_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11293_ net14 net1045 net1034 net2555 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__o22a_1
X_13032_ clknet_leaf_13_clk _00024_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10244_ net1055 _05170_ net699 vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_91_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09200__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1102 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10091__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ net200 _04812_ _05093_ net1250 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__o31a_1
Xfanout1123 net1124 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_2
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07762__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1145 net1146 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_4
Xfanout1156 net1158 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_4
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout180 net183 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06970__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1180 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_4
Xfanout191 _05548_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1189 net1199 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13934_ clknet_leaf_116_clk _00821_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07514__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ clknet_leaf_3_clk _00752_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12816_ net236 net2101 net557 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__mux2_1
X_13796_ clknet_leaf_14_clk _00683_ net1115 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__C _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12746__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12747_ net249 net1928 net565 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12678_ net2140 net261 net431 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
XANTENNA__08525__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11629_ screen.counter.currentCt\[9\] screen.counter.currentCt\[8\] screen.counter.currentCt\[11\]
+ screen.counter.currentCt\[10\] vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__or4_1
X_14417_ clknet_leaf_27_clk _01304_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ clknet_leaf_31_clk _01235_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10585__A1 _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold606 datapath.rf.registers\[30\]\[25\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 datapath.rf.registers\[20\]\[15\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 datapath.rf.registers\[17\]\[11\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12481__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold639 datapath.rf.registers\[22\]\[8\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ clknet_leaf_21_clk _01166_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08840_ net364 _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__and3_1
XANTENNA__07753__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08771_ net334 _03684_ net635 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__o21a_1
X_07722_ datapath.rf.registers\[10\]\[13\] net916 net868 datapath.rf.registers\[27\]\[13\]
+ _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ datapath.rf.registers\[13\]\[14\] net795 net766 datapath.rf.registers\[3\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06604_ datapath.ru.latched_instruction\[8\] _01472_ _01511_ _01415_ _01533_ vssd1
+ vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a221o_1
X_07584_ datapath.rf.registers\[24\]\[16\] net906 net887 datapath.rf.registers\[9\]\[16\]
+ _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09323_ _04151_ _04152_ net374 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__a21o_1
X_06535_ _01407_ _01464_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__and2_1
XANTENNA__12656__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ net335 _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__nor2_1
XANTENNA__10812__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08205_ datapath.rf.registers\[3\]\[2\] net964 net960 datapath.rf.registers\[16\]\[2\]
+ _03131_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a221o_1
X_09185_ net638 _04096_ _04110_ _04111_ net655 vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09415__C1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_A _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__C1 _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ net507 _03061_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__A1 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12391__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ datapath.rf.registers\[26\]\[5\] net940 net932 datapath.rf.registers\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__a22o_1
XANTENNA__10904__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ datapath.rf.registers\[23\]\[29\] net934 net859 datapath.rf.registers\[15\]\[29\]
+ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_73_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout873_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07744__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__inv_2
XANTENNA__06952__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ datapath.multiplication_module.multiplier_i\[0\] datapath.mulitply_result\[0\]
+ datapath.multiplication_module.multiplicand_i\[0\] net350 vssd1 vssd1 vccd1 vccd1
+ _06268_ sky130_fd_sc_hd__a31o_1
X_10931_ net283 net2131 net590 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10862_ net283 net2361 net598 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__mux2_1
X_13650_ clknet_leaf_101_clk _00588_ net1223 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12601_ net1505 net182 net440 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13581_ clknet_leaf_79_clk _00531_ net1233 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10793_ datapath.mulitply_result\[10\] net426 net658 vssd1 vssd1 vccd1 vccd1 _05627_
+ sky130_fd_sc_hd__a21oi_2
XANTENNA__12566__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ net2473 net170 net454 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ net188 net2200 net462 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11414_ screen.register.currentYbus\[26\] net130 _05892_ net159 vssd1 vssd1 vccd1
+ vccd1 _00384_ sky130_fd_sc_hd__a22o_1
X_14202_ clknet_leaf_23_clk _01089_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12394_ net209 net1942 net470 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ clknet_leaf_28_clk _01020_ net1130 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11345_ mmio.memload_or_instruction\[24\] net1058 net307 net311 datapath.ru.latched_instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__a32o_1
XANTENNA__10814__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07983__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ clknet_leaf_0_clk _00951_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11276_ net27 net1047 net1036 net1531 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__a22o_1
XANTENNA__11516__B1 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ clknet_leaf_44_clk _00007_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10227_ net1277 net1310 _05151_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10158_ net833 _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nor2_1
Xhold3 keypad.debounce.debounce\[9\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06943__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ _04817_ _04819_ _04821_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13917_ clknet_leaf_33_clk _00804_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11295__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__C net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13848_ clknet_leaf_40_clk _00735_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12476__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13779_ clknet_leaf_49_clk _00666_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08255__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07120__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold403 datapath.rf.registers\[4\]\[27\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold414 datapath.rf.registers\[18\]\[8\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 datapath.rf.registers\[23\]\[3\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10724__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold436 datapath.rf.registers\[8\]\[16\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 datapath.rf.registers\[15\]\[26\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 datapath.rf.registers\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold469 datapath.rf.registers\[5\]\[13\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ datapath.PC\[31\] net1312 _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__buf_4
Xfanout916 net919 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_4
Xfanout927 _01825_ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_4
X_09872_ _04797_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_5_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07187__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout938 _01817_ vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_4
XFILLER_0_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout949 net951 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__buf_4
Xhold1103 datapath.mulitply_result\[28\] vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ net417 _03614_ _03749_ net317 vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__a211o_1
Xhold1114 datapath.rf.registers\[6\]\[23\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1125 datapath.rf.registers\[30\]\[21\] vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1136 datapath.rf.registers\[29\]\[17\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 datapath.rf.registers\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net368 _03679_ _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__and3_1
Xhold1158 datapath.rf.registers\[12\]\[23\] vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 datapath.rf.registers\[28\]\[10\] vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ datapath.rf.registers\[8\]\[13\] net737 _02628_ _02630_ _02631_ vssd1 vssd1
+ vccd1 vccd1 _02632_ sky130_fd_sc_hd__a2111o_2
X_08685_ _03460_ _03480_ net341 vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_92_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08151__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ datapath.rf.registers\[24\]\[15\] net905 net886 datapath.rf.registers\[9\]\[15\]
+ _02562_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07567_ datapath.rf.registers\[20\]\[16\] net803 net753 datapath.rf.registers\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a22o_1
XANTENNA__12386__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout719_A _01782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10246__B1 _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09306_ net419 net414 net317 _04121_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__or4_1
X_06518_ columns.count\[0\] _01447_ _01448_ _01449_ vssd1 vssd1 vccd1 vccd1 _01450_
+ sky130_fd_sc_hd__or4_2
XFILLER_0_118_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07498_ datapath.rf.registers\[11\]\[18\] net970 net933 datapath.rf.registers\[23\]\[18\]
+ _02416_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ net513 _02812_ net356 vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09939__B1 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ net383 _04092_ _04094_ net332 vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__a211o_1
X_08119_ datapath.rf.registers\[18\]\[4\] net792 net778 datapath.rf.registers\[9\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a22o_1
X_09099_ net498 net495 net517 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a21o_1
X_11130_ _05717_ net1020 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__nor2_1
XANTENNA__07965__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold970 datapath.rf.registers\[18\]\[30\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 datapath.rf.registers\[26\]\[26\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08331__C _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold992 datapath.rf.registers\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ net1300 net1301 _05698_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or3_2
XANTENNA__07178__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07717__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ net1057 _04938_ _04937_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06925__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ net239 net2032 net581 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__mux2_1
XANTENNA__08142__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_83_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[19\]
+ net1258 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ net214 net2318 net596 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__mux2_1
X_11894_ _05879_ _06263_ net149 net1423 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__a22o_1
XANTENNA__07350__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10845_ net1698 net214 net603 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__mux2_1
X_13633_ clknet_leaf_39_clk _00571_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12296__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ clknet_leaf_89_clk _00514_ net1216 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10776_ _01470_ net709 _05612_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__o21a_2
XFILLER_0_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07102__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12515_ net2137 net253 net452 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__mux2_1
X_13495_ clknet_leaf_80_clk net1383 net1239 vssd1 vssd1 vccd1 vccd1 screen.screenEdge.enable3
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08850__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ net267 net2152 net460 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12377_ net279 net1761 net468 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__mux2_1
XANTENNA__11201__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11328_ _01470_ net1028 net307 net311 datapath.ru.latched_instruction\[7\] vssd1
+ vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__a32o_1
X_14116_ clknet_leaf_17_clk _01003_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11259_ net530 _05844_ net140 net1463 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14047_ clknet_leaf_38_clk _00934_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07169__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07708__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08470_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07341__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07352_ datapath.rf.registers\[31\]\[21\] net818 _02262_ _02270_ _02278_ vssd1 vssd1
+ vccd1 vccd1 _02279_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07283_ net694 _02196_ _02197_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__or4_1
XANTENNA__12934__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ net392 _03856_ _03857_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold200 keypad.apps.button\[3\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 datapath.rf.registers\[10\]\[3\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold222 datapath.rf.registers\[7\]\[14\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold233 net44 vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 net73 vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 datapath.rf.registers\[6\]\[4\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 datapath.rf.registers\[3\]\[7\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 datapath.rf.registers\[4\]\[8\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 datapath.rf.registers\[22\]\[18\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 datapath.rf.registers\[31\]\[7\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlymetal6s2s_1
X_09924_ datapath.PC\[29\] net628 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nor2_1
Xfanout713 _06097_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1111_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_4
Xfanout735 _01777_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
Xfanout746 _01773_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_4
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 net758 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
X_09855_ _04770_ _04781_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout571_A _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_4
Xfanout779 net781 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_4
XANTENNA_fanout669_A _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08806_ net422 _03482_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__or2_1
X_09786_ datapath.PC\[10\] _02784_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__and2_1
X_06998_ datapath.rf.registers\[14\]\[29\] net801 net757 datapath.rf.registers\[24\]\[29\]
+ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_29_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ net529 net528 net405 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_65_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout836_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08124__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _03359_ _03360_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_101_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ net647 net423 net626 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08599_ net384 _03525_ _03524_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10630_ net1276 datapath.PC\[13\] _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_81_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09624__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08326__C _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10561_ keypad.apps.button\[3\] net1032 vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12844__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap1019 _06096_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_1
X_12300_ net1935 net165 net482 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__mux2_1
X_13280_ clknet_leaf_92_clk _00270_ net1202 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
X_10492_ net1050 _05399_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ net172 net2584 net576 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__mux2_1
XANTENNA__09388__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07399__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08342__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _06407_ _06411_ _06415_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a21oi_1
X_11113_ net1023 _05731_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_112_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12093_ _06357_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ net1024 _05691_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08899__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output121_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12995_ net1538 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_56_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08115__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09312__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11946_ net631 _05669_ _05671_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__or3_4
XFILLER_0_143_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07323__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ screen.counter.ack3 screen.counter.ack2 vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13616_ clknet_leaf_1_clk _00554_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ datapath.PC\[15\] _05489_ datapath.PC\[16\] vssd1 vssd1 vccd1 vccd1 _05656_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_119_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12754__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11422__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ clknet_leaf_90_clk _00497_ net1209 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10759_ datapath.PC\[5\] _05482_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_99_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13478_ clknet_leaf_84_clk _00431_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09379__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12429_ net1846 net195 net465 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08252__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06601__A2 _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ datapath.rf.registers\[26\]\[7\] net940 net864 datapath.rf.registers\[13\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a22o_1
X_06921_ net1000 net983 net979 _01801_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_147_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08354__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06852_ net973 _01741_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__and2_1
X_09640_ _01992_ net685 net682 _01993_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__o22a_1
XANTENNA__10303__A _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ _03747_ _03785_ _04474_ _04496_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__and4b_1
X_06783_ _01590_ _01659_ net977 datapath.ru.latched_instruction\[20\] _01709_ vssd1
+ vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a221o_1
XANTENNA__10022__B _03785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08106__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09303__A1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ _03444_ _03447_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__nand2_4
XANTENNA__07314__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08453_ _02634_ _02655_ _02700_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07404_ datapath.rf.registers\[12\]\[20\] net890 net850 datapath.rf.registers\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a22o_1
X_08384_ _03249_ _03288_ _03307_ _03248_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07335_ datapath.rf.registers\[20\]\[21\] net802 net752 datapath.rf.registers\[22\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a22o_1
XANTENNA__12664__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1159_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07266_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__inv_2
XANTENNA__07093__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09005_ net523 net356 _03929_ net389 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07197_ _02119_ _02121_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__or3_1
XANTENNA__08162__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A1 screen.screenLogic.currentWrx vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_A _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10912__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 _02951_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
Xfanout521 _02520_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_4
X_09907_ _04669_ _04773_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__or2_1
Xfanout532 _02038_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_4
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_8
Xfanout565 _06465_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_8
Xfanout576 _06446_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_4
X_09838_ _04687_ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__nand2_1
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07506__B _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout598 _05668_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_4
XANTENNA__10213__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ datapath.PC\[15\] net632 _04694_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__or3_1
XANTENNA__12839__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
X_11800_ _04663_ _05630_ net302 _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_83_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ net251 net1864 net561 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11731_ screen.counter.ct\[11\] _06077_ _06082_ _06098_ vssd1 vssd1 vccd1 vccd1 _06160_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10860__A0 _05590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14450_ clknet_leaf_34_clk _01337_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11662_ screen.counter.currentCt\[8\] _06114_ net667 vssd1 vssd1 vccd1 vccd1 _06117_
+ sky130_fd_sc_hd__o21ai_1
X_13401_ clknet_leaf_77_clk _00002_ net1246 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10613_ net1521 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[25\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12574__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14381_ clknet_leaf_0_clk _01268_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11593_ _01437_ net1294 net1284 net1282 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_12_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10544_ net1050 net1026 net1025 _05441_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__or4_1
X_13332_ clknet_leaf_97_clk net1375 net1230 vssd1 vssd1 vccd1 vccd1 mmio.key_en2 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09449__A _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07084__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10475_ screen.register.currentYbus\[9\] screen.register.currentYbus\[8\] screen.register.currentYbus\[11\]
+ screen.register.currentYbus\[10\] vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__or4_1
X_13263_ clknet_leaf_110_clk _00253_ net1104 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08569__C1 _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ net259 net2374 net573 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13194_ clknet_leaf_12_clk _00186_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12145_ _06403_ _06404_ _06402_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__o21ai_1
X_12076_ datapath.mulitply_result\[16\] datapath.multiplication_module.multiplicand_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
X_11027_ _05266_ _05271_ _05677_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__or3_2
XANTENNA__10679__B1 _05529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__A1 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12749__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ net248 net2295 net607 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ net154 _05881_ net129 screen.register.currentXbus\[15\] vssd1 vssd1 vccd1
+ vccd1 _00526_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12484__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ datapath.rf.registers\[17\]\[26\] net763 net756 datapath.rf.registers\[24\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a22o_1
XANTENNA__07075__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07051_ datapath.rf.registers\[29\]\[28\] net878 _01973_ _01975_ _01977_ vssd1 vssd1
+ vccd1 vccd1 _01978_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_140_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07783__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ net513 _02879_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__and2_1
X_06904_ net999 net985 net978 _01812_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__and4_4
X_07884_ net694 _02801_ _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__or3_1
XANTENNA__11331__A1 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ net318 _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__nand2_1
X_06835_ net997 _01754_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__and2_1
XANTENNA__11882__A2 _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12659__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06766_ datapath.ru.latched_instruction\[1\] _01587_ _01607_ datapath.ru.latched_instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ net421 _04480_ net318 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08505_ _02084_ _03428_ _03429_ _03362_ _02082_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__o311a_1
XANTENNA__07299__C1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06697_ mmio.memload_or_instruction\[14\] net1063 net1008 datapath.ru.latched_instruction\[14\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__a32o_4
X_09485_ net636 _04397_ _04408_ _04404_ net611 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout534_A _01950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08436_ _02105_ net531 vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11799__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08367_ datapath.rf.registers\[27\]\[0\] net868 _03289_ _03291_ _03293_ vssd1 vssd1
+ vccd1 vccd1 _03294_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__12394__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08799__C1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ datapath.rf.registers\[3\]\[22\] net966 net954 datapath.rf.registers\[22\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
X_08298_ datapath.rf.registers\[14\]\[1\] net995 _01752_ vssd1 vssd1 vccd1 vccd1 _03225_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10070__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ datapath.rf.registers\[20\]\[23\] net802 net731 datapath.rf.registers\[16\]\[23\]
+ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10260_ net505 _03207_ net360 vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__mux2_1
XANTENNA__06556__C_N mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ _05116_ _05117_ net1056 vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1305 net1307 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout340 _03509_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_2
Xfanout351 _05332_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_2
X_13950_ clknet_leaf_50_clk _00837_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout373 _03538_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_2
Xfanout384 net387 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_2
XANTENNA__07526__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11322__B2 _01464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net397 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_2
X_12901_ net1671 net292 net548 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
XANTENNA__12569__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13831__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ clknet_leaf_60_clk _00768_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12832_ net180 net1745 net556 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12763_ net168 net2274 net567 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14502_ clknet_leaf_106_clk _01389_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11714_ net1296 net663 _06149_ net712 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12694_ net1874 net188 net434 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14433_ clknet_leaf_41_clk _01320_ net1162 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11645_ net666 _06103_ _06105_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07057__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ clknet_leaf_54_clk _01251_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11576_ net1012 _06032_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a21o_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput37 gpio_in[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XFILLER_0_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13315_ clknet_leaf_110_clk _00305_ net1103 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_10527_ _05431_ _05432_ _05435_ _05399_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__o221a_1
X_14295_ clknet_leaf_45_clk _01182_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ clknet_leaf_75_clk _00236_ net1251 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
X_10458_ net527 net526 net524 _02389_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10389_ net1288 net1283 net1279 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__or3_1
X_13177_ clknet_leaf_48_clk _00169_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07765__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ net323 _06390_ _06391_ net327 net1820 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a32o_1
X_12059_ _06331_ _06332_ _06330_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_127_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07517__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A1 datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06620_ _01493_ _01497_ _01547_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06740__A1 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06551_ net1305 net1303 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ _01481_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_47_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09270_ net320 _03841_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06482_ datapath.ru.latched_instruction\[13\] vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
XANTENNA__07296__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08221_ datapath.rf.registers\[0\]\[2\] net827 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_60_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08152_ datapath.rf.registers\[11\]\[3\] net969 net857 datapath.rf.registers\[15\]\[3\]
+ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a221o_1
XANTENNA__07048__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10052__A1 _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ datapath.rf.registers\[31\]\[27\] net950 net946 datapath.rf.registers\[19\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ datapath.rf.registers\[6\]\[5\] net813 net774 datapath.rf.registers\[11\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12942__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07034_ datapath.rf.registers\[24\]\[28\] net756 net752 datapath.rf.registers\[22\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07756__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _01633_ net688 net492 vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout484_A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ datapath.rf.registers\[22\]\[8\] net754 net745 datapath.rf.registers\[21\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a22o_1
XANTENNA__12389__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ datapath.rf.registers\[16\]\[9\] net962 net897 datapath.rf.registers\[6\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__a22o_1
XANTENNA__08181__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09606_ net339 _04399_ net315 vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06818_ datapath.rf.registers\[7\]\[31\] net825 net821 datapath.rf.registers\[26\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a22o_1
X_07798_ datapath.rf.registers\[12\]\[11\] net888 net860 datapath.rf.registers\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XANTENNA__06731__A1 _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net654 _04459_ _04461_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or4b_1
XFILLER_0_149_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06749_ _01672_ _01674_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout916_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09130__C1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ _02764_ _02786_ net683 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08419_ _02085_ _02127_ _03343_ _02081_ _02039_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o311a_1
X_09399_ net403 _03992_ _04325_ net336 vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07039__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11430_ _05716_ _05809_ _05813_ net1293 vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08334__C _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11361_ _03285_ net669 vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__and2_1
XANTENNA__11240__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07995__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ net1278 _04278_ net536 vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__mux2_1
X_13100_ clknet_leaf_30_clk _00092_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11292_ net12 net1046 net1035 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1
+ vccd1 _00306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14080_ clknet_leaf_46_clk _00967_ net1195 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10243_ net1278 datapath.PC\[3\] vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__xor2_1
X_13031_ clknet_leaf_25_clk _00023_ net1144 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07747__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1125 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_2
X_10174_ net203 _05096_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__or3_1
XANTENNA__07211__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 net1115 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_4
Xfanout1124 net1125 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_2
Xfanout1135 net1200 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_2
Xfanout1146 net1149 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_4
Xfanout1157 net1158 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_4
Xfanout1168 net1171 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout170 _05569_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_2
Xfanout181 net183 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_2
Xfanout192 _05544_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
X_13933_ clknet_leaf_119_clk _00820_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12299__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__B _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864_ clknet_leaf_105_clk _00751_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12815_ net240 net2633 net559 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13795_ clknet_leaf_107_clk _00682_ net1110 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10806__B1 _05636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12746_ net254 net2105 net565 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__mux2_1
XANTENNA__07278__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09401__S net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12677_ net2565 net265 net431 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14416_ clknet_leaf_3_clk _01303_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11628_ screen.counter.currentCt\[13\] screen.counter.currentCt\[12\] screen.counter.currentCt\[15\]
+ screen.counter.currentCt\[14\] vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09424__B1 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11231__B1 _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ clknet_leaf_68_clk _01234_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12762__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11559_ screen.register.currentXbus\[7\] _05720_ _05735_ screen.register.currentYbus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 datapath.mulitply_result\[26\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 datapath.rf.registers\[20\]\[22\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 datapath.rf.registers\[12\]\[10\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ clknet_leaf_106_clk _01165_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07450__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09188__C1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13229_ clknet_leaf_90_clk _00220_ net1211 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11534__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07202__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ net706 _03638_ net623 vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__a21o_1
X_07721_ datapath.rf.registers\[23\]\[13\] net932 net888 datapath.rf.registers\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XANTENNA__11298__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11407__A _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ datapath.rf.registers\[2\]\[14\] net726 net722 datapath.rf.registers\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XANTENNA__06713__A1 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09522__D _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06603_ datapath.ru.latched_instruction\[19\] _01494_ _01507_ datapath.ru.latched_instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07583_ datapath.rf.registers\[10\]\[16\] net918 net850 datapath.rf.registers\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12937__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06534_ mmio.key_data\[1\] mmio.memload_or_instruction\[1\] net1060 vssd1 vssd1 vccd1
+ vccd1 _01464_ sky130_fd_sc_hd__mux2_2
X_09322_ net370 _04129_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or2_1
XANTENNA__07269__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__B1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09253_ _04175_ _04179_ net402 vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08435__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ datapath.rf.registers\[6\]\[2\] net899 net884 datapath.rf.registers\[9\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09184_ _04103_ _04105_ _03505_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08135_ net647 _03060_ _03041_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12672__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ datapath.rf.registers\[8\]\[5\] net925 net884 datapath.rf.registers\[9\]\[5\]
+ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a221o_1
XANTENNA__07441__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ datapath.rf.registers\[4\]\[29\] net931 net927 datapath.rf.registers\[8\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nand2_1
X_07919_ datapath.rf.registers\[8\]\[8\] net925 net851 datapath.rf.registers\[1\]\[8\]
+ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__a221o_1
XANTENNA__11828__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08154__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ net707 _03786_ net623 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_3_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10930_ net294 net2160 net591 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07901__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ net295 net2296 net600 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12600_ _05575_ _05671_ _06445_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_27_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ clknet_leaf_89_clk _00530_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10792_ _04416_ _05624_ net844 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__mux2_2
XFILLER_0_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12531_ net1975 net171 net453 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12462_ net193 net2214 net461 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
X_14201_ clknet_leaf_47_clk _01088_ net1197 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ _02059_ net668 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__and2_1
XANTENNA__11213__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12582__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ net213 net2480 net469 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
XANTENNA__07968__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ clknet_leaf_115_clk _01019_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09457__A _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _01503_ net1027 net308 net312 datapath.ru.latched_instruction\[23\] vssd1
+ vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__a32o_1
XANTENNA__07432__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14063_ clknet_leaf_7_clk _00950_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11275_ net24 net1046 net1035 mmio.memload_or_instruction\[2\] vssd1 vssd1 vccd1
+ vccd1 _00289_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09185__A2 _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ clknet_leaf_24_clk _00006_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10226_ net204 _04804_ _05152_ net1309 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a31oi_1
X_10157_ _04081_ _04417_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__xor2_1
Xhold4 keypad.debounce.debounce\[11\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
X_10088_ net834 _03909_ _04449_ _04965_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__o311a_1
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08145__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13916_ clknet_leaf_58_clk _00803_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07499__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ clknet_leaf_45_clk _00734_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12757__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08448__A1 _02457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13778_ clknet_leaf_35_clk _00665_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12729_ net172 net2445 net572 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08255__B net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07671__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11204__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12492__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold404 datapath.rf.registers\[13\]\[19\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09367__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 datapath.mulitply_result\[4\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 datapath.rf.registers\[15\]\[14\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 datapath.rf.registers\[14\]\[25\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 datapath.rf.registers\[9\]\[7\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _04611_ net201 _04667_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a31oi_1
Xhold459 datapath.rf.registers\[13\]\[30\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ _04722_ _04747_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__xnor2_1
Xfanout917 net919 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_4
Xfanout928 _01820_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 _01817_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
XFILLER_0_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08822_ net415 _03603_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nor2_1
Xhold1104 datapath.rf.registers\[14\]\[31\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 datapath.rf.registers\[16\]\[6\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 datapath.rf.registers\[18\]\[18\] vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 datapath.rf.registers\[14\]\[10\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net497 net494 net529 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__a21o_1
Xhold1148 datapath.rf.registers\[0\]\[31\] vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout182_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09333__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _02617_ _02618_ _02625_ _02627_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__or4_1
XANTENNA__07334__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08684_ _03477_ _03479_ net409 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06698__A0 datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07635_ datapath.rf.registers\[22\]\[15\] net953 net870 datapath.rf.registers\[27\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
XANTENNA__12667__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1189_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ datapath.rf.registers\[11\]\[16\] net776 net764 datapath.rf.registers\[17\]\[16\]
+ _02492_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__a221o_1
XANTENNA__08446__A _02457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09305_ _04225_ _04227_ _04231_ _04194_ net674 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__o32a_2
X_06517_ columns.count\[5\] columns.count\[4\] vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07497_ _02418_ _02420_ _02422_ _02423_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ net399 _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07662__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10915__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ net382 _03887_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ datapath.rf.registers\[12\]\[4\] net736 net728 datapath.rf.registers\[2\]\[4\]
+ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__a221o_1
XANTENNA__08611__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ net502 net619 net496 net518 vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a211o_1
X_08049_ _02973_ net510 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07509__B _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13604__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold960 datapath.rf.registers\[7\]\[23\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 datapath.rf.registers\[27\]\[14\] vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _05698_ _05702_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__or2_1
Xhold982 datapath.rf.registers\[28\]\[31\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 datapath.rf.registers\[11\]\[15\] vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08375__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ datapath.PC\[25\] _04518_ net539 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__mux2_1
XANTENNA__10650__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08127__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07244__B _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ net247 net1742 net580 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13701_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[18\]
+ net1258 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ net217 net2552 net597 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__mux2_1
XANTENNA__12577__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ net1425 _05878_ net156 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14560__1333 vssd1 vssd1 vccd1 vccd1 _14560__1333/HI net1333 sky130_fd_sc_hd__conb_1
X_13632_ clknet_leaf_51_clk _00570_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10844_ net2081 net217 net604 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10237__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13563_ clknet_leaf_89_clk _00513_ net1231 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10775_ datapath.mulitply_result\[7\] net430 _05608_ _05611_ net659 vssd1 vssd1 vccd1
+ vccd1 _05612_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12514_ net2169 net257 net452 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13494_ clknet_leaf_80_clk net1372 net1239 vssd1 vssd1 vccd1 vccd1 screen.screenEdge.enable2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07653__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08850__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12445_ net272 net1852 net461 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XANTENNA__06861__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07405__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ _05607_ net2242 net468 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14115_ clknet_leaf_105_clk _01002_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11327_ datapath.ru.latched_instruction\[6\] net313 net309 _01582_ vssd1 vssd1 vccd1
+ vccd1 _00329_ sky130_fd_sc_hd__a22o_1
XANTENNA__13345__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07419__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14046_ clknet_leaf_53_clk _00933_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11258_ net1455 net140 net134 _02191_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08366__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ _04817_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_66_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11189_ mmio.key_data\[4\] net220 _05829_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_50_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08118__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09072__D _03998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07420_ _02324_ net524 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09618__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07351_ _02271_ _02275_ _02276_ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_75_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ datapath.rf.registers\[18\]\[23\] net914 net901 datapath.rf.registers\[20\]\[23\]
+ _02208_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07644__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09021_ _02567_ net687 net679 _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08054__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 datapath.rf.registers\[7\]\[0\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 datapath.rf.registers\[27\]\[1\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 datapath.rf.registers\[25\]\[30\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06604__B1 _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold234 net87 vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 datapath.rf.registers\[28\]\[1\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12950__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07329__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold256 datapath.rf.registers\[21\]\[25\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold267 datapath.rf.registers\[20\]\[2\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 datapath.rf.registers\[12\]\[21\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _04844_ _04847_ _04842_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__o21a_1
Xhold289 datapath.rf.registers\[30\]\[0\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 _01721_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_2
Xfanout714 screen.counter.ack vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_84_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout725 _01780_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
Xfanout736 _01777_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_4
X_09854_ datapath.PC\[21\] net629 _04672_ _04769_ vssd1 vssd1 vccd1 vccd1 _04781_
+ sky130_fd_sc_hd__a211oi_2
Xfanout747 _01773_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_4
Xfanout758 _01770_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_4
Xfanout769 _01766_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
X_08805_ net639 _03720_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a21bo_1
X_09785_ datapath.PC\[11\] net627 _04709_ _04710_ vssd1 vssd1 vccd1 vccd1 _04712_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_147_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08109__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ datapath.rf.registers\[4\]\[29\] net811 net747 datapath.rf.registers\[21\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ net414 _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08667_ net1057 _03593_ net705 vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout731_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ datapath.rf.registers\[0\]\[15\] net828 _02544_ vssd1 vssd1 vccd1 vccd1 _02545_
+ sky130_fd_sc_hd__o21ai_2
XANTENNA__09609__B1 _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08598_ _03288_ _03507_ _01861_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10219__A1 _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ datapath.rf.registers\[0\]\[17\] net690 _02463_ _02475_ vssd1 vssd1 vccd1
+ vccd1 _02476_ sky130_fd_sc_hd__o22a_4
XFILLER_0_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07096__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net1050 _05467_ keypad.alpha vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__mux2_1
XANTENNA__07635__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ net379 _04132_ _04145_ net332 vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _05399_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net184 net2543 net575 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08342__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12860__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ datapath.mulitply_result\[30\] datapath.multiplication_module.multiplicand_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08060__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11112_ net1023 _05731_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12092_ net321 _06360_ _06361_ net325 net1967 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_112_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold790 datapath.rf.registers\[23\]\[8\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _05313_ _05322_ _05684_ _05693_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__and4_1
XANTENNA__07020__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_12994_ net1409 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__clkbuf_1
X_11945_ net153 _05897_ net128 net2606 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876_ datapath.PC\[1\] net177 _06261_ _05183_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__o22a_1
XANTENNA__07874__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13615_ clknet_leaf_1_clk _00553_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10827_ net841 _03946_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13546_ clknet_leaf_88_clk _00496_ net1209 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ net839 _04336_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__nand2_1
XANTENNA__07626__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13477_ clknet_leaf_83_clk _00430_ net1237 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10689_ datapath.PC\[26\] _05532_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12428_ net1710 net196 net466 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08587__A0 _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12770__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ net2147 net218 net474 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14029_ clknet_leaf_118_clk _00916_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_06920_ net1000 net983 net980 _01801_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__and4_1
XANTENNA__07011__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11894__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ _01731_ _01758_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__and2_1
XANTENNA__10303__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09570_ _04475_ _04477_ _04495_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__or3_1
X_06782_ _01410_ net1009 _01582_ _01671_ _01708_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08521_ _03444_ _03447_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__and2_2
XFILLER_0_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11415__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08452_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07403_ datapath.rf.registers\[5\]\[20\] net854 _02325_ _02327_ _02329_ vssd1 vssd1
+ vccd1 vccd1 _02330_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_148_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12945__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _03288_ _03307_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout145_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07078__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07334_ datapath.rf.registers\[0\]\[21\] net828 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07265_ net652 _02191_ net627 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout312_A _05859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08443__B _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ net522 net356 _03930_ net385 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07196_ datapath.rf.registers\[17\]\[25\] net882 net859 datapath.rf.registers\[15\]\[25\]
+ _02122_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a221o_1
XANTENNA__12680__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1221_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout681_A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
XANTENNA_fanout779_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _02951_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_2
X_09906_ _04780_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__and2_1
Xfanout522 _02476_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_4
Xfanout533 _01991_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
Xfanout544 _06471_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_8
Xfanout566 _06465_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_4
Xfanout577 _06445_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
X_09837_ _04688_ _04691_ _04762_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__or3_1
Xfanout588 net589 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_8
Xfanout599 _05668_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14055__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ net632 _04694_ datapath.PC\[15\] vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__o21a_1
X_08719_ _03642_ _03645_ net413 vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _04586_ _04625_ _03504_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11730_ screen.counter.ct\[10\] net663 _06159_ net712 vssd1 vssd1 vccd1 vccd1 _00433_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08337__C _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11661_ screen.counter.currentCt\[8\] _06114_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__and2_1
XANTENNA__12855__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13400_ clknet_leaf_77_clk _00001_ net1246 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10612_ net1490 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[24\]
+ sky130_fd_sc_hd__and2_1
X_14380_ clknet_leaf_30_clk _01267_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08805__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ net1293 _05752_ _06055_ net1292 vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_12_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13331_ clknet_leaf_95_clk net1302 net1218 vssd1 vssd1 vccd1 vccd1 mmio.key_en3 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ _05432_ _05443_ _05452_ _05397_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13262_ clknet_leaf_63_clk _00252_ net1271 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ screen.register.currentYbus\[1\] screen.register.currentYbus\[0\] screen.register.currentYbus\[3\]
+ screen.register.currentYbus\[2\] vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_114_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12213_ net262 net2521 net573 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12590__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08033__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ clknet_leaf_12_clk _00185_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12144_ _06402_ _06403_ _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_94_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12075_ datapath.mulitply_result\[16\] datapath.multiplication_module.multiplicand_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nand2_1
X_11026_ _05269_ _05270_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12977_ net251 net1709 net606 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ net154 _05880_ net129 net2483 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__a22o_1
XANTENNA__07847__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ _05552_ net176 _06249_ net179 vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10603__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13529_ clknet_leaf_86_clk _00479_ net1232 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11800__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08272__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07050_ datapath.rf.registers\[17\]\[28\] net881 net853 datapath.rf.registers\[5\]\[28\]
+ _01976_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a221o_1
XANTENNA__07480__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__08024__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_140_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07232__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08980__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ net650 _02875_ _02878_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a21oi_1
X_06903_ net999 net985 net978 net976 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__and4_4
X_07883_ _02803_ _02805_ _02807_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or4_1
X_09622_ _03834_ _04548_ net418 vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__mux2_1
X_06834_ net996 _01733_ _01735_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__and3_2
X_09553_ _04452_ _04479_ net411 vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06765_ datapath.ru.latched_instruction\[23\] _01656_ _01690_ _01691_ vssd1 vssd1
+ vccd1 vccd1 _01692_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_65_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08504_ _02084_ _03428_ _03429_ _02082_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__o31a_1
XANTENNA__07838__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _03321_ net613 _04388_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06696_ mmio.memload_or_instruction\[14\] net1063 net1008 datapath.ru.latched_instruction\[14\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08435_ _02019_ net532 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12675__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A _02255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ datapath.rf.registers\[4\]\[0\] net929 net895 datapath.rf.registers\[14\]\[0\]
+ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__a221o_1
XANTENNA__11799__B _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14577__1347 vssd1 vssd1 vccd1 vccd1 _14577__1347/HI net1347 sky130_fd_sc_hd__conb_1
XFILLER_0_151_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07317_ datapath.rf.registers\[2\]\[22\] net922 net854 datapath.rf.registers\[5\]\[22\]
+ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a221o_1
X_08297_ datapath.rf.registers\[12\]\[1\] net996 _01776_ vssd1 vssd1 vccd1 vccd1 _03224_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08263__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07471__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ datapath.rf.registers\[7\]\[23\] net826 net720 datapath.rf.registers\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout896_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08015__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ net648 _02104_ net626 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07223__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ net1276 _03576_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_76_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1306 mmio.key_en3 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__clkbuf_2
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_2
Xfanout341 _03456_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
Xfanout385 net387 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
X_12900_ net2076 net300 net548 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13880_ clknet_leaf_39_clk _00767_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08629__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ net631 _06451_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ net174 net2377 net568 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__mux2_1
XANTENNA__07829__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ clknet_leaf_95_clk _01388_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ net1296 _05715_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12585__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12693_ net1813 net194 net433 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__mux2_1
X_14432_ clknet_leaf_50_clk _01319_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11644_ _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14363_ clknet_leaf_52_clk _01250_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_30_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ _06038_ _06039_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nand2_1
XANTENNA__09451__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ clknet_leaf_110_clk _00304_ net1103 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput38 gpio_in[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_96_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10526_ net1048 _05404_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__or3_1
X_14294_ clknet_leaf_9_clk _01181_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13245_ clknet_leaf_75_clk _00235_ net1250 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08006__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ _05362_ _05363_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__or3_1
XANTENNA__10833__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06637__A_N mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07214__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ clknet_leaf_42_clk _00168_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10388_ net1292 net1285 _05299_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__o21a_1
XANTENNA__06568__A2 _01456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _06382_ _06389_ _06388_ _06387_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__o211ai_2
X_12058_ _06330_ _06331_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_127_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08714__A0 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11009_ net234 net2415 net582 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06550_ net1306 net1302 mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ _01480_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_47_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06481_ datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XANTENNA__12495__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ net847 _01644_ _01726_ _01639_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ datapath.rf.registers\[23\]\[3\] net935 net891 datapath.rf.registers\[12\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__a22o_1
XANTENNA__09978__C1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07102_ datapath.rf.registers\[21\]\[27\] net938 net882 datapath.rf.registers\[17\]\[27\]
+ _02028_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10052__A2 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08082_ _03002_ _03004_ _03006_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07033_ datapath.rf.registers\[26\]\[28\] net821 net775 datapath.rf.registers\[11\]\[28\]
+ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07205__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08984_ net655 _01633_ net641 net675 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07935_ _02860_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout477_A _06452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__inv_2
X_09605_ _03530_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or2_1
X_06817_ net987 _01743_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07797_ datapath.rf.registers\[10\]\[11\] net916 net880 datapath.rf.registers\[17\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XANTENNA__08168__B _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ net315 _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__or2_1
X_06748_ datapath.ru.latched_instruction\[17\] net1037 vssd1 vssd1 vccd1 vccd1 _01675_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ net420 _04392_ _04393_ net319 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__o211ai_2
X_06679_ mmio.memload_or_instruction\[30\] net1063 net1010 datapath.ru.latched_instruction\[30\]
+ net1040 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a32oi_4
XANTENNA_fanout811_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout909_A _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08418_ _02085_ _02127_ _03343_ _02081_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o31a_1
XANTENNA__07692__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ net392 _04100_ _04324_ net400 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08349_ datapath.rf.registers\[30\]\[0\] net990 _01752_ net974 _01731_ vssd1 vssd1
+ vccd1 vccd1 _03276_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11360_ _05260_ _05689_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_78_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07444__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__A2 _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__B2 _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ net844 _04661_ _04788_ net835 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__o211ai_2
XANTENNA__10653__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ net11 net1046 net1035 mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1
+ vccd1 _00305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13030_ clknet_leaf_114_clk _00022_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07528__A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ net699 _04278_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1103 net1105 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
X_10173_ net1054 _05097_ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a21oi_1
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
Xfanout1125 _00004_ vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
Xfanout1136 net1144 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input38_A gpio_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1149 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
Xfanout160 _05261_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10889__A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1158 net1163 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_2
Xfanout171 net174 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
Xfanout1169 net1171 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06970__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout193 _05544_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_1
X_13932_ clknet_leaf_31_clk _00819_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13863_ clknet_leaf_15_clk _00750_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12814_ net247 net2604 net558 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13794_ clknet_leaf_43_clk _00681_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10806__A1 _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10267__C1 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12745_ net257 net1739 net565 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12676_ net1617 net271 net433 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14415_ clknet_leaf_6_clk _01302_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11627_ screen.counter.currentCt\[0\] screen.counter.currentCt\[3\] screen.counter.currentCt\[2\]
+ screen.counter.currentCt\[1\] vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__or4b_1
XFILLER_0_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14346_ clknet_leaf_9_clk _01233_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07435__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ net1011 _06023_ _06006_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__a21o_1
Xhold608 datapath.rf.registers\[4\]\[12\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _05407_ _05419_ _05396_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__a21oi_1
X_14277_ clknet_leaf_107_clk _01164_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold619 datapath.rf.registers\[8\]\[15\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ screen.register.currentYbus\[11\] _05736_ _05955_ _05958_ vssd1 vssd1 vccd1
+ vccd1 _05959_ sky130_fd_sc_hd__a211o_1
X_13228_ clknet_leaf_88_clk _00219_ net1212 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13159_ clknet_leaf_10_clk _00151_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07157__B _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06961__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ datapath.rf.registers\[25\]\[13\] net872 net852 datapath.rf.registers\[5\]\[13\]
+ _02637_ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a221o_1
X_14576__1346 vssd1 vssd1 vccd1 vccd1 _14576__1346/HI net1346 sky130_fd_sc_hd__conb_1
XANTENNA__11298__B2 mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11407__B _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ datapath.rf.registers\[19\]\[14\] net759 net755 datapath.rf.registers\[24\]\[14\]
+ _02576_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06602_ _01465_ _01471_ _01506_ _01531_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__or4_1
X_07582_ datapath.rf.registers\[22\]\[16\] net954 net866 datapath.rf.registers\[13\]\[16\]
+ _02508_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09321_ net369 _04150_ _04246_ net378 vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__o211a_1
X_06533_ datapath.ru.latched_instruction\[28\] _01460_ _01462_ datapath.ru.latched_instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__o22a_1
XANTENNA__11423__A _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _04176_ _04178_ net395 vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07674__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08856__A1_N net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ datapath.rf.registers\[12\]\[2\] net891 net867 datapath.rf.registers\[13\]\[2\]
+ _03129_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a221o_1
XANTENNA__09415__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09183_ _02835_ net683 _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__o21a_1
XANTENNA__12953__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_A _05512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ net646 _03060_ _03041_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__o21a_1
XANTENNA__07426__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11773__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ datapath.rf.registers\[27\]\[5\] net869 net851 datapath.rf.registers\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07016_ datapath.rf.registers\[22\]\[29\] net954 net850 datapath.rf.registers\[1\]\[29\]
+ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout594_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1242_A mmio.memload_or_instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07067__B _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ net524 net355 _03855_ net390 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06952__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ datapath.rf.registers\[16\]\[8\] net961 net861 datapath.rf.registers\[28\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__a22o_1
X_08898_ _01717_ _03824_ net493 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a21o_1
X_07849_ datapath.rf.registers\[26\]\[10\] net820 net770 datapath.rf.registers\[30\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a22o_1
X_10860_ _05590_ net1552 net599 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ net675 _04440_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_27_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10791_ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__inv_2
XANTENNA__08626__B _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ net1893 net186 net454 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07665__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08345__C _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12461_ net198 net2199 net462 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
XANTENNA__08209__A2 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14200_ clknet_leaf_39_clk _01087_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11412_ screen.register.currentYbus\[25\] net131 _05891_ net160 vssd1 vssd1 vccd1
+ vccd1 _00383_ sky130_fd_sc_hd__a22o_1
XANTENNA__10016__A2 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net219 net2086 net470 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14131_ clknet_leaf_48_clk _01018_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11343_ _01485_ net1027 net308 net312 datapath.ru.latched_instruction\[22\] vssd1
+ vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_104_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14062_ clknet_leaf_116_clk _00949_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11274_ net13 net1047 net1036 mmio.memload_or_instruction\[1\] vssd1 vssd1 vccd1
+ vccd1 _00288_ sky130_fd_sc_hd__a22o_1
XANTENNA__11516__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ clknet_leaf_28_clk _00005_ net1130 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ _04801_ _04803_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__or2_1
XANTENNA__07196__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ _04808_ _05082_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06943__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 screen.counter.ack1 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ net1054 _05013_ _05012_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a21o_1
XANTENNA__08089__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06569__C_N mmio.memload_or_instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13915_ clknet_leaf_55_clk _00802_ net1175 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_113_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13846_ clknet_leaf_25_clk _00733_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13777_ clknet_leaf_7_clk _00664_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10989_ net167 net2376 net588 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10255__A2 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12728_ net187 net2102 net571 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__mux2_1
XANTENNA__07120__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12773__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12659_ net198 net1803 net438 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07408__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold405 datapath.rf.registers\[7\]\[10\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08081__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14329_ clknet_leaf_47_clk _01216_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold416 datapath.rf.registers\[13\]\[12\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 datapath.rf.registers\[14\]\[2\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold438 datapath.mulitply_result\[11\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold449 datapath.rf.registers\[14\]\[19\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout907 _01833_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _04792_ _04794_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_55_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_4
XANTENNA__09030__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10715__B1 _05560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout929 _01820_ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_2
XANTENNA__07187__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09383__A _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ _02303_ _02304_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__nor2_2
XANTENNA__09581__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 datapath.rf.registers\[20\]\[27\] vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 datapath.rf.registers\[9\]\[23\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net502 net618 _03543_ net531 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a211o_1
Xhold1127 datapath.rf.registers\[12\]\[29\] vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 datapath.rf.registers\[24\]\[4\] vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 datapath.rf.registers\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ datapath.rf.registers\[3\]\[13\] net766 net765 datapath.rf.registers\[17\]\[13\]
+ _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a221o_1
X_08683_ _01952_ net681 net678 _03596_ _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o221a_1
XANTENNA__12948__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10041__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06698__A1 _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ datapath.rf.registers\[3\]\[15\] net965 net897 datapath.rf.registers\[6\]\[15\]
+ _02560_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a221o_1
XANTENNA__07895__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ datapath.rf.registers\[14\]\[16\] net801 net794 datapath.rf.registers\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09304_ net638 _04209_ _04223_ _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__o211a_1
X_06516_ columns.count\[1\] columns.count\[3\] columns.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _01448_ sky130_fd_sc_hd__nand3_1
XANTENNA__07647__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ datapath.rf.registers\[2\]\[18\] net921 net873 datapath.rf.registers\[25\]\[18\]
+ _02421_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07111__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__C _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ net396 _04160_ _04161_ _04159_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__a31o_1
XANTENNA__12683__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout607_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09166_ net381 _03884_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nand2_1
X_08117_ datapath.rf.registers\[20\]\[4\] net802 net752 datapath.rf.registers\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08072__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09097_ net498 net495 _02608_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08611__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ net510 _02973_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold950 datapath.rf.registers\[5\]\[21\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 datapath.rf.registers\[14\]\[15\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 datapath.rf.registers\[29\]\[18\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10931__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold983 datapath.rf.registers\[3\]\[28\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 datapath.rf.registers\[28\]\[2\] vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07178__A2 _02104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ net1057 _03587_ _04936_ net845 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a31o_1
X_09999_ _01432_ _03584_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__nor2_1
XANTENNA__06925__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11961_ net251 net2589 net578 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__mux2_1
XANTENNA__12858__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ clknet_leaf_68_clk datapath.multiplication_module.multiplicand_i_n\[17\]
+ net1258 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10912_ net223 net2285 net596 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07886__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net1467 _05877_ net156 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
XANTENNA__07350__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ clknet_leaf_32_clk _00569_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10843_ net1779 net223 net603 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13562_ clknet_leaf_89_clk _00512_ net1214 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ net841 _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07102__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ net2551 net261 net452 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13493_ clknet_leaf_80_clk screen.screenEdge.enableIn net1239 vssd1 vssd1 vccd1 vccd1
+ screen.screenEdge.enable1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12593__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ net274 net1981 net462 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14575__1345 vssd1 vssd1 vccd1 vccd1 _14575__1345/HI net1345 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_117_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08063__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ net283 net2558 net468 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11002__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14114_ clknet_leaf_51_clk _01001_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11326_ datapath.ru.latched_instruction\[5\] net313 net309 _01501_ vssd1 vssd1 vccd1
+ vccd1 _00328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07810__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10126__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ clknet_leaf_32_clk _00932_ net1139 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10841__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ _02234_ _05844_ net146 net1600 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_130_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07169__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _04812_ _04813_ _04816_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__a21o_1
X_11188_ net1566 _05828_ _05833_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__a21o_1
XANTENNA__10173__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _04795_ _04796_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_50_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12768__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ clknet_leaf_107_clk _00716_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ datapath.rf.registers\[15\]\[21\] net806 net738 datapath.rf.registers\[8\]\[21\]
+ _02263_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a221o_1
XANTENNA__07629__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07281_ datapath.rf.registers\[23\]\[23\] net933 net893 datapath.rf.registers\[14\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09020_ _03376_ _03377_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08282__A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold202 datapath.rf.registers\[13\]\[24\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold213 datapath.rf.registers\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 datapath.rf.registers\[21\]\[24\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10400__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 datapath.rf.registers\[13\]\[23\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 datapath.rf.registers\[5\]\[24\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 screen.counter.currentCt\[15\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold268 datapath.rf.registers\[11\]\[24\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09922_ _04837_ _04840_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__and3_1
Xhold279 datapath.rf.registers\[22\]\[9\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09003__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 _01721_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_2
XFILLER_0_111_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout715 _01783_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_4
Xfanout726 net729 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_8
Xfanout737 _01775_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
X_09853_ _04773_ _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__or2_1
XANTENNA__06530__A mmio.memload_or_instruction\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout748 _01772_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_8
Xfanout759 net762 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_A _05590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net337 _03730_ net315 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__o21bai_1
X_09784_ net627 _04709_ _04710_ datapath.PC\[11\] vssd1 vssd1 vccd1 vccd1 _04711_
+ sky130_fd_sc_hd__o31a_1
X_06996_ datapath.rf.registers\[5\]\[29\] net785 net741 datapath.rf.registers\[1\]\[29\]
+ _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a221o_1
XANTENNA__07580__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _03660_ _03661_ net409 vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__mux2_1
XANTENNA__12678__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ datapath.PC\[31\] _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07868__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ net832 _02535_ _02541_ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__or4_1
X_08597_ _03247_ _03507_ _03511_ _03521_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout724_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _02458_ _02459_ _02472_ _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_81_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10926__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ _02396_ _02399_ _02404_ _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__or4_1
X_09218_ _04139_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10490_ net121 net123 net124 net122 vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__or4b_2
XFILLER_0_63_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06705__A _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09149_ _04050_ _04051_ _04075_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__or3b_1
XANTENNA__09242__C1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07399__A2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ datapath.mulitply_result\[30\] datapath.multiplication_module.multiplicand_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__nand2_1
X_11111_ _05717_ _05719_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nand2_1
X_12091_ _06353_ _06359_ _06358_ _06357_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__o211ai_1
Xhold780 datapath.mulitply_result\[27\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 datapath.rf.registers\[4\]\[13\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net1292 net1285 _05692_ net1012 vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07571__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ net1828 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__clkbuf_1
X_11944_ net154 _05896_ net129 net2641 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__a22o_1
XANTENNA__08520__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ net835 _05208_ net177 vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13614_ clknet_leaf_32_clk _00552_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10826_ net1860 net246 net603 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13545_ clknet_leaf_88_clk _00495_ net1211 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10836__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ net1722 net295 net603 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13476_ clknet_leaf_83_clk _00429_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ datapath.PC\[26\] _05532_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08036__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ net1591 net209 net466 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08587__A1 _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ net2316 net225 net473 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11309_ net122 _05407_ _05851_ vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
X_12289_ net2315 net232 net483 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14028_ clknet_leaf_35_clk _00915_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_06850_ net995 _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_147_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07562__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire525_A _02323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ _01482_ _01498_ _01508_ _01707_ net1005 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__o41a_1
XFILLER_0_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12498__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06770__B1 _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _03061_ net992 _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_2
XANTENNA__08277__A datapath.rf.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07314__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ _02634_ _02655_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__nor2_1
XANTENNA__11415__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07402_ datapath.rf.registers\[7\]\[20\] net958 net922 datapath.rf.registers\[2\]\[20\]
+ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08382_ _03287_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07333_ _02258_ _02259_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_34_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08814__A2 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_A _05840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ datapath.rf.registers\[0\]\[23\] _02190_ net829 vssd1 vssd1 vccd1 vccd1 _02191_
+ sky130_fd_sc_hd__mux2_8
X_09003_ net500 net621 net488 net521 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08027__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12961__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ datapath.rf.registers\[31\]\[25\] net950 net915 datapath.rf.registers\[18\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout501 _03287_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 _02905_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
X_09905_ _04782_ _04829_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__and3_1
Xfanout523 _02389_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_4
Xfanout534 _01950_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
Xfanout545 net548 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout674_A _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 _06468_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11885__A1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ _04691_ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__or2_1
Xfanout567 _06465_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_8
Xfanout578 _06266_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_4
Xfanout589 _05674_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_4
XANTENNA_fanout841_A _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _01653_ _04678_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nor2_1
X_06979_ _01885_ _01904_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__nand2_1
X_14574__1344 vssd1 vssd1 vccd1 vccd1 _14574__1344/HI net1344 sky130_fd_sc_hd__conb_1
XANTENNA_fanout939_A _01817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ _03643_ _03644_ net410 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__mux2_1
X_09698_ _03598_ _04544_ _04565_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_83_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08649_ datapath.PC\[11\] _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__or2_1
X_11660_ net667 _06113_ _06115_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__and3_1
X_10611_ net1398 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[23\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__08266__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_115_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11591_ screen.counter.ct\[11\] net1288 net1281 net1287 vssd1 vssd1 vccd1 vccd1 _06055_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_135_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08634__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ clknet_leaf_78_clk mmio.WEN net1246 vssd1 vssd1 vccd1 vccd1 mmio.WEN1 sky130_fd_sc_hd__dfrtp_1
X_10542_ net1049 _05426_ _05439_ _05451_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08018__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ clknet_leaf_63_clk _00251_ net1271 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12871__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10473_ screen.register.currentYbus\[5\] screen.register.currentYbus\[4\] screen.register.currentYbus\[7\]
+ screen.register.currentYbus\[6\] vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_114_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08569__A1 datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12212_ net265 net2489 net573 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ clknet_leaf_14_clk _00184_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12143_ datapath.mulitply_result\[27\] datapath.multiplication_module.multiplicand_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07792__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ net322 _06345_ _06346_ net326 net1858 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__a32o_1
X_11025_ net1292 screen.counter.ct\[8\] net1287 net1288 vssd1 vssd1 vccd1 vccd1 _05676_
+ sky130_fd_sc_hd__or4_1
XANTENNA__07544__A2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12976_ net255 net2223 net606 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11927_ net154 _05879_ net129 screen.register.currentXbus\[13\] vssd1 vssd1 vccd1
+ vccd1 _00524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11950__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11858_ net836 _04848_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_106_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10809_ _05488_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__nor2_1
XANTENNA__08257__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_19 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14577_ net1347 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11789_ datapath.PC\[8\] net303 _06197_ _06199_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ clknet_leaf_80_clk net1500 net1239 vssd1 vssd1 vccd1 vccd1 screen.counter.currentEnable
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11800__A1 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08009__B1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12781__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ clknet_leaf_77_clk _00415_ net1247 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09206__C1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07783__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08980__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ net650 _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__nor2_1
XANTENNA__10119__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06991__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06902_ net969 _01804_ _01824_ net924 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ datapath.rf.registers\[10\]\[9\] net917 net905 datapath.rf.registers\[24\]\[9\]
+ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11867__B2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ net991 _01739_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__and2_2
X_09621_ _03478_ _03487_ net411 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_1
X_09552_ _03660_ _03665_ net341 vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__mux2_1
X_06764_ datapath.ru.latched_instruction\[19\] _01640_ _01679_ datapath.ru.latched_instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08503_ _03428_ _03429_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09483_ net625 _04389_ _04390_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06695_ _01591_ _01621_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__or2_1
XANTENNA__12956__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ _02019_ net532 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08365_ datapath.rf.registers\[26\]\[0\] net943 net864 datapath.rf.registers\[13\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__C1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11161__A _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08454__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ datapath.rf.registers\[16\]\[22\] net963 net902 datapath.rf.registers\[20\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a22o_1
X_08296_ datapath.rf.registers\[6\]\[1\] net816 _03220_ _03221_ _03222_ vssd1 vssd1
+ vccd1 vccd1 _03223_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_150_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08173__C _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ datapath.rf.registers\[26\]\[23\] net821 net771 datapath.rf.registers\[30\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12691__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ net648 _02104_ net626 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout791_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout889_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13442__SET_B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1307 mmio.key_en3 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_1
Xfanout320 _03483_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
Xfanout331 _03534_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_2
Xfanout353 net358 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_4
Xfanout364 _03541_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_2
Xfanout375 _03538_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07526__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_2
X_09819_ _04726_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand2_1
Xfanout397 _03518_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08629__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ net163 net2577 net558 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12866__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ net184 net1862 net567 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__mux2_1
X_14500_ clknet_leaf_17_clk _01387_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11712_ net1297 net663 _06148_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a21o_1
X_12692_ net1677 net198 net434 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14431_ clknet_leaf_38_clk _01318_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11643_ screen.counter.currentCt\[1\] screen.counter.currentCt\[2\] _06100_ vssd1
+ vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _05722_ _05788_ net1017 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__o21ai_1
X_14362_ clknet_leaf_52_clk _01249_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10597__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_13313_ clknet_leaf_112_clk _00303_ net1098 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_10525_ _05396_ _05435_ _05407_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__mux2_1
Xinput39 nrst vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ clknet_leaf_28_clk _01180_ net1130 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ clknet_leaf_76_clk _00234_ net1247 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
X_10456_ _05365_ _05366_ _05367_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ clknet_leaf_43_clk _00167_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10387_ _05299_ _05307_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__nand2_1
XANTENNA__11010__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ _06387_ _06388_ _06389_ _06382_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__a211o_1
XANTENNA__06973__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ datapath.mulitply_result\[13\] datapath.multiplication_module.multiplicand_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07517__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ net241 net2619 net584 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08190__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ net186 net2632 net543 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__mux2_1
XANTENNA__12776__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06480_ datapath.ru.latched_instruction\[9\] vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XANTENNA__10824__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__C1 _04353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ datapath.rf.registers\[24\]\[3\] net904 net877 datapath.rf.registers\[29\]\[3\]
+ _03076_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07101_ datapath.rf.registers\[4\]\[27\] net930 net879 datapath.rf.registers\[29\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ datapath.rf.registers\[16\]\[5\] net733 net726 datapath.rf.registers\[2\]\[5\]
+ _03007_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_155_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14573__1343 vssd1 vssd1 vccd1 vccd1 _14573__1343/HI net1343 sky130_fd_sc_hd__conb_1
X_07032_ datapath.rf.registers\[27\]\[28\] net723 net720 datapath.rf.registers\[28\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06803__A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06522__B datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07756__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ _02526_ _03413_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06964__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ datapath.rf.registers\[25\]\[8\] net798 net721 datapath.rf.registers\[28\]\[8\]
+ _02859_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a221o_1
X_07865_ net515 _02786_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08449__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ net332 net379 _04247_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__or3_1
X_06816_ _01638_ _01646_ net982 net977 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__and4_4
X_07796_ _02722_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08168__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06747_ datapath.ru.latched_instruction\[17\] net1037 vssd1 vssd1 vccd1 vccd1 _01674_
+ sky130_fd_sc_hd__and2_1
X_09535_ _04256_ _04257_ net339 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12686__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ net412 _04122_ net418 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06678_ datapath.ru.latched_instruction\[25\] net1040 _01604_ vssd1 vssd1 vccd1 vccd1
+ _01606_ sky130_fd_sc_hd__a21o_1
XANTENNA__07141__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08417_ _02085_ _02127_ _03343_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ _04322_ _04323_ net392 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout804_A _01751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08348_ datapath.rf.registers\[16\]\[0\] net733 _03261_ _03266_ _03271_ vssd1 vssd1
+ vccd1 vccd1 _03275_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10579__A1 _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10934__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _03203_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__nand2_2
XFILLER_0_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10310_ _05181_ _05211_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07995__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09296__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net10 net1046 net1035 mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1
+ vccd1 _00304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10241_ _05166_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07747__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ net1056 _03577_ _05098_ net701 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a31o_1
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_2
Xfanout1115 net1124 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_2
Xfanout1126 net1130 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_4
Xfanout1137 net1144 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_2
Xfanout150 _06264_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout1148 net1149 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout161 _05261_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout1159 net1163 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_4
Xfanout172 net174 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout183 _05579_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_2
X_13931_ clknet_leaf_56_clk _00818_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
X_13862_ clknet_leaf_114_clk _00749_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07380__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ net251 net1826 net557 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__mux2_1
XANTENNA__12596__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13793_ clknet_leaf_40_clk _00680_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10267__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12744_ net261 net1994 net565 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__mux2_1
XANTENNA__10806__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13339__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ net1630 net273 net432 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XANTENNA__11005__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14414_ clknet_leaf_116_clk _01301_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ screen.counter.currentCt\[5\] screen.counter.currentCt\[4\] screen.counter.currentCt\[7\]
+ screen.counter.currentCt\[6\] vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14345_ clknet_leaf_12_clk _01232_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11231__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ screen.register.currentXbus\[31\] _05700_ _05776_ screen.register.currentYbus\[15\]
+ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10844__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07986__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10508_ _05415_ _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__or3_1
Xhold609 datapath.rf.registers\[10\]\[29\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
X_11488_ screen.register.currentYbus\[27\] _05742_ _05956_ _05957_ vssd1 vssd1 vccd1
+ vccd1 _05958_ sky130_fd_sc_hd__a211o_1
X_14276_ clknet_leaf_14_clk _01163_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13227_ clknet_leaf_88_clk _00218_ net1212 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10439_ screen.register.currentXbus\[9\] screen.register.currentXbus\[8\] screen.register.currentXbus\[11\]
+ screen.register.currentXbus\[10\] vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__or4_1
XANTENNA_max_cap435_A _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ clknet_leaf_106_clk _00150_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10742__A1 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06946__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12109_ _06373_ _06374_ _06372_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__o21ai_1
X_13089_ clknet_leaf_45_clk _00081_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11298__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ datapath.rf.registers\[26\]\[14\] net820 net789 datapath.rf.registers\[18\]\[14\]
+ _02569_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07371__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ _01410_ _01457_ _01517_ _01523_ _01524_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07910__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ datapath.rf.registers\[19\]\[16\] net946 net922 datapath.rf.registers\[2\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a22o_1
X_09320_ net369 _04150_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__o21ai_1
X_06532_ net1306 net1302 mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ _01462_ sky130_fd_sc_hd__or3b_2
XFILLER_0_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07123__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__A2 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ net389 _03690_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__o21a_1
X_08202_ datapath.rf.registers\[7\]\[2\] net959 net869 datapath.rf.registers\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ net679 _04082_ _04107_ net317 _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__o221a_1
X_08133_ datapath.rf.registers\[0\]\[4\] net828 _03050_ _03059_ vssd1 vssd1 vccd1
+ vccd1 _03060_ sky130_fd_sc_hd__o22a_4
XANTENNA__10754__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout218_A _05519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08064_ _02984_ _02986_ _02988_ _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07015_ datapath.rf.registers\[16\]\[29\] net963 net890 datapath.rf.registers\[12\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10733__A1 _05234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _02431_ net354 _03892_ net386 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a211o_1
X_07917_ datapath.rf.registers\[22\]\[8\] net955 net867 datapath.rf.registers\[13\]\[8\]
+ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a221o_1
X_08897_ net656 _03799_ _03811_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_95_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08154__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09351__B2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ datapath.rf.registers\[28\]\[10\] net718 _02773_ _02774_ vssd1 vssd1 vccd1
+ vccd1 _02775_ sky130_fd_sc_hd__a211o_1
XANTENNA__07362__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10929__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ datapath.rf.registers\[15\]\[11\] net805 net751 datapath.rf.registers\[22\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09518_ _04421_ _04439_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10790_ _05486_ _05623_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__or2_1
XANTENNA__08195__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09449_ _03505_ _04371_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ net210 net1760 net462 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11411_ net424 net714 vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__nor2_1
XANTENNA__08614__A0 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11213__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ net222 net2400 net469 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11342_ mmio.memload_or_instruction\[21\] net1061 net307 net311 datapath.ru.latched_instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__a32o_1
XANTENNA__07968__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14130_ clknet_leaf_34_clk _01017_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14061_ clknet_leaf_119_clk _00948_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11273_ net2 net1044 net1033 net2616 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10224_ net833 _05148_ _05150_ net204 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a211o_1
X_13012_ net2514 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11921__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ _04805_ _04807_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 screen.screenEdge.enable1 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _01430_ _03909_ net537 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__mux2_1
XANTENNA__10412__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08145__A2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ clknet_leaf_23_clk _00801_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_14572__1342 vssd1 vssd1 vccd1 vccd1 _14572__1342/HI net1342 sky130_fd_sc_hd__conb_1
X_13845_ clknet_leaf_28_clk _00732_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10839__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13776_ clknet_leaf_4_clk _00663_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07105__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10988_ net174 net2001 net589 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12727_ net190 net2556 net572 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__mux2_1
XANTENNA__11452__A2 _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ net210 net1952 net438 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ screen.counter.ct\[13\] screen.counter.ct\[15\] net1289 _06071_ vssd1 vssd1
+ vccd1 vccd1 _06072_ sky130_fd_sc_hd__and4_1
XFILLER_0_154_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12589_ net1644 net224 net445 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_152_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14328_ clknet_leaf_40_clk _01215_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold406 datapath.rf.registers\[4\]\[30\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 datapath.rf.registers\[6\]\[18\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 datapath.rf.registers\[10\]\[24\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 datapath.rf.registers\[5\]\[30\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ clknet_leaf_48_clk _01146_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 _01831_ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_4
Xfanout919 _01827_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08384__A2 _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ net673 _03705_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09383__B _04277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 datapath.rf.registers\[2\]\[6\] vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 screen.register.currentXbus\[14\] vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 datapath.rf.registers\[3\]\[18\] vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _02080_ net359 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_77_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
Xhold1139 datapath.rf.registers\[14\]\[4\] vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_07702_ datapath.rf.registers\[4\]\[13\] net809 net740 datapath.rf.registers\[1\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a22o_1
X_08682_ _01951_ net685 vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__or2_1
XANTENNA__07344__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ datapath.rf.registers\[10\]\[15\] net917 net853 datapath.rf.registers\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_1
X_07564_ _02486_ _02488_ _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__or3_1
XANTENNA__09097__B1 _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06515_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09303_ net623 _04228_ _04229_ _04197_ net656 vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_24_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12964__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ datapath.rf.registers\[26\]\[18\] net941 net938 datapath.rf.registers\[21\]\[18\]
+ _02415_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09234_ net522 net356 _03930_ net389 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08743__A _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09165_ net372 _03982_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08116_ datapath.rf.registers\[31\]\[4\] _01747_ net743 datapath.rf.registers\[1\]\[4\]
+ _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a221o_1
X_09096_ net502 net618 net496 _02566_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08047_ net510 _02973_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__nand2_1
Xhold940 datapath.rf.registers\[23\]\[23\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold951 datapath.rf.registers\[30\]\[31\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 datapath.rf.registers\[13\]\[10\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold973 datapath.rf.registers\[11\]\[14\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold984 datapath.rf.registers\[1\]\[24\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 datapath.rf.registers\[26\]\[5\] vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A _01848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11903__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12204__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net538 _04496_ _04924_ net1057 vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a211o_1
XANTENNA__07583__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ net421 _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_68_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08127__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ net255 net2059 net578 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__mux2_1
XANTENNA__07335__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ net230 net2130 net597 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__mux2_1
X_11891_ net1475 _05876_ net156 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13630_ clknet_leaf_53_clk _00568_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09088__A0 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ net2407 net231 net603 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ clknet_leaf_86_clk _00511_ net1232 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11434__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12874__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _05484_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ net2114 net266 net452 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06872__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ clknet_leaf_80_clk _00445_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ net277 net2545 net460 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XANTENNA__06861__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12374_ net294 net1621 net469 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__mux2_1
XANTENNA__09260__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14113_ clknet_leaf_42_clk _01000_ net1162 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11325_ _01477_ net1029 net309 net313 datapath.ru.latched_instruction\[4\] vssd1
+ vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_10_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14044_ clknet_leaf_57_clk _00931_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11256_ net342 _05844_ net147 net2645 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06536__C_N mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06901__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08366__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ datapath.PC\[8\] net1253 _05130_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_
+ sky130_fd_sc_hd__o22a_1
X_11187_ mmio.key_data\[3\] net220 _05829_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__and3_1
X_10138_ net698 _05064_ _05062_ net203 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_59_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11953__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ net842 _04662_ _04826_ _04995_ net704 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a221oi_1
XANTENNA__07326__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13828_ clknet_leaf_14_clk _00715_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12784__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ clknet_leaf_37_clk _00646_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ datapath.rf.registers\[16\]\[23\] net962 net941 datapath.rf.registers\[26\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 datapath.rf.registers\[5\]\[1\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold214 net42 vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold225 datapath.rf.registers\[7\]\[24\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 datapath.rf.registers\[12\]\[4\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 datapath.rf.registers\[15\]\[5\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 datapath.rf.registers\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 datapath.rf.registers\[23\]\[0\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07907__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09921_ _04844_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06811__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 _01721_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_2
Xfanout716 _01783_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_4
X_09852_ _04671_ _04674_ _04772_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__and3_1
Xfanout727 net729 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_4
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
Xfanout749 _01772_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_4
XANTENNA__07565__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08803_ _03527_ _03729_ net401 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__mux2_1
XANTENNA__12959__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ _01650_ net672 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nor2_1
X_06995_ datapath.rf.registers\[13\]\[29\] net794 net739 datapath.rf.registers\[8\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout285_A _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08109__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _02431_ net522 net404 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__mux2_1
XANTENNA__07317__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08665_ datapath.PC\[30\] _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout452_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _02530_ _02531_ _02533_ _02542_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__or4_1
X_08596_ _03247_ _03507_ _03521_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08176__C _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07547_ datapath.rf.registers\[30\]\[17\] net908 net852 datapath.rf.registers\[5\]\[17\]
+ _02473_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a221o_1
XANTENNA__08817__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12694__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout717_A _01783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ datapath.rf.registers\[31\]\[18\] net818 net763 datapath.rf.registers\[17\]\[18\]
+ _02394_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a221o_1
XANTENNA__07096__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09217_ _03538_ _04140_ _04143_ net382 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09148_ net708 _04074_ net491 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06559__C_N mmio.memload_or_instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10942__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ _03999_ _04004_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o21ai_1
X_14571__1341 vssd1 vssd1 vccd1 vccd1 _14571__1341/HI net1341 sky130_fd_sc_hd__conb_1
X_11110_ net1296 net1295 _01437_ net1294 vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__or4_1
X_12090_ _06357_ _06358_ _06359_ _06353_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_141_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold770 datapath.rf.registers\[28\]\[29\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 datapath.rf.registers\[5\]\[22\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net1282 net1279 _05323_ _05324_ _05300_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a41o_1
XANTENNA__08348__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold792 datapath.rf.registers\[31\]\[12\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11352__A1 _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09751__B net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ net1996 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07308__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__A _02457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ net153 _05895_ net128 screen.register.currentXbus\[29\] vssd1 vssd1 vccd1
+ vccd1 _00540_ sky130_fd_sc_hd__a22o_1
XANTENNA__07859__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__A0 _05607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11874_ datapath.PC\[0\] _06260_ net177 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__mux2_1
X_13613_ clknet_leaf_56_clk _00551_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ _01461_ net710 _05652_ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__o22a_2
XANTENNA__08808__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13544_ clknet_leaf_96_clk _00494_ net1219 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10756_ _05594_ _05595_ _01477_ net710 vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__08383__A _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13475_ clknet_leaf_83_clk _00428_ net1237 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ net198 net1658 net608 vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__mux2_1
XANTENNA__11013__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ net2326 net216 net466 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09784__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11948__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12357_ net2089 net231 net474 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__mux2_1
XANTENNA__10852__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ net121 _05449_ _05851_ vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12288_ net1666 net227 net480 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14027_ clknet_leaf_101_clk _00914_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11239_ net1468 net141 net136 _03060_ vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__a22o_1
XANTENNA__07547__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07011__A2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06780_ net1028 _01705_ _01706_ _01474_ _01467_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08277__B net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ _02547_ net520 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nand2_1
X_07401_ datapath.rf.registers\[26\]\[20\] net942 net863 datapath.rf.registers\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08381_ datapath.rf.registers\[0\]\[0\] net691 net643 _03306_ vssd1 vssd1 vccd1 vccd1
+ _03308_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_147_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07332_ _02236_ _02255_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07078__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06806__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07263_ datapath.rf.registers\[9\]\[23\] net779 _02186_ _02188_ _02189_ vssd1 vssd1
+ vccd1 vccd1 _02190_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_155_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09002_ net500 net620 net488 _02431_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__o211a_1
X_07194_ datapath.rf.registers\[25\]\[25\] net874 net850 datapath.rf.registers\[1\]\[25\]
+ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout200_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07250__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ _04771_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__xnor2_1
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_2
Xfanout513 _02855_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 _02343_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07538__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout557 net560 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_8
X_09835_ _04693_ _04696_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__and3_1
XANTENNA__07002__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12689__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _06465_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_4
Xfanout579 _06266_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09571__B _03785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _04691_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__nor2_1
X_06978_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__inv_2
X_08717_ _03146_ _03207_ net407 vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09697_ _03638_ _04502_ _04521_ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_83_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__C1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ net1277 datapath.PC\[10\] _03574_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07710__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10937__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ net689 _03504_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__or2_2
XFILLER_0_92_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10610_ net2201 net345 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[22\]
+ sky130_fd_sc_hd__and2_1
X_11590_ net1290 net1291 net1285 screen.counter.ct\[10\] vssd1 vssd1 vccd1 vccd1 _06054_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_107_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ _05404_ _05413_ _05449_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13260_ clknet_leaf_63_clk _00250_ net1271 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10472_ mmio.wishbone.curr_state\[1\] _01434_ _05255_ mmio.wishbone.curr_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09215__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12211_ net270 net2609 net575 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
X_13191_ clknet_leaf_16_clk _00183_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07777__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12142_ datapath.mulitply_result\[27\] datapath.multiplication_module.multiplicand_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12073_ _06335_ _06340_ _06344_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__nand3_1
XANTENNA__11325__A1 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ net1396 _01442_ net1032 net1496 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__a22o_1
XANTENNA__11876__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12599__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ net259 net2108 net606 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__mux2_1
XANTENNA__11008__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11926_ net154 _05878_ net129 screen.register.currentXbus\[12\] vssd1 vssd1 vccd1
+ vccd1 _00523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ net705 _04584_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__nand2_1
XANTENNA__10847__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ net1276 _05487_ datapath.PC\[13\] vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a21oi_1
X_14576_ net1346 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
X_11788_ _05615_ net175 _06198_ net177 vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11261__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13527_ clknet_leaf_73_clk _00477_ net1245 vssd1 vssd1 vccd1 vccd1 datapath.PC\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10739_ datapath.mulitply_result\[1\] net426 _05580_ _05581_ net659 vssd1 vssd1 vccd1
+ vccd1 _05582_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ clknet_leaf_77_clk _00414_ net1247 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07480__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ net1861 net281 net464 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
X_13389_ clknet_leaf_109_clk net1387 net1202 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__07768__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__C1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07232__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07950_ _01612_ _01727_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nor2_1
X_06901_ net968 _01804_ _01824_ net924 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nor4_1
XANTENNA__11867__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ datapath.rf.registers\[22\]\[9\] net953 net901 datapath.rf.registers\[20\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a22o_1
X_09620_ net421 _03836_ _04052_ _03448_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o211ai_2
X_06832_ _01741_ net972 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__and2_1
XANTENNA__07940__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _02260_ _03338_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__xor2_1
X_06763_ datapath.ru.latched_instruction\[22\] _01638_ _01645_ datapath.ru.latched_instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08502_ _03366_ _03425_ _03367_ _02171_ _03364_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_19_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06694_ _01591_ _01621_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_65_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09482_ net638 _04408_ _04404_ net655 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07299__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14570__1340 vssd1 vssd1 vccd1 vccd1 _14570__1340/HI net1340 sky130_fd_sc_hd__conb_1
XFILLER_0_148_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08433_ _01931_ net534 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nor2_1
XANTENNA__10757__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout248_A _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ datapath.rf.registers\[11\]\[0\] net969 net909 datapath.rf.registers\[30\]\[0\]
+ _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11252__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ datapath.rf.registers\[26\]\[22\] net942 net931 datapath.rf.registers\[4\]\[22\]
+ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12972__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ datapath.rf.registers\[30\]\[1\] net992 _01752_ vssd1 vssd1 vccd1 vccd1 _03222_
+ sky130_fd_sc_hd__and3_1
X_07246_ datapath.rf.registers\[23\]\[23\] net788 net775 datapath.rf.registers\[11\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
XANTENNA__07471__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ datapath.rf.registers\[0\]\[25\] net829 _02098_ _02103_ vssd1 vssd1 vccd1
+ vccd1 _02104_ sky130_fd_sc_hd__o22ai_4
XANTENNA__07759__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__A2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout784_A _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1308 net72 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__buf_2
Xfanout310 _05860_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_2
Xfanout332 net333 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_2
Xfanout354 net358 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
Xfanout365 _03540_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_2
Xfanout376 net379 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
X_09818_ _04741_ _04743_ _04727_ _04729_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a211o_1
Xfanout387 _03523_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12212__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 _03515_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_2
XANTENNA__06734__A1 _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08198__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _04672_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_107_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ net188 net2171 net567 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _05715_ _06098_ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and3_1
X_12691_ net1606 net209 net434 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
X_14430_ clknet_leaf_50_clk _01317_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11642_ screen.counter.currentCt\[0\] screen.counter.currentCt\[1\] _06087_ screen.counter.currentCt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14361_ clknet_leaf_60_clk _01248_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12882__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11573_ _05304_ _05782_ _06031_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o211a_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_13312_ clknet_leaf_112_clk _00302_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ net1026 _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14292_ clknet_leaf_114_clk _01179_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07462__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ clknet_leaf_75_clk _00233_ net1250 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ _02368_ _05368_ _05369_ net423 vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4b_1
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ clknet_leaf_26_clk _00166_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07214__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10386_ _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__or2_1
XANTENNA__10415__B datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ _06377_ _06381_ _06383_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__a21oi_1
X_12056_ datapath.mulitply_result\[13\] datapath.multiplication_module.multiplicand_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_144_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11007_ net247 net1758 net584 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06725__A1 _01461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11961__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ net190 net2495 net542 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__mux2_1
XANTENNA__09675__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _05894_ _06263_ net149 net1464 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12889_ net209 net1590 net552 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14559_ net1332 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__12792__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07989__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ datapath.rf.registers\[8\]\[27\] net927 net859 datapath.rf.registers\[15\]\[27\]
+ _02026_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a221o_1
X_08080_ datapath.rf.registers\[23\]\[5\] net786 net734 datapath.rf.registers\[12\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a22o_1
XANTENNA__07453__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08571__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07031_ datapath.rf.registers\[18\]\[28\] net790 net779 datapath.rf.registers\[9\]\[28\]
+ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09386__B net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07205__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08982_ net672 _03906_ _03908_ _03903_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__o22a_2
XFILLER_0_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ datapath.rf.registers\[20\]\[8\] net803 _01760_ datapath.rf.registers\[23\]\[8\]
+ _02856_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout198_A _05537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _02790_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ net319 _04529_ _04525_ _04523_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06815_ _01639_ _01656_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__nor2_1
X_07795_ net652 _02721_ net627 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a21o_1
XANTENNA__12967__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _03540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ net637 _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__nor2_1
X_06746_ _01452_ _01577_ _01579_ _01480_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a211o_1
XANTENNA__09666__A0 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09465_ _04119_ _04391_ net412 vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__mux2_1
X_06677_ net1040 _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout532_A _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08416_ _02172_ _02214_ _03340_ _02169_ _02126_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__o311a_1
XANTENNA__07692__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ net390 _04211_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__or2_1
XANTENNA__11225__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ datapath.rf.registers\[21\]\[0\] net745 _03254_ _03262_ _03264_ vssd1 vssd1
+ vccd1 vccd1 _03274_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11776__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ datapath.rf.registers\[0\]\[1\] net693 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07444__A2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07229_ datapath.rf.registers\[11\]\[24\] net971 net874 datapath.rf.registers\[25\]\[24\]
+ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a221o_1
XANTENNA__09296__B _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12207__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10240_ _05123_ _05134_ _05145_ _05165_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_91_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10171_ net1276 _03576_ datapath.PC\[13\] vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10950__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1105 net1111 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1116 net1119 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_4
Xfanout1127 net1130 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
Xfanout140 net148 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout1138 net1144 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_4
Xfanout151 net155 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
Xfanout1149 net1164 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_2
Xfanout162 _05261_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
X_13930_ clknet_leaf_12_clk _00817_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_1
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_2
Xfanout195 _05544_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlymetal6s2s_1
X_13861_ clknet_leaf_95_clk _00748_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12877__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ net255 net1897 net557 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ clknet_leaf_46_clk _00679_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ net265 net2364 net565 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12674_ net2209 net279 net431 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
X_14413_ clknet_leaf_119_clk _01300_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11625_ screen.counter.currentEnable _06081_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06891__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ clknet_leaf_15_clk _01231_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09487__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__A_N net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire530 _02147_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_4
X_11556_ screen.register.currentXbus\[15\] _05709_ _06019_ _06021_ vssd1 vssd1 vccd1
+ vccd1 _06022_ sky130_fd_sc_hd__a211o_1
XANTENNA__07435__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ net1026 net1025 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14275_ clknet_leaf_105_clk _01162_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11487_ screen.register.currentXbus\[11\] net1016 net1014 screen.register.currentXbus\[19\]
+ _05734_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__a221o_1
XANTENNA__11021__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_90_clk _00217_ net1211 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10438_ screen.register.currentXbus\[13\] screen.register.currentXbus\[12\] screen.register.currentXbus\[15\]
+ screen.register.currentXbus\[14\] vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11956__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10860__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ clknet_leaf_109_clk _00149_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10369_ _05275_ _05276_ _05284_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__or3_1
X_12108_ _06372_ _06373_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__or3_1
X_13088_ clknet_leaf_46_clk _00080_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08148__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _06315_ _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nand2_1
XANTENNA__12787__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ datapath.ru.latched_instruction\[4\] _01476_ _01522_ _01529_ _01474_ vssd1
+ vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a2111oi_1
X_07580_ datapath.rf.registers\[7\]\[16\] net958 _02502_ _02504_ _02506_ vssd1 vssd1
+ vccd1 vccd1 _02507_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06531_ mmio.memload_or_instruction\[15\] net1058 vssd1 vssd1 vccd1 vccd1 _01461_
+ sky130_fd_sc_hd__and2_1
X_09250_ net528 net357 _03814_ net385 vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07674__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08201_ datapath.rf.registers\[19\]\[2\] net947 net877 datapath.rf.registers\[29\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11207__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09181_ _02836_ _03494_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__nand2_1
X_08132_ _03052_ _03054_ _03056_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07426__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06814__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ datapath.rf.registers\[4\]\[5\] net928 net860 datapath.rf.registers\[28\]\[5\]
+ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07014_ datapath.rf.registers\[31\]\[29\] net950 net946 datapath.rf.registers\[19\]\[29\]
+ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10770__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11265__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ net499 net620 net488 net522 vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout482_A _06449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ datapath.rf.registers\[18\]\[8\] net913 net895 datapath.rf.registers\[14\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08896_ net315 _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__or2_1
X_07847_ datapath.rf.registers\[24\]\[10\] net755 net740 datapath.rf.registers\[1\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__a22o_1
XANTENNA__12697__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ datapath.rf.registers\[8\]\[11\] net737 net718 datapath.rf.registers\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09517_ _04438_ _04441_ _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_104_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06729_ datapath.ru.latched_instruction\[23\] net1039 net1007 _01655_ vssd1 vssd1
+ vccd1 vccd1 _01656_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_149_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08195__B _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_A _01830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ _04372_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07665__A2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06873__B1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ net625 _04293_ _04294_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a31o_1
XANTENNA__10945__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11410_ net2630 net131 _05890_ net160 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ net230 net2023 net470 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ _01505_ net1028 net307 net311 datapath.ru.latched_instruction\[20\] vssd1
+ vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__a32o_1
XANTENNA__08090__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14060_ clknet_leaf_31_clk _00947_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ net1308 net1047 mmio.wishbone.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05848_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13011_ net1598 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__clkbuf_1
X_10223_ net700 _04386_ _05149_ _04385_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_18_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10680__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__B1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07050__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ _05048_ _05058_ _05069_ _05079_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__or4_1
Xhold7 screen.register.cFill1 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net1056 _03580_ _05011_ net702 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a31o_1
XANTENNA__09770__A _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13913_ clknet_leaf_48_clk _00800_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08550__A0 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13844_ clknet_leaf_115_clk _00731_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12400__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_27_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13775_ clknet_leaf_9_clk _00662_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ net185 net1719 net587 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__mux2_1
XANTENNA__11016__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12726_ net194 net2206 net571 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07656__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06864__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ net215 net2420 net437 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11608_ screen.counter.ct\[11\] screen.counter.ct\[10\] net1291 _06070_ vssd1 vssd1
+ vccd1 vccd1 _06071_ sky130_fd_sc_hd__and4_1
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07408__A2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ net1848 net231 net446 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ clknet_leaf_44_clk _01214_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11539_ _05978_ _05996_ net975 vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__or3b_1
XANTENNA__08081__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold407 datapath.rf.registers\[10\]\[21\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 mmio.wishbone.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 datapath.rf.registers\[30\]\[19\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ clknet_leaf_36_clk _01145_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_36_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08369__B1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ clknet_leaf_47_clk _00201_ net1196 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_14189_ clknet_leaf_119_clk _01076_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout909 _01831_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07041__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08384__A3 _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08750_ net532 net359 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__or2_1
Xhold1107 datapath.rf.registers\[10\]\[30\] vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 datapath.rf.registers\[26\]\[2\] vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 datapath.rf.registers\[23\]\[27\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ datapath.rf.registers\[20\]\[13\] net804 net751 datapath.rf.registers\[22\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08681_ _03448_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__nand2_1
XANTENNA__08541__A0 _02997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ datapath.rf.registers\[19\]\[15\] net945 net926 datapath.rf.registers\[8\]\[15\]
+ _02558_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a221o_1
XANTENNA__12310__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07895__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ datapath.rf.registers\[31\]\[16\] net819 net732 datapath.rf.registers\[16\]\[16\]
+ _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__a221o_1
XANTENNA__11979__A1 datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09302_ net689 _04193_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ columns.count\[9\] columns.count\[10\] _01445_ vssd1 vssd1 vccd1 vccd1 _01446_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07647__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ datapath.rf.registers\[7\]\[18\] net957 net910 datapath.rf.registers\[30\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ net385 _04014_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout230_A _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ net374 _04089_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06607__B1 _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08115_ datapath.rf.registers\[30\]\[4\] net773 net730 datapath.rf.registers\[16\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a22o_1
XANTENNA__12980__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08072__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ net339 _04021_ _04020_ _04019_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08002__A_N net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _02971_ _02972_ net646 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_2
XANTENNA__07280__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold930 datapath.rf.registers\[26\]\[4\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold941 datapath.rf.registers\[29\]\[6\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 datapath.rf.registers\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 datapath.rf.registers\[30\]\[14\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 datapath.rf.registers\[15\]\[12\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 datapath.rf.registers\[11\]\[3\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold996 datapath.rf.registers\[6\]\[31\] vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__CLK clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ datapath.PC\[22\] net538 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout864_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _03601_ _03612_ _03454_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__mux2_1
XANTENNA__09590__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ _03801_ _03802_ net368 vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__a21o_1
X_10910_ net226 net2055 net594 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__mux2_1
XANTENNA__12220__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _05875_ _06263_ net149 net1443 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10841_ net1659 net227 net603 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__mux2_1
XANTENNA__09088__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10487__D_N net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07099__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ clknet_leaf_79_clk _00510_ net1244 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ datapath.PC\[6\] _05483_ datapath.PC\[7\] vssd1 vssd1 vccd1 vccd1 _05609_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ net2037 net270 net454 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
X_13491_ clknet_leaf_80_clk _00444_ net1239 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12442_ net280 net2530 net460 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12373_ net292 net2444 net471 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__mux2_1
XANTENNA__08063__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14112_ clknet_leaf_48_clk _00999_ net1195 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11324_ datapath.ru.latched_instruction\[3\] net313 net309 _01456_ vssd1 vssd1 vccd1
+ vccd1 _00326_ sky130_fd_sc_hd__a22o_1
XANTENNA__07271__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14043_ clknet_leaf_21_clk _00930_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09484__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11255_ net525 _05844_ net147 net2648 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__a2bb2o_1
X_10206_ net204 _05132_ net1310 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a21o_1
X_11186_ net1400 _05828_ _05832_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__a21o_1
X_10137_ _04338_ _05063_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ _04784_ _04822_ _04825_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08523__A0 _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__A datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ clknet_leaf_104_clk _00714_ net1121 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ clknet_leaf_49_clk _00645_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07629__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ net271 net1932 net571 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10585__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[6\] net1224
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08054__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold204 datapath.rf.registers\[10\]\[4\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 datapath.rf.registers\[15\]\[0\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 datapath.rf.registers\[29\]\[3\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold237 datapath.rf.registers\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 datapath.rf.registers\[25\]\[14\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _04773_ _04774_ _04846_ _04845_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold259 datapath.rf.registers\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12305__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06811__B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net708 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_2
XANTENNA__07014__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 _01783_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
X_09851_ _04776_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__or2_1
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
Xfanout739 _01775_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
XANTENNA__08762__A0 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08802_ net394 _03727_ _03728_ _03724_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a31o_1
X_09782_ net977 _04678_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06994_ datapath.rf.registers\[6\]\[29\] net815 net736 datapath.rf.registers\[12\]\[29\]
+ _01920_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a221o_1
X_08733_ net524 net523 net405 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_53_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout180_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08514__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout278_A _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__A1_N net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ datapath.PC\[29\] _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__or2_1
XANTENNA__07868__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ datapath.rf.registers\[17\]\[15\] net763 net723 datapath.rf.registers\[27\]\[15\]
+ _02534_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a221o_1
XANTENNA__12975__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _03247_ _03507_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout445_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ datapath.rf.registers\[25\]\[17\] net872 net864 datapath.rf.registers\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a22o_1
XANTENNA__08900__A1_N net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ datapath.rf.registers\[25\]\[18\] net797 net760 datapath.rf.registers\[19\]\[18\]
+ _02400_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ net366 _04141_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ net653 _04065_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07253__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ net613 _03997_ _04001_ _04003_ net491 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout981_A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ datapath.rf.registers\[7\]\[6\] net824 net740 datapath.rf.registers\[1\]\[6\]
+ _02954_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a221o_1
XANTENNA__12215__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07817__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold760 datapath.rf.registers\[28\]\[6\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06635__B_N mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold771 datapath.rf.registers\[10\]\[13\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 datapath.rf.registers\[14\]\[26\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07005__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _01440_ _05284_ _05348_ _05680_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_112_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold793 datapath.rf.registers\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08753__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ net1532 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07308__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ net153 _05894_ net128 screen.register.currentXbus\[28\] vssd1 vssd1 vccd1
+ vccd1 _00539_ sky130_fd_sc_hd__a22o_1
XANTENNA__07552__B net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__A2 _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12885__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ net203 _05212_ _05234_ net699 vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__a22o_1
X_13612_ clknet_leaf_10_clk _00550_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10824_ datapath.mulitply_result\[15\] net428 net662 vssd1 vssd1 vccd1 vccd1 _05653_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13543_ clknet_leaf_87_clk _00493_ net1220 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10755_ datapath.mulitply_result\[4\] net428 net662 vssd1 vssd1 vccd1 vccd1 _05595_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08383__B _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13474_ clknet_leaf_83_clk _00427_ net1237 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07492__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10686_ _01483_ net710 _05535_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__o22a_2
XFILLER_0_152_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12425_ net2440 net219 net466 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__mux2_1
XANTENNA__08036__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12356_ net1681 net226 net473 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__mux2_1
XANTENNA__06598__A2 _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _01449_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__nor2_4
XFILLER_0_121_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12287_ net2494 net242 net482 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14026_ clknet_leaf_8_clk _00913_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11238_ net1527 net142 net134 _03118_ vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11964__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _05806_ _05761_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_147_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12795__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07400_ datapath.rf.registers\[21\]\[20\] net939 net887 datapath.rf.registers\[9\]\[20\]
+ _02326_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ net643 _03306_ datapath.rf.registers\[0\]\[0\] net691 vssd1 vssd1 vccd1 vccd1
+ _03307_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07331_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06806__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07262_ _02176_ _02177_ _02183_ _02185_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ net657 _03927_ _03916_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__a21o_1
XANTENNA__08027__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07193_ datapath.rf.registers\[8\]\[25\] net927 net871 datapath.rf.registers\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07235__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09903_ _01432_ _01614_ _01727_ _04770_ _04781_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__o32a_1
Xfanout503 _03287_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout514 _02812_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11874__S net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ _04700_ _04702_ _04758_ _04698_ _04695_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a311o_1
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1102_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net560 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_4
Xfanout569 _06464_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_8
X_09765_ datapath.PC\[16\] net632 _04690_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__nor3_1
X_06977_ datapath.rf.registers\[0\]\[30\] net693 _01889_ _01903_ vssd1 vssd1 vccd1
+ vccd1 _01904_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout562_A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ net507 _03087_ net407 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__mux2_1
X_09696_ _04476_ _03705_ _03780_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__and4b_1
XFILLER_0_68_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08647_ datapath.PC\[8\] _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout827_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ net688 _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07529_ datapath.rf.registers\[0\]\[17\] net827 _02448_ _02455_ vssd1 vssd1 vccd1
+ vccd1 _02456_ sky130_fd_sc_hd__o22a_4
XANTENNA__08266__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10540_ net1048 _05419_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__nor2_1
XANTENNA__07474__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10471_ net1784 _01434_ _05256_ datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 _00002_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08018__A2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10953__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12210_ net273 net1958 net574 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
XANTENNA__07226__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ clknet_leaf_108_clk _00182_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08974__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ _06397_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__and2_1
X_12072_ _06335_ _06340_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a21o_1
Xhold590 datapath.rf.registers\[7\]\[18\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08726__A0 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net163 net2317 net584 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ net264 net2065 net606 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__mux2_1
X_11925_ net152 _05877_ net127 net2617 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_142_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _06247_ datapath.PC\[27\] net305 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10807_ net2129 net259 net602 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14575_ net1345 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11787_ net700 _04800_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08257__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10738_ datapath.PC\[1\] net839 vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__or2_1
X_13526_ clknet_leaf_73_clk _00476_ net1245 vssd1 vssd1 vccd1 vccd1 datapath.PC\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07465__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11261__B2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11959__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ clknet_leaf_81_clk _00413_ net1242 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08009__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ _05520_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12408_ net1651 net285 net464 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XANTENNA__07217__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06642__A mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_92_clk net1368 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
X_12339_ net2528 net299 net475 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08717__A0 _03146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ net1001 net986 net979 _01801_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__and4_1
X_14009_ clknet_leaf_48_clk _00896_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06991__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ datapath.rf.registers\[23\]\[9\] net933 net878 datapath.rf.registers\[29\]\[9\]
+ _02806_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a221o_1
XANTENNA__08193__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13756__RESET_B net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ _01638_ net991 _01656_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__and3_1
X_09550_ net676 _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__and2_1
X_06762_ _01417_ net1005 _01680_ _01685_ _01688_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__a311o_1
X_08501_ _03363_ _03365_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09481_ net332 _04405_ _04406_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o31a_1
XFILLER_0_144_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06693_ _01593_ _01600_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_65_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08432_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ datapath.rf.registers\[31\]\[0\] net948 net923 datapath.rf.registers\[2\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout143_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07314_ datapath.rf.registers\[19\]\[22\] net946 net695 _02240_ vssd1 vssd1 vccd1
+ vccd1 _02241_ sky130_fd_sc_hd__a211o_1
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07456__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__B2 _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ datapath.rf.registers\[8\]\[1\] net996 _01731_ _01742_ vssd1 vssd1 vccd1
+ vccd1 _03221_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07245_ _02170_ _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout310_A _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1052_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07208__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ net832 _02088_ _02090_ _02102_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1160_A datapath.rf.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout300 _05586_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
Xfanout311 _05859_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_2
Xfanout1309 net1311 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__clkbuf_4
Xfanout322 net324 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
Xfanout333 net334 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06698__S net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net358 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_1
Xfanout366 _03540_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_1
X_09817_ _04741_ _04743_ _04729_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a21o_1
Xfanout377 net379 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_2
Xfanout388 _03522_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout944_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XANTENNA__08198__B _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ datapath.PC\[20\] net629 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__nor2_1
XANTENNA__10279__C1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _04597_ _04600_ _04603_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a31o_1
XANTENNA__10948__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ net1300 screen.counter.ct\[0\] net1298 screen.counter.ct\[3\] vssd1 vssd1
+ vccd1 vccd1 _06147_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_124_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10294__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07695__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ net2465 net213 net433 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
X_11641_ net2621 _06100_ _06102_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08239__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07447__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ clknet_leaf_42_clk _01247_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11572_ screen.controlBus\[7\] _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nand2_1
XANTENNA__11243__B2 _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13311_ clknet_leaf_111_clk _00301_ net1098 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_10523_ _05406_ net1026 vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__nor2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_14291_ clknet_leaf_49_clk _01178_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13242_ clknet_leaf_77_clk _00232_ net1247 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
X_10454_ _02234_ net342 net525 vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nand3_1
XANTENNA__09739__A2 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10203__C1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ clknet_leaf_30_clk _00165_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10385_ _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12124_ datapath.mulitply_result\[24\] datapath.multiplication_module.multiplicand_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06973__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _06326_ _06328_ _06325_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__a21boi_1
XANTENNA__11808__A _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__B _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12403__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ net251 net2329 net582 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11019__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10858__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ net195 net2546 net543 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ net1484 _05893_ net156 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
X_12888_ net215 net2228 net552 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ _05516_ net176 _06235_ net179 vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07438__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14558_ net1331 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__11785__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ clknet_leaf_74_clk _00459_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_153_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14489_ clknet_leaf_47_clk _01376_ net1197 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08571__B _03496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07030_ datapath.rf.registers\[3\]\[28\] net767 net727 datapath.rf.registers\[2\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08290__C _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10606__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07610__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08981_ _03900_ _03907_ _03905_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06964__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ datapath.rf.registers\[12\]\[8\] net736 net724 datapath.rf.registers\[27\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XANTENNA__12313__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ net515 _02786_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__and2_1
X_06814_ net998 _01682_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nor2_2
X_09602_ _04453_ _04528_ net418 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
X_07794_ datapath.rf.registers\[0\]\[11\] net827 _02713_ _02720_ vssd1 vssd1 vccd1
+ vccd1 _02721_ sky130_fd_sc_hd__o22a_4
X_09533_ net331 _04251_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nand2_1
X_06745_ _01453_ _01576_ _01580_ _01479_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout260_A _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _03640_ _03657_ net341 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__mux2_1
X_06676_ _01483_ net1029 net1008 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__and3_1
XANTENNA__08874__C1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07141__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ _02172_ _02214_ _03340_ _02169_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__o31a_1
XFILLER_0_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09395_ net511 net352 _04215_ net386 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1267_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ datapath.rf.registers\[1\]\[0\] net973 _01735_ vssd1 vssd1 vccd1 vccd1 _03273_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07429__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ datapath.rf.registers\[0\]\[1\] net693 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07228_ datapath.rf.registers\[16\]\[24\] net963 net898 datapath.rf.registers\[6\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07159_ datapath.rf.registers\[9\]\[25\] net780 net753 datapath.rf.registers\[22\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ _01428_ _04007_ net540 vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__mux2_1
XANTENNA__07601__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1106 net1108 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
Xfanout1117 net1119 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12223__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 _05865_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_4
Xfanout141 net148 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_2
Xfanout1139 net1143 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_4
Xfanout152 net155 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout163 net166 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout174 _05562_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_2
Xfanout185 _05555_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_126_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout196 _05537_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_2
X_13860_ clknet_leaf_14_clk _00747_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08937__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ net259 net1847 net557 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09657__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ clknet_leaf_38_clk _00678_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11363__A _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10267__A2 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12742_ net269 net1945 net567 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__mux2_1
XANTENNA__08865__C1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12893__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12673_ net2436 net282 net431 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
X_11624_ screen.counter.ct\[21\] screen.counter.ct\[22\] _06086_ vssd1 vssd1 vccd1
+ vccd1 _06087_ sky130_fd_sc_hd__nand3_1
X_14412_ clknet_leaf_31_clk _01299_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ screen.register.currentYbus\[7\] _05772_ _06020_ vssd1 vssd1 vccd1 vccd1
+ _06021_ sky130_fd_sc_hd__a21o_1
X_14343_ clknet_leaf_19_clk _01230_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09290__C1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10506_ net38 _05345_ _05411_ net37 vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07840__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ clknet_leaf_43_clk _01161_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ screen.register.currentXbus\[27\] net1013 _05737_ screen.register.currentYbus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a22o_1
X_13225_ clknet_leaf_88_clk _00216_ net1211 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ screen.register.currentXbus\[25\] screen.register.currentXbus\[24\] screen.register.currentXbus\[27\]
+ screen.register.currentXbus\[26\] vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__or4_1
XANTENNA__09042__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09593__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ clknet_leaf_17_clk _00148_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ _05287_ _05289_ _05274_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06946__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13348__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ datapath.mulitply_result\[21\] datapath.multiplication_module.multiplicand_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nor2_1
X_13087_ clknet_leaf_39_clk _00079_ net1152 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10299_ net365 _04239_ _05224_ _05225_ net373 vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__o221a_1
X_12038_ datapath.mulitply_result\[10\] datapath.multiplication_module.multiplicand_i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__or2_1
XANTENNA__11972__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07371__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13989_ clknet_leaf_108_clk _00876_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08566__B _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06530_ mmio.memload_or_instruction\[28\] net1059 vssd1 vssd1 vccd1 vccd1 _01460_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08320__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07123__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08285__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08200_ _03124_ _03125_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09180_ net419 _03874_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ datapath.rf.registers\[29\]\[4\] net717 _03057_ net831 vssd1 vssd1 vccd1
+ vccd1 _03058_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08084__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12308__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06814__B _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08062_ datapath.rf.registers\[16\]\[5\] net961 net852 datapath.rf.registers\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07831__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07013_ datapath.rf.registers\[30\]\[29\] net910 net902 datapath.rf.registers\[20\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09033__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ _03629_ _03757_ net394 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__mux2_1
X_07915_ datapath.rf.registers\[29\]\[8\] net877 net857 datapath.rf.registers\[15\]\[8\]
+ _02837_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__a221o_1
X_08895_ net339 _03813_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__nor3_1
XANTENNA__12978__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ datapath.rf.registers\[5\]\[10\] net782 net722 datapath.rf.registers\[27\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a22o_1
XANTENNA__07898__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07362__A2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ datapath.rf.registers\[18\]\[11\] net789 net770 datapath.rf.registers\[30\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06728_ datapath.ru.latched_instruction\[23\] _01503_ net1027 vssd1 vssd1 vccd1 vccd1
+ _01655_ sky130_fd_sc_hd__mux2_1
X_09516_ net615 _04436_ _04442_ net676 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_104_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07114__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09447_ _02880_ _03494_ net680 _02885_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__a221o_1
X_06659_ _01501_ net1009 net1042 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06873__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ net639 _04291_ _04304_ _04282_ net653 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__a2111o_1
X_08329_ datapath.rf.registers\[23\]\[0\] net988 _01739_ vssd1 vssd1 vccd1 vccd1 _03256_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08075__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ mmio.memload_or_instruction\[19\] net1058 net307 net311 datapath.ru.latched_instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__a32o_1
XANTENNA__07822__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10961__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ net1308 mmio.wishbone.prev_BUSY_O net1045 vssd1 vssd1 vccd1 vccd1 _05847_
+ sky130_fd_sc_hd__and3b_1
X_13010_ net1466 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
X_10222_ net700 _04116_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__and2_1
X_10153_ _05058_ _05069_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_7_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ datapath.PC\[17\] _03579_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__nand2_1
XANTENNA__12888__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 keypad.debounce.debounce\[8\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
X_13912_ clknet_leaf_42_clk _00799_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ clknet_leaf_61_clk _00730_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13774_ clknet_leaf_116_clk _00661_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10986_ net188 net2562 net588 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__mux2_1
XANTENNA__07105__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12725_ net198 net2265 net572 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08606__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ net217 net2106 net438 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11607_ screen.counter.ct\[9\] net1293 _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__and3_1
XANTENNA__08066__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09263__C1 _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ net1712 net226 net445 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06634__B mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07813__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06616__B2 datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14326_ clknet_leaf_24_clk _01213_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11538_ net1413 _06005_ _05901_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11967__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold408 datapath.rf.registers\[5\]\[9\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold419 datapath.mulitply_result\[13\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ screen.register.currentXbus\[26\] _05700_ _05777_ screen.register.currentYbus\[26\]
+ _05780_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a221o_1
XANTENNA__10871__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14257_ clknet_leaf_27_clk _01144_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ clknet_leaf_39_clk _00200_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14188_ clknet_leaf_31_clk _01075_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ clknet_leaf_61_clk _00131_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1108 datapath.rf.registers\[9\]\[26\] vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 datapath.rf.registers\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07700_ datapath.rf.registers\[6\]\[13\] net813 net805 datapath.rf.registers\[15\]\[13\]
+ _02626_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a221o_1
X_08680_ _03603_ _03606_ net421 vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__mux2_1
XANTENNA__08577__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07344__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ datapath.rf.registers\[4\]\[15\] net930 net893 datapath.rf.registers\[14\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XANTENNA__06809__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ datapath.rf.registers\[2\]\[16\] net728 net724 datapath.rf.registers\[27\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a22o_1
X_09301_ net641 _04226_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__nor2_1
X_06513_ columns.count\[7\] columns.count\[6\] columns.count\[8\] vssd1 vssd1 vccd1
+ vccd1 _01445_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07493_ datapath.rf.registers\[4\]\[18\] net930 net914 datapath.rf.registers\[18\]\[18\]
+ _02419_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ net389 _03816_ _04158_ net391 vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06825__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08057__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ net367 _04066_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ net650 _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__or2_1
XANTENNA__07804__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09094_ net398 _03812_ _03516_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08045_ _01613_ _01727_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold920 datapath.rf.registers\[7\]\[12\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 datapath.rf.registers\[27\]\[27\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold942 datapath.rf.registers\[14\]\[21\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 datapath.rf.registers\[23\]\[1\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 datapath.rf.registers\[13\]\[1\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 datapath.rf.registers\[9\]\[17\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11364__B1 _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout592_A _05673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 datapath.rf.registers\[26\]\[17\] vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold997 datapath.rf.registers\[28\]\[26\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07375__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _04921_ _04922_ _04497_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_4_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07583__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _03602_ _03604_ net413 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout857_A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _03803_ _03804_ net363 vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a21o_1
XANTENNA__07335__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08532__A1 _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ datapath.rf.registers\[3\]\[10\] net964 net900 datapath.rf.registers\[20\]\[10\]
+ _02752_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a221o_1
X_10840_ net1808 net244 net603 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ net839 _04359_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__nand2_1
XANTENNA__10956__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12510_ net2539 net274 net453 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__mux2_1
X_13490_ clknet_leaf_80_clk _00443_ net1239 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12441_ net284 net2210 net463 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10257__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12372_ net299 net1951 net468 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11323_ datapath.ru.latched_instruction\[2\] net313 net309 _01478_ vssd1 vssd1 vccd1
+ vccd1 _00325_ sky130_fd_sc_hd__a22o_1
X_14111_ clknet_leaf_38_clk _00998_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ net1441 net142 net135 _02368_ vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__a22o_1
X_14042_ clknet_leaf_22_clk _00929_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10205_ _04801_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or2_1
X_11185_ mmio.key_data\[2\] net220 _05829_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ _04192_ _04337_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__and2_1
XANTENNA__11816__A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12411__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ net1052 _04991_ _04993_ net704 vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_50_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08523__A1 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13826_ clknet_leaf_43_clk _00713_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13757_ clknet_leaf_23_clk _00644_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10866__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10969_ net267 net2176 net586 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ net273 net1898 net570 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[5\] net1228
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11264__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ net285 net2382 net436 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ clknet_leaf_107_clk _01196_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold205 datapath.rf.registers\[10\]\[7\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 datapath.rf.registers\[5\]\[7\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 datapath.rf.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 datapath.rf.registers\[11\]\[1\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 datapath.rf.registers\[25\]\[11\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08211__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlymetal6s2s_1
X_09850_ _04775_ _04668_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__and2b_1
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_4
Xfanout729 _01779_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07565__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__A1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09691__A _03288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ _02079_ net352 _03725_ net388 vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__a211o_1
X_09781_ _04706_ _04707_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__nor2_1
X_06993_ datapath.rf.registers\[2\]\[29\] net728 net721 datapath.rf.registers\[28\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XANTENNA__12321__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08732_ _03655_ _03658_ net413 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__mux2_1
XANTENNA__08514__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ datapath.PC\[28\] _03589_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07614_ datapath.rf.registers\[18\]\[15\] net790 _02536_ _02538_ _02540_ vssd1 vssd1
+ vccd1 vccd1 _02541_ sky130_fd_sc_hd__a2111o_1
X_08594_ _01646_ _03507_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_101_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ _02465_ _02467_ _02469_ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout438_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ datapath.rf.registers\[24\]\[18\] net756 _02397_ _02402_ vssd1 vssd1 vccd1
+ vccd1 _02403_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_81_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06555__A mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09215_ net498 net495 net515 vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09146_ net638 _04072_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ net642 _04003_ _04002_ net625 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_116_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ datapath.rf.registers\[25\]\[6\] net796 net770 datapath.rf.registers\[30\]\[6\]
+ _02953_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a221o_1
Xhold750 datapath.rf.registers\[19\]\[30\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold761 datapath.rf.registers\[22\]\[6\] vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold772 datapath.rf.registers\[22\]\[20\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 screen.register.currentXbus\[5\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08202__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11888__A1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 datapath.rf.registers\[28\]\[4\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07556__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__B1 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__B1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _04837_ _04840_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__or2_1
XANTENNA__12231__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ net2410 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07308__A2 _02234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ net152 _05893_ net127 screen.register.currentXbus\[27\] vssd1 vssd1 vccd1
+ vccd1 _00538_ sky130_fd_sc_hd__a22o_1
XANTENNA__10312__A1 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11872_ _06259_ datapath.PC\[31\] net305 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__mux2_1
X_13611_ clknet_leaf_2_clk _00549_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08269__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ _03977_ _05651_ net846 vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_118_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08808__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11371__A _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ clknet_leaf_87_clk _00492_ net1219 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ _04309_ _05592_ net844 vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ clknet_leaf_84_clk _00426_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10685_ datapath.mulitply_result\[25\] net429 net661 vssd1 vssd1 vccd1 vccd1 _05536_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12424_ net2282 net224 net465 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12406__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ net2184 net243 net473 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__mux2_1
XANTENNA__11310__S _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__A2 _02721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _01446_ _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__nand2_2
X_12286_ net1746 net237 net480 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14025_ clknet_leaf_2_clk _00912_ net1075 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11237_ net1488 net141 net136 _03176_ vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07547__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__B1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ net1051 _05043_ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10450__A _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ net1287 net1288 vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07180__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ clknet_leaf_8_clk _00696_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_109_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ _02236_ net527 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08293__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07261_ datapath.rf.registers\[4\]\[23\] net810 net741 datapath.rf.registers\[1\]\[23\]
+ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09000_ net334 _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10328__C _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ _02112_ _02114_ _02116_ _02118_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__or4_1
XANTENNA__08590__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12316__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06822__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06994__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09902_ _04826_ _04828_ _04783_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 _03178_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_4
Xfanout515 _02763_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_4
XANTENNA__07538__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout526 _02301_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_4
Xfanout537 net540 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
X_09833_ _04700_ _04702_ _04758_ _04698_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a31o_1
Xfanout548 _06470_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_4
XANTENNA_fanout290_A _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_8
X_09764_ net632 _04690_ datapath.PC\[16\] vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__o21a_1
X_06976_ _01898_ _01900_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__or3_1
X_08715_ _03640_ _03641_ net408 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__mux2_1
X_09695_ _03786_ _03833_ _04450_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08646_ _01426_ _03572_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07710__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout722_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ net1003 _03443_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__or2_4
XFILLER_0_64_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ net831 _02452_ _02453_ _02454_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__or4_1
X_07459_ datapath.rf.registers\[9\]\[19\] net886 net853 datapath.rf.registers\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10470_ _05384_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.zero_multi
+ sky130_fd_sc_hd__inv_2
XFILLER_0_150_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09129_ net398 _03854_ _03516_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_131_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12226__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08974__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ net323 _06400_ _06401_ net327 net1973 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a32o_1
XANTENNA__06985__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ _06342_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__or2_1
Xhold580 datapath.rf.registers\[7\]\[17\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07529__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 datapath.rf.registers\[29\]\[19\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ net169 net2635 net584 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
XANTENNA__08726__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06737__B1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ net267 net2622 net606 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__mux2_1
XANTENNA__12896__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1280 datapath.ru.latched_instruction\[25\] vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11924_ net151 _05876_ net126 screen.register.currentXbus\[10\] vssd1 vssd1 vccd1
+ vccd1 _00521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07162__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11855_ net836 _04561_ _04664_ _05545_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _01509_ net709 _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__o22a_2
XFILLER_0_83_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14574_ net1344 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
X_11786_ net700 _04383_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ clknet_leaf_63_clk _00475_ net1271 vssd1 vssd1 vccd1 vccd1 datapath.PC\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_153_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11261__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ net839 _05208_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13456_ clknet_leaf_77_clk _00412_ net1238 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10668_ datapath.PC\[23\] _05514_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__nor2_1
XANTENNA__08614__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12407_ net1638 net295 net465 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13387_ clknet_leaf_92_clk net1376 net1201 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10599_ net1587 net516 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[11\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06642__B mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__07768__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
X_12338_ net1569 net288 net472 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_81_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11975__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12269_ net1625 net182 net481 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__mux2_1
XANTENNA__08717__A1 _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ clknet_leaf_42_clk _00895_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08193__A2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ net993 _01756_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__and2_2
XANTENNA__07940__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ _01411_ _01649_ _01687_ net1004 _01686_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a221o_1
X_08500_ _02170_ _03426_ _02171_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a21bo_1
X_06692_ _01606_ _01619_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__nand2_1
X_09480_ net331 net376 _04247_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_19_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08431_ _01931_ net534 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06817__B _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ datapath.rf.registers\[24\]\[0\] net907 net899 datapath.rf.registers\[6\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a22o_1
X_07313_ datapath.rf.registers\[8\]\[22\] net927 net871 datapath.rf.registers\[27\]\[22\]
+ _02239_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11252__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ datapath.rf.registers\[16\]\[1\] _01731_ net972 vssd1 vssd1 vccd1 vccd1 _03220_
+ sky130_fd_sc_hd__and3_1
X_07244_ _02148_ _02167_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07175_ datapath.rf.registers\[20\]\[25\] net803 _02099_ _02101_ vssd1 vssd1 vccd1
+ vccd1 _02102_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout303_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06967__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1212_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 _05859_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_2
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout334 _03533_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout672_A _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08184__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_2
X_09816_ _04729_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nor2_1
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_2
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_2
XANTENNA__07392__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ net629 _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_129_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06959_ datapath.rf.registers\[10\]\[30\] net917 net906 datapath.rf.registers\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout937_A _01817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ net615 _04597_ _04604_ net676 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_38_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ net655 net616 vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_124_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ screen.counter.currentCt\[1\] _06100_ net664 vssd1 vssd1 vccd1 vccd1 _06102_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_64_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11571_ _05728_ _05806_ _05810_ _05725_ _05730_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__o221a_1
XANTENNA__10964__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13310_ clknet_leaf_112_clk _00300_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_10522_ _05410_ _05422_ net1025 vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_138_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14290_ clknet_leaf_34_clk _01177_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ _02059_ _02191_ _05361_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or3_1
X_13241_ clknet_leaf_77_clk _00231_ net1247 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10384_ _05304_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__nand2_1
X_13172_ clknet_leaf_114_clk _00164_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ datapath.mulitply_result\[24\] datapath.multiplication_module.multiplicand_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nand2_1
X_12054_ net2476 net325 net321 _06329_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a22o_1
XANTENNA__09372__A1 _02742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ net256 net1940 net582 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07383__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_4
X_12956_ net198 net2187 net542 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__mux2_1
XANTENNA__07135__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ net1482 _05892_ net156 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
X_12887_ net219 net2107 net552 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11838_ net837 _04782_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__nand2_1
XANTENNA__09427__A2 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10874__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14557_ net1330 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_60_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11769_ datapath.PC\[3\] net302 _06180_ _06184_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ clknet_leaf_75_clk _00458_ net1251 vssd1 vssd1 vccd1 vccd1 datapath.PC\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07989__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14488_ clknet_leaf_39_clk _01375_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13439_ clknet_leaf_85_clk _00395_ net1231 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12195__B1 _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06949__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08980_ net708 _03906_ net624 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_58_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07931_ datapath.rf.registers\[7\]\[8\] net824 net817 datapath.rf.registers\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a22o_1
X_07862_ net515 _02786_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__or2_1
XANTENNA__07913__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _04479_ _04527_ net411 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_1
X_06813_ net996 _01739_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__and2_4
X_07793_ _02715_ _02716_ _02717_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__or4_1
XANTENNA__09115__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09115__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _04455_ _04457_ _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nand3_1
X_06744_ datapath.ru.n_memwrite2 datapath.ru.n_memread2 vssd1 vssd1 vccd1 vccd1 _01671_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07126__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09463_ net641 _04387_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__nand2_1
X_06675_ net709 vssd1 vssd1 vccd1 vccd1 datapath.MemRead sky130_fd_sc_hd__inv_2
XFILLER_0_148_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08414_ _02214_ _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__nor2_1
X_09394_ net329 _03772_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08345_ datapath.rf.registers\[29\]\[0\] net988 _01756_ vssd1 vssd1 vccd1 vccd1 _03272_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1162_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A _02654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ net691 _03184_ net645 net644 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_78_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07227_ datapath.rf.registers\[13\]\[24\] net866 net850 datapath.rf.registers\[1\]\[24\]
+ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08929__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ _02083_ _02084_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout887_A _01841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ datapath.rf.registers\[0\]\[27\] net829 _02015_ vssd1 vssd1 vccd1 vccd1 _02016_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_100_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_4
Xfanout131 _05865_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_2
Xfanout1129 net1130 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
Xfanout142 net148 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout164 net166 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07365__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout186 _05555_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_2
Xfanout197 _05537_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_1
XANTENNA__10959__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12810_ net261 net2192 net557 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07117__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13790_ clknet_leaf_50_clk _00677_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__D1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11363__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ net274 net1988 net566 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10672__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12672_ net1613 net285 net431 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14411_ clknet_leaf_101_clk _01298_ net1226 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_146_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11623_ net1281 net1283 net1280 _06085_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__and4_1
XANTENNA__06891__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14342_ clknet_leaf_114_clk _01229_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11554_ screen.register.currentYbus\[23\] _05775_ _05777_ screen.register.currentYbus\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10505_ _05345_ net37 net38 _05411_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_137_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14273_ clknet_leaf_40_clk _01160_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11485_ screen.register.currentXbus\[3\] _05720_ _05735_ screen.register.currentYbus\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ clknet_leaf_91_clk _00215_ net1211 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10436_ screen.register.currentXbus\[29\] screen.register.currentXbus\[28\] screen.register.currentXbus\[31\]
+ screen.register.currentXbus\[30\] vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__or4_1
XANTENNA__10727__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ clknet_leaf_104_clk _00147_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12414__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ _01441_ _05279_ _05284_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or4_1
X_12106_ datapath.mulitply_result\[21\] datapath.multiplication_module.multiplicand_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_155_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13086_ clknet_leaf_52_clk _00078_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10298_ _03307_ net360 net361 vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a21o_1
XANTENNA__08148__A2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
X_12037_ datapath.mulitply_result\[10\] datapath.multiplication_module.multiplicand_i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nand2_1
XANTENNA__07356__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10869__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13988_ clknet_leaf_16_clk _00875_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07108__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ net273 net2156 net544 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08320__A2 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08608__A0 _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11207__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ datapath.rf.registers\[15\]\[4\] net805 net782 datapath.rf.registers\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08061_ datapath.rf.registers\[22\]\[5\] net952 net895 datapath.rf.registers\[14\]\[5\]
+ _02987_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__a221o_1
X_07012_ datapath.rf.registers\[21\]\[29\] net939 net879 datapath.rf.registers\[29\]\[29\]
+ _01938_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12324__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06830__B _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08963_ net638 _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07914_ datapath.rf.registers\[17\]\[8\] net882 net871 datapath.rf.registers\[27\]\[8\]
+ _02840_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a221o_1
XANTENNA__07347__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ net395 _03691_ _03819_ net402 vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__o211a_1
X_07845_ datapath.rf.registers\[13\]\[10\] net795 net766 datapath.rf.registers\[3\]\[10\]
+ _02771_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout468_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ datapath.rf.registers\[23\]\[11\] net786 net730 datapath.rf.registers\[16\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a22o_1
XANTENNA__06558__A mmio.memload_or_instruction\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09515_ net635 _04429_ _04437_ net610 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a22o_1
X_06727_ datapath.ru.latched_instruction\[15\] net1037 net1004 _01652_ vssd1 vssd1
+ vccd1 vccd1 _01654_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08311__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09446_ net513 _02879_ net684 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o21a_1
X_06658_ _01586_ _01587_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout802_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06873__A2 _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ net340 _04295_ _04301_ _04302_ net640 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o311a_1
XFILLER_0_148_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06589_ net1306 net1302 mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ _01519_ sky130_fd_sc_hd__or3b_1
X_08328_ datapath.rf.registers\[11\]\[0\] net994 _01763_ vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09272__B1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08259_ datapath.rf.registers\[11\]\[1\] net969 net899 datapath.rf.registers\[6\]\[1\]
+ _03185_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12159__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ mmio.wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11906__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _05146_ _05147_ net1056 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__mux2_1
XANTENNA__07586__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _05075_ _05078_ datapath.PC\[5\] net1243 vssd1 vssd1 vccd1 vccd1 _05079_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07050__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ datapath.PC\[17\] net1311 vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__nand2_1
XANTENNA__07338__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 mmio.key_en1 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ clknet_leaf_44_clk _00798_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_35_clk _00729_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11093__B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ clknet_leaf_119_clk _00660_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10985_ net194 net2464 net587 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__B1 _05500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ net209 net2135 net571 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06864__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12655_ net222 net2308 net437 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XANTENNA__12409__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11606_ screen.counter.ct\[7\] net1294 _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12586_ net1880 net243 net445 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
XANTENNA__06634__C mmio.memload_or_instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14325_ clknet_leaf_28_clk _01212_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11537_ _05930_ _05995_ _05996_ _06004_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__or4_1
XFILLER_0_151_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 datapath.rf.registers\[27\]\[8\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ clknet_leaf_4_clk _01143_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11468_ net1535 _05902_ _05939_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__a21o_1
XANTENNA__06931__A _01849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ clknet_leaf_45_clk _00199_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08369__A2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ net347 _05338_ vssd1 vssd1 vccd1 vccd1 datapath.ack_mul sky130_fd_sc_hd__nor2_1
XANTENNA__10453__A _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14187_ clknet_leaf_17_clk _01074_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11399_ _02368_ net668 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__and2_1
XANTENNA__07577__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07041__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ clknet_leaf_36_clk _00130_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13069_ clknet_leaf_0_clk _00061_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
Xhold1109 datapath.rf.registers\[2\]\[23\] vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07630_ datapath.rf.registers\[15\]\[15\] net858 net849 datapath.rf.registers\[1\]\[15\]
+ _02556_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a221o_1
X_07561_ datapath.rf.registers\[8\]\[16\] net739 net716 datapath.rf.registers\[29\]\[16\]
+ _02487_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a221o_1
X_09300_ net491 _04226_ net674 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06512_ keypad.alpha vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07492_ datapath.rf.registers\[13\]\[18\] net865 net849 datapath.rf.registers\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ _02389_ net356 _03929_ net385 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__a211o_1
XANTENNA__12319__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06825__B _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09162_ _04087_ _04088_ net364 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ net847 _01665_ _01726_ net992 vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ net402 _04018_ net339 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout216_A _05526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net831 _02968_ _02970_ _02952_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__o31a_4
XFILLER_0_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07280__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 datapath.rf.registers\[19\]\[24\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold921 datapath.rf.registers\[24\]\[29\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 datapath.rf.registers\[20\]\[20\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 datapath.rf.registers\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold954 datapath.rf.registers\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1125_A _00004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 datapath.rf.registers\[10\]\[19\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 datapath.rf.registers\[17\]\[19\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 datapath.rf.registers\[19\]\[22\] vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold998 datapath.rf.registers\[17\]\[10\] vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ net704 _04496_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout585_A _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08946_ _02478_ _02479_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_4_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ net497 net494 net524 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout752_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07828_ _02747_ _02748_ _02753_ _02754_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__or4_1
XANTENNA__07740__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ datapath.rf.registers\[2\]\[12\] net920 net876 datapath.rf.registers\[29\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07099__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ net1714 net282 net602 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09429_ net613 _04352_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or2_1
XANTENNA__12229__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ net294 net1801 net461 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10972__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net289 net2643 net471 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14110_ clknet_leaf_50_clk _00997_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11322_ datapath.ru.latched_instruction\[1\] net313 net309 _01464_ vssd1 vssd1 vccd1
+ vccd1 _00324_ sky130_fd_sc_hd__a22o_1
XANTENNA__07271__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ clknet_leaf_60_clk _00928_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11253_ net2134 net142 net135 _02410_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__a22o_1
XANTENNA__07559__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10204_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__and2_1
XANTENNA__06901__D net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ net1407 _05828_ _05831_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__a21o_1
XANTENNA__08220__B2 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12899__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ net1055 _05059_ _05061_ net835 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__o211a_1
X_10066_ _03582_ _04992_ net1054 vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_50_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11308__S _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06534__A1 mmio.memload_or_instruction\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13825_ clknet_leaf_42_clk _00712_ net1162 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13756_ clknet_leaf_58_clk _00643_ net1261 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10968_ net269 net2042 net587 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12707_ net279 net1620 net569 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__mux2_1
XANTENNA__09302__A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10448__A _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13687_ clknet_leaf_70_clk datapath.multiplication_module.multiplicand_i_n\[4\] net1228
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[4\] sky130_fd_sc_hd__dfrtp_1
X_10899_ net274 net1775 net597 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12638_ net295 net2505 net437 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11978__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12569_ net1546 net290 net444 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14308_ clknet_leaf_104_clk _01195_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold206 datapath.rf.registers\[23\]\[2\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 datapath.rf.registers\[4\]\[11\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 net80 vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold239 datapath.rf.registers\[10\]\[16\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ clknet_leaf_38_clk _01126_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11346__A1 _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07014__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout708 _01716_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_2
Xfanout719 _01782_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13332__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08800_ net529 net352 _03726_ net384 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__a211o_1
XANTENNA__09691__B _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ net1276 net632 _04705_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__nor3_1
XANTENNA__12602__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ _01913_ _01915_ _01916_ _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__or4_1
XANTENNA__07970__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ _03656_ _03657_ net408 vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__mux2_1
Xfanout1290 screen.counter.ct\[13\] vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10122__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ datapath.PC\[27\] _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__or2_1
XANTENNA__07722__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ datapath.rf.registers\[23\]\[15\] net787 net741 datapath.rf.registers\[1\]\[15\]
+ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ _03512_ net393 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout166_A _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07544_ datapath.rf.registers\[3\]\[17\] net967 net912 datapath.rf.registers\[18\]\[17\]
+ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06836__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10085__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ datapath.rf.registers\[5\]\[18\] net784 net738 datapath.rf.registers\[8\]\[18\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1075_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ net502 net618 net496 net516 vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09145_ net332 _04069_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__o31a_1
XANTENNA__10792__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07789__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09076_ _03324_ _03979_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07253__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08027_ datapath.rf.registers\[18\]\[6\] net789 net730 datapath.rf.registers\[16\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold740 datapath.rf.registers\[14\]\[22\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11337__A1 _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold751 datapath.rf.registers\[19\]\[28\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 datapath.rf.registers\[20\]\[10\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07005__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold773 datapath.rf.registers\[15\]\[29\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 datapath.rf.registers\[28\]\[13\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 datapath.rf.registers\[2\]\[30\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12512__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net836 _04904_ _04903_ net201 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o211a_1
XANTENNA__07961__B1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08929_ net524 net355 _03855_ net386 vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a211o_1
X_11940_ net151 _05892_ net126 screen.register.currentXbus\[26\] vssd1 vssd1 vccd1
+ vccd1 _00537_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07713__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14279__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _04610_ _06258_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__nand2_1
X_13610_ clknet_leaf_12_clk _00548_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10822_ datapath.PC\[15\] _05489_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13541_ clknet_leaf_97_clk _00491_ net1220 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11371__B _05695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10753_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__inv_2
XANTENNA__11812__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ clknet_leaf_84_clk _00425_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07492__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ _04518_ _05534_ net845 vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ net2398 net232 net466 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12354_ net1904 net234 net472 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06481__A datapath.ru.latched_instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11305_ columns.count\[1\] columns.count\[0\] columns.count\[3\] columns.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13293__CLK clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12285_ datapath.rf.registers\[3\]\[16\] net241 net482 vssd1 vssd1 vccd1 vccd1 _00730_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14024_ clknet_leaf_14_clk _00911_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11236_ net1446 net140 net134 _03244_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__a22o_1
X_11167_ _05323_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__nand2_1
XANTENNA__10731__A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ net1055 _03571_ _05044_ net698 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_147_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10450__B _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11098_ _01437_ net1294 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__nand2_1
X_10049_ _04964_ _04975_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10877__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13808_ clknet_leaf_0_clk _00695_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11264__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13739_ clknet_leaf_101_clk _00626_ net1226 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07260_ datapath.rf.registers\[3\]\[23\] net767 net746 datapath.rf.registers\[21\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09209__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10328__D _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07191_ datapath.rf.registers\[11\]\[25\] net971 net863 datapath.rf.registers\[28\]\[25\]
+ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10775__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ _04768_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout505 _03146_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_4
XFILLER_0_10_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout516 _02742_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
X_09832_ _04702_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nand2_1
Xfanout527 _02255_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12332__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout538 net540 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
Xfanout549 _06469_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07943__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _01662_ _04678_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__nor2_1
X_06975_ datapath.rf.registers\[11\]\[30\] net970 net942 datapath.rf.registers\[26\]\[30\]
+ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout283_A _05602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ net510 net509 net404 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__mux2_1
X_09694_ _04620_ _03906_ _03910_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__and3b_1
X_08645_ datapath.PC\[5\] datapath.PC\[6\] _03571_ vssd1 vssd1 vccd1 vccd1 _03572_
+ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout450_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1192_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ _03475_ _03501_ _03502_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07527_ datapath.rf.registers\[14\]\[17\] _01753_ net717 datapath.rf.registers\[29\]\[17\]
+ _02438_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a221o_1
XANTENNA__11255__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A _01783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07474__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07458_ _02379_ _02380_ _02382_ _02384_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_33_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12507__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07389_ datapath.rf.registers\[26\]\[20\] net822 net750 datapath.rf.registers\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a22o_1
XANTENNA__11558__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09128_ net680 _04048_ _04053_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__a211o_1
XANTENNA__07226__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ net329 net377 _03623_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__o31a_1
XFILLER_0_102_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10781__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12070_ datapath.mulitply_result\[15\] datapath.multiplication_module.multiplicand_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06572__C_N mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 datapath.rf.registers\[0\]\[7\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 datapath.rf.registers\[13\]\[6\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 datapath.rf.registers\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net173 net2541 net585 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07954__A_N net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ net269 net2487 net607 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__mux2_1
Xhold1270 screen.register.currentXbus\[23\] vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net151 _05875_ net126 screen.register.currentXbus\[9\] vssd1 vssd1 vccd1
+ vccd1 _00520_ sky130_fd_sc_hd__a22o_1
Xhold1281 datapath.mulitply_result\[7\] vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10697__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ net206 _04840_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11246__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ datapath.mulitply_result\[12\] net426 net658 vssd1 vssd1 vccd1 vccd1 _05637_
+ sky130_fd_sc_hd__a21o_1
X_14573_ net1343 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_11785_ datapath.PC\[7\] net302 _06194_ _06196_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09454__A3 _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ clknet_leaf_63_clk _00474_ net1272 vssd1 vssd1 vccd1 vccd1 datapath.PC\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_45_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ net1748 net182 net602 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13455_ clknet_leaf_81_clk _00411_ net1242 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12417__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ datapath.PC\[23\] _05514_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12406_ net1765 net291 net467 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07217__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ clknet_leaf_92_clk net1380 net1202 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10445__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ net2196 net515 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[10\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12337_ datapath.rf.registers\[5\]\[0\] net180 net472 vssd1 vssd1 vccd1 vccd1 _00778_
+ sky130_fd_sc_hd__mux2_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12268_ _06445_ _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nor2_4
X_14007_ clknet_leaf_44_clk _00894_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11219_ net1461 net145 net139 _04998_ vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__a22o_1
XANTENNA__10461__A _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__A1 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ _01602_ _01621_ net840 _01665_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__a31o_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__07925__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ _01406_ _01458_ net1028 _01493_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a31o_1
XANTENNA__09678__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07770__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06691_ _01608_ _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08350__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ _01620_ _01633_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11237__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ net651 _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a21o_2
XFILLER_0_129_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08102__B1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ datapath.rf.registers\[11\]\[22\] net971 net863 datapath.rf.registers\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
X_08292_ datapath.rf.registers\[19\]\[1\] net762 _03216_ _03217_ _03218_ vssd1 vssd1
+ vccd1 vccd1 _03219_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07456__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07243_ _02148_ net529 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12327__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06833__B _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout129_A _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07208__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07174_ datapath.rf.registers\[27\]\[25\] net724 net716 datapath.rf.registers\[29\]\[25\]
+ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a221o_1
XANTENNA__10748__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1038_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout498_A _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 _05859_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
XANTENNA__06719__A1 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 _06270_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1205_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 _03510_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
Xfanout346 _05333_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
XANTENNA__07916__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ datapath.PC\[4\] _03040_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nor2_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
Xfanout368 _03540_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
Xfanout379 _03536_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_1
X_09746_ datapath.PC\[20\] datapath.PC\[21\] datapath.PC\[22\] datapath.PC\[23\] vssd1
+ vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__or4_1
X_06958_ net648 net344 _01730_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_97_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07680__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09677_ net635 _04599_ _04601_ net611 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a22o_1
X_06889_ net999 net985 net979 _01801_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout832_A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ net655 net616 vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07695__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11228__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ net531 net529 net405 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__mux2_1
X_11570_ _06032_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07447__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10521_ _05401_ _05416_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12237__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13240_ clknet_leaf_76_clk _00230_ net1249 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ _02831_ _02876_ _03118_ _05360_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__or4b_1
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10739__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10980__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ clknet_leaf_53_clk _00163_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10383_ _05291_ screen.controlBus\[5\] screen.controlBus\[4\] _05296_ vssd1 vssd1
+ vccd1 vccd1 _05305_ sky130_fd_sc_hd__or4bb_1
X_12122_ net323 _06385_ _06386_ net327 net2220 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a32o_1
XANTENNA__07080__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__A _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ _06327_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__xnor2_1
X_11004_ net260 net1733 net582 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout880 net883 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_8
Xfanout891 _01839_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_4
XANTENNA__12700__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12955_ net209 net1715 net542 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ _05891_ _06263_ net149 net1438 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ net222 net1949 net551 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XANTENNA__06637__C mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11219__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ _06234_ datapath.PC\[21\] net304 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__mux2_1
XANTENNA__06894__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14556_ net1329 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__07438__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11768_ _06181_ net177 net175 _05170_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06934__A _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13507_ clknet_leaf_74_clk _00457_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10719_ _05563_ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14487_ clknet_leaf_45_clk _01374_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07843__C1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ screen.counter.currentCt\[20\] _06138_ screen.counter.currentCt\[21\] vssd1
+ vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13438_ clknet_leaf_90_clk _00394_ net1209 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13369_ clknet_leaf_70_clk _00354_ net1228 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07071__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07610__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07930_ datapath.rf.registers\[5\]\[8\] net783 net748 datapath.rf.registers\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__a22o_1
XANTENNA__08299__C _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__inv_2
X_09600_ _03664_ _04526_ _03456_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_1
X_06812_ _01639_ _01646_ _01656_ _01682_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__and4_4
XANTENNA__12610__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07792_ datapath.rf.registers\[29\]\[11\] net717 _02718_ net831 vssd1 vssd1 vccd1
+ vccd1 _02719_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _03449_ net419 net413 _04121_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__or4_1
X_06743_ _01604_ _01605_ datapath.ru.latched_instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ _01670_ sky130_fd_sc_hd__mux2_1
XANTENNA__06828__B _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__B1 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09462_ _03321_ _04388_ net641 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__a21o_1
X_06674_ _01594_ _01602_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__or2_1
XANTENNA__10130__B1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08413_ _02260_ _02304_ _03337_ _02256_ _02213_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o311a_1
X_09393_ net378 _03983_ _04319_ net332 vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ datapath.rf.registers\[10\]\[0\] net995 _01743_ vssd1 vssd1 vccd1 vccd1 _03271_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07429__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ net691 _03184_ _03195_ net644 vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__and4_1
XFILLER_0_116_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06563__B _01492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07226_ datapath.rf.registers\[30\]\[24\] net911 net890 datapath.rf.registers\[12\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11896__S net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14549__1360 vssd1 vssd1 vccd1 vccd1 net1360 _14549__1360/LO sky130_fd_sc_hd__conb_1
X_07157_ _02060_ _02079_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07088_ _01999_ _02000_ _02014_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__or3_1
XANTENNA__07601__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1111 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
Xfanout1119 net1124 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_2
Xfanout132 _05865_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
XFILLER_0_100_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout143 net144 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
XANTENNA__09354__A2 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 _05263_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08562__A0 _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_2
Xfanout176 _06183_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout187 _05555_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_1
XANTENNA__12520__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout198 _05537_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_2
X_09729_ _01908_ _03435_ _01864_ _01907_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ net278 net2207 net565 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__mux2_1
XANTENNA__07668__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12671_ net1927 net294 net431 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XANTENNA__10975__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12949__A0 _05496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14410_ clknet_leaf_15_clk _01297_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11622_ net1287 net1284 net1286 _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__and4_1
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ clknet_leaf_109_clk _01228_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11553_ screen.register.currentXbus\[7\] _05704_ _05707_ screen.register.currentXbus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ _05412_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14272_ clknet_leaf_45_clk _01159_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07840__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11484_ screen.register.currentXbus\[27\] _05700_ _05709_ screen.register.currentXbus\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13223_ clknet_leaf_91_clk _00214_ net1211 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10435_ screen.register.currentXbus\[17\] screen.register.currentXbus\[16\] screen.register.currentXbus\[19\]
+ screen.register.currentXbus\[18\] vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__or4_1
XFILLER_0_111_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09042__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13154_ clknet_leaf_43_clk _00146_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ screen.controlBus\[0\] _05285_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12105_ _06367_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__and2_1
X_13085_ clknet_leaf_23_clk _00077_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10297_ _03206_ net360 vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__nor2_1
X_12036_ net321 _06313_ _06314_ net325 net1838 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a32o_1
XANTENNA__08553__A0 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12430__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13987_ clknet_leaf_105_clk _00874_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12938_ net278 net2084 net541 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__mux2_1
XANTENNA__06867__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10885__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ net296 net1796 net550 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08608__A1 _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ net1326 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XANTENNA__08084__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08060_ datapath.rf.registers\[11\]\[5\] net968 net876 datapath.rf.registers\[29\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a22o_1
XANTENNA__07292__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07831__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07011_ datapath.rf.registers\[24\]\[29\] net906 net882 datapath.rf.registers\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a22o_1
XANTENNA__12605__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08962_ net330 _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__nand2_1
XANTENNA__06633__C_N mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07913_ datapath.rf.registers\[6\]\[8\] net898 _02839_ net695 vssd1 vssd1 vccd1 vccd1
+ _02840_ sky130_fd_sc_hd__a211o_1
X_08893_ net395 _03691_ _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o21a_1
XANTENNA__08544__A0 _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A _05537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ datapath.rf.registers\[7\]\[10\] net824 net737 datapath.rf.registers\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__a22o_1
XANTENNA__12340__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ _02700_ _02701_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__and2b_2
XANTENNA__06558__B _01455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ _01717_ _04440_ net625 vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__o21ai_1
X_06726_ datapath.ru.latched_instruction\[15\] net1037 net1004 _01652_ vssd1 vssd1
+ vccd1 vccd1 _01653_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_88_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09445_ net419 _03646_ _03649_ net319 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06858__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06657_ datapath.ru.latched_instruction\[1\] net1042 _01464_ net1009 vssd1 vssd1
+ vccd1 vccd1 _01587_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1272_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ net492 _04292_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__nand2_1
X_06588_ mmio.memload_or_instruction\[11\] net1062 vssd1 vssd1 vccd1 vccd1 _01518_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08327_ datapath.rf.registers\[25\]\[0\] net990 _01754_ vssd1 vssd1 vccd1 vccd1 _03254_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08075__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ datapath.rf.registers\[3\]\[1\] net967 net925 datapath.rf.registers\[8\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__a22o_1
XANTENNA__07822__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07209_ datapath.rf.registers\[11\]\[24\] net776 net757 datapath.rf.registers\[24\]\[24\]
+ _02135_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a221o_1
XANTENNA__12515__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ datapath.rf.registers\[21\]\[3\] net745 _03090_ _03091_ _03105_ vssd1 vssd1
+ vccd1 vccd1 _03116_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07035__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ net1277 _03574_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__xnor2_1
X_10151_ net203 _05077_ net1309 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ _05005_ _05008_ datapath.PC\[26\] net1271 vssd1 vssd1 vccd1 vccd1 _05009_
+ sky130_fd_sc_hd__o2bb2a_1
X_13910_ clknet_leaf_26_clk _00797_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12250__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ clknet_leaf_27_clk _00728_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11093__C _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ clknet_leaf_35_clk _00659_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ net196 net2143 net588 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__mux2_1
X_12723_ net215 net2090 net572 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ net233 net1963 net438 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _05715_ _05752_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12585_ net1754 net236 net444 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__mux2_1
XANTENNA__08066__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09263__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14324_ clknet_leaf_105_clk _01211_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06634__D mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ _05904_ _05994_ _06002_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__a211o_1
XANTENNA__07274__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07813__A2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14255_ clknet_leaf_5_clk _01142_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11467_ net975 _05812_ _05929_ _05938_ _05901_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__o221a_1
XANTENNA__12425__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06931__B _01852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07026__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ clknet_leaf_25_clk _00198_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10418_ _05334_ _05335_ _05336_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__or4_1
X_14186_ clknet_leaf_12_clk _01073_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11398_ screen.register.currentYbus\[18\] net130 _05884_ net159 vssd1 vssd1 vccd1
+ vccd1 _00376_ sky130_fd_sc_hd__a22o_1
XANTENNA__10453__B _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13467__D net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ clknet_leaf_8_clk _00129_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10349_ screen.counter.ct\[7\] net1294 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or2_1
X_13068_ clknet_leaf_29_clk _00060_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12019_ datapath.mulitply_result\[7\] datapath.multiplication_module.multiplicand_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ datapath.rf.registers\[23\]\[16\] net788 net747 datapath.rf.registers\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__a22o_1
XANTENNA__08829__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06511_ screen.screenEdge.enable3 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
X_07491_ datapath.rf.registers\[19\]\[18\] net945 net881 datapath.rf.registers\[17\]\[18\]
+ _02417_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a221o_1
X_09230_ net634 _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06825__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ net498 net495 net514 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a21o_1
XANTENNA__08057__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _03025_ _03028_ _03038_ net692 datapath.rf.registers\[0\]\[4\] vssd1 vssd1
+ vccd1 vccd1 _03039_ sky130_fd_sc_hd__o32a_2
XANTENNA__07265__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09092_ net402 _03820_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__nor2_1
XANTENNA__07804__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08043_ _02958_ _02962_ _02963_ _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold900 datapath.rf.registers\[13\]\[8\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12335__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold911 datapath.mulitply_result\[2\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 datapath.rf.registers\[30\]\[10\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07017__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09557__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 datapath.rf.registers\[8\]\[29\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 datapath.rf.registers\[31\]\[27\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 datapath.rf.registers\[14\]\[3\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 datapath.rf.registers\[29\]\[21\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 datapath.rf.registers\[0\]\[26\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold988 datapath.rf.registers\[15\]\[2\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net837 _04475_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__or2_1
Xhold999 datapath.rf.registers\[21\]\[29\] vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07953__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout480_A _06449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ net503 net619 _03543_ net526 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__a211o_1
X_07827_ datapath.rf.registers\[14\]\[10\] net892 net860 datapath.rf.registers\[28\]\[10\]
+ _02749_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a221o_1
XANTENNA__11194__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ datapath.rf.registers\[1\]\[12\] net848 _02680_ _02682_ _02684_ vssd1 vssd1
+ vccd1 vccd1 _02685_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08784__A _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06709_ _01636_ vssd1 vssd1 vccd1 vccd1 datapath.MUL_EN sky130_fd_sc_hd__inv_2
XFILLER_0_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout912_A _01830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ datapath.rf.registers\[26\]\[13\] net820 net744 datapath.rf.registers\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XANTENNA__08296__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ net653 _04342_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09359_ net365 _04133_ _04134_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12370_ net180 net2302 net471 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11321_ _01458_ net1029 net309 net313 datapath.ru.latched_instruction\[0\] vssd1
+ vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12245__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ clknet_leaf_37_clk _00927_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07008__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11252_ net1545 net140 net134 _02456_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _05124_ _05125_ _05129_ net200 vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__o211a_1
X_11183_ mmio.key_data\[1\] net220 _05829_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _03572_ _05060_ net1055 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07863__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ net1275 _03580_ datapath.PC\[19\] vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10315__B1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ clknet_leaf_47_clk _00711_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ net276 net2006 net588 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__mux2_1
X_13755_ clknet_leaf_54_clk _00642_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12706_ net280 net2481 net569 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__mux2_1
XANTENNA__07495__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11291__B2 mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08692__C1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10898_ net278 net1680 net594 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__mux2_1
X_13686_ clknet_leaf_70_clk datapath.multiplication_module.multiplicand_i_n\[3\] net1229
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10448__B _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12637_ net291 net2321 net436 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__mux2_1
XANTENNA__08039__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07247__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ net2070 net181 net447 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08995__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ clknet_leaf_105_clk _01194_ net1101 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11519_ _05814_ _05987_ _05986_ _05901_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10464__A _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ net167 net2250 net457 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__mux2_1
Xhold207 net65 vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 datapath.rf.registers\[18\]\[3\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 datapath.rf.registers\[4\]\[3\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ clknet_leaf_50_clk _01125_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14169_ clknet_leaf_60_clk _01056_ net1266 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08211__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net711 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
X_06991_ datapath.rf.registers\[15\]\[29\] net807 net780 datapath.rf.registers\[9\]\[29\]
+ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08730_ _02763_ net514 net404 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__mux2_1
Xfanout1280 screen.counter.ct\[20\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__clkbuf_2
Xfanout1291 screen.counter.ct\[12\] vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_2
X_08661_ datapath.PC\[26\] _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__or2_1
XANTENNA__07183__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ datapath.rf.registers\[7\]\[15\] net825 net749 datapath.rf.registers\[10\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a22o_1
X_08592_ net504 net622 _03517_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_85_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07543_ datapath.rf.registers\[31\]\[17\] net948 net856 datapath.rf.registers\[15\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06836__B _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout159_A _05261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__B2 mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ datapath.rf.registers\[10\]\[18\] net749 net735 datapath.rf.registers\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09213_ net361 _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07238__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ net330 net378 _03844_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or3b_1
XFILLER_0_115_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06852__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09075_ net642 _04000_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_116_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1235_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08026_ datapath.rf.registers\[5\]\[6\] net782 net765 datapath.rf.registers\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a22o_1
XANTENNA__11189__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold730 datapath.rf.registers\[27\]\[9\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 datapath.rf.registers\[21\]\[22\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__A0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout695_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 datapath.rf.registers\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 datapath.rf.registers\[25\]\[12\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08202__A2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold774 datapath.rf.registers\[15\]\[11\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 datapath.rf.registers\[20\]\[8\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 datapath.rf.registers\[6\]\[29\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net221 _04561_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout862_A _01851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06764__A2 _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__S net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net499 net620 net488 net523 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08859_ _02349_ _03420_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_28_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11870_ net201 _05571_ _06257_ net705 vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10821_ net1614 net252 net602 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__mux2_1
XANTENNA__09403__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08269__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13540_ clknet_leaf_88_clk _00490_ net1218 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10752_ _05482_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__or2_1
XANTENNA__07477__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13471_ clknet_leaf_84_clk _00424_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10983__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10683_ _05532_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nor2_1
XANTENNA__07229__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ net1917 net228 net465 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ net1695 net240 net474 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11304_ net26 net1045 net1034 net2575 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__o22a_1
X_12284_ net2618 net245 net482 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08729__A0 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14023_ clknet_leaf_15_clk _00910_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11235_ net1610 net142 net135 _03285_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12703__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07401__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _05716_ _05801_ _05814_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09941__A2 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net1278 datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _05044_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_147_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11097_ net1023 _05713_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nor2_1
X_10048_ net205 _04972_ _04974_ net1251 vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__o211a_1
Xhold90 screen.controlBus\[31\] vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07180__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ clknet_leaf_7_clk _00694_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10459__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _06282_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07468__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ clknet_leaf_10_clk _00625_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11264__B2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10893__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13669_ clknet_leaf_79_clk net1397 net1238 vssd1 vssd1 vccd1 vccd1 datapath.pc_module.i_ack1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07190_ datapath.rf.registers\[3\]\[25\] net966 net922 datapath.rf.registers\[2\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09983__A _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06994__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09900_ _04675_ _04767_ _04672_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12613__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout506 _03087_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _04708_ _04712_ _04755_ _04706_ _04703_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a311o_1
Xfanout517 _02698_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_4
Xfanout528 _02212_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09762_ _04688_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__inv_2
X_06974_ datapath.rf.registers\[16\]\[30\] net962 net930 datapath.rf.registers\[4\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
X_08713_ net513 net512 net404 vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__mux2_1
X_09693_ _03252_ _04615_ _04619_ _04617_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__or4b_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08644_ datapath.PC\[2\] datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1
+ _03571_ sky130_fd_sc_hd__or3_2
XANTENNA__07950__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06847__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ net319 _03492_ net686 _01863_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout1185_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ datapath.rf.registers\[24\]\[17\] net755 net737 datapath.rf.registers\[8\]\[17\]
+ _02439_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a221o_1
XANTENNA__07459__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ datapath.rf.registers\[7\]\[19\] net957 net917 datapath.rf.registers\[10\]\[19\]
+ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06582__A mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07388_ datapath.rf.registers\[25\]\[20\] net798 net791 datapath.rf.registers\[18\]\[20\]
+ _02314_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09127_ _02743_ net683 _03494_ _02744_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_98_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07631__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ net330 _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__nand2_1
X_08009_ datapath.rf.registers\[31\]\[6\] net948 net916 datapath.rf.registers\[10\]\[6\]
+ _02933_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__a221o_1
XANTENNA__06985__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 datapath.rf.registers\[11\]\[28\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
X_14527__1349 vssd1 vssd1 vccd1 vccd1 net1349 _14527__1349/LO sky130_fd_sc_hd__conb_1
Xhold571 datapath.rf.registers\[17\]\[16\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net186 net2529 net584 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
Xhold582 datapath.rf.registers\[16\]\[22\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 datapath.rf.registers\[16\]\[11\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06737__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ net274 net1675 net608 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__mux2_1
XANTENNA__10978__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1260 datapath.rf.registers\[16\]\[5\] vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 datapath.rf.registers\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ net152 _05874_ net127 screen.register.currentXbus\[8\] vssd1 vssd1 vccd1
+ vccd1 _00519_ sky130_fd_sc_hd__a22o_1
Xhold1282 net85 vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07162__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _06243_ _06244_ _06245_ net305 datapath.PC\[26\] vssd1 vssd1 vccd1 vccd1
+ _00470_ sky130_fd_sc_hd__a32o_1
X_10804_ _04047_ _05635_ net844 vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__mux2_1
X_14572_ net1342 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__11246__B2 _02721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11784_ _05610_ net175 _06195_ net177 vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__a22o_1
XANTENNA__11797__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13523_ clknet_leaf_63_clk _00473_ net1272 vssd1 vssd1 vccd1 vccd1 datapath.PC\[29\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_45_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10735_ _01458_ net711 _05577_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_45_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13454_ clknet_leaf_81_clk _00410_ net1238 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07870__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ net218 net2244 net608 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12405_ net2408 net297 net467 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
X_13385_ clknet_leaf_92_clk net1377 net1202 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597_ net1685 net514 net349 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[9\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10445__C net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
X_12336_ _05575_ _06445_ _06450_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__nor3_1
XANTENNA__07622__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12433__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ _05669_ _06443_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ net1437 net145 net138 _04976_ vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__a22o_1
X_14006_ clknet_leaf_26_clk _00893_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12198_ _01643_ _01666_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__nand2_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XANTENNA__10461__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
X_11149_ _05299_ net1014 _05767_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__or3_1
XANTENNA__09127__B1 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07689__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ _01611_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08360_ net651 _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a21oi_4
X_07311_ datapath.rf.registers\[31\]\[22\] net950 net939 datapath.rf.registers\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11788__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ datapath.rf.registers\[25\]\[1\] net990 _01754_ vssd1 vssd1 vccd1 vccd1 _03218_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_144_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12608__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06664__A1 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ _02148_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07173_ datapath.rf.registers\[26\]\[25\] net822 net747 datapath.rf.registers\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_113_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07613__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06967__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12343__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout303 net306 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_4
Xfanout314 _05859_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_2
Xfanout336 _03510_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
X_09814_ _04731_ _04740_ _04730_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a21o_1
Xfanout358 _03626_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout1100_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _03539_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_2
XANTENNA__07392__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ datapath.PC\[20\] net629 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and2_1
X_06957_ datapath.rf.registers\[0\]\[30\] net828 _01883_ vssd1 vssd1 vccd1 vccd1 _01884_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout658_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ net706 _04586_ net623 vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a21o_1
X_06888_ datapath.rf.registers\[31\]\[31\] net949 net945 datapath.rf.registers\[19\]\[31\]
+ _01811_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a221o_1
XANTENNA__07144__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08627_ _01634_ _03552_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout825_A _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08558_ net532 _02079_ net406 vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__mux2_1
X_07509_ _02411_ _02431_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08489_ _03376_ _03412_ _03377_ _02525_ _03374_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__o2111a_1
XANTENNA__12518__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10827__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10520_ _05396_ _05415_ net1025 vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06655__A1 _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07852__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ _02017_ _03176_ _03244_ _03285_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13475__RESET_B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ clknet_leaf_35_clk _00162_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07604__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ screen.controlBus\[3\] _05292_ _05301_ screen.controlBus\[2\] vssd1 vssd1
+ vccd1 vccd1 _05304_ sky130_fd_sc_hd__or4bb_1
XANTENNA__08575__A1_N net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ _06377_ _06381_ _06384_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__nand3_1
XANTENNA__06958__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12253__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _06320_ _06321_ _06322_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__o21bai_1
XANTENNA__11377__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 datapath.rf.registers\[30\]\[3\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net263 net1855 net582 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
XANTENNA__09109__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 _01848_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
XANTENNA__07383__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout881 net883 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_4
Xfanout892 net895 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11393__A _02499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ net215 net2306 net542 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
Xhold1090 datapath.rf.registers\[28\]\[8\] vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ _05890_ _06263_ net149 net1460 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ net232 datapath.rf.registers\[21\]\[20\] net552 vssd1 vssd1 vccd1 vccd1 _01310_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06637__D mmio.memload_or_instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ net201 _04828_ _05509_ _04664_ _04949_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__o221ai_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14555_ net1366 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__08096__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net204 net303 vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12428__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ clknet_leaf_76_clk _00456_ net1250 vssd1 vssd1 vccd1 vccd1 datapath.PC\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ datapath.PC\[30\] _05556_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ clknet_leaf_24_clk _01373_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11698_ net1508 _06138_ _06140_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13437_ clknet_leaf_89_clk _00393_ net1210 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10649_ _05503_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13368_ clknet_leaf_71_clk _00353_ net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06949__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net1672 net247 net478 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
X_13299_ clknet_leaf_110_clk _00289_ net1104 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08020__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _02764_ _02786_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__or2_1
XANTENNA__07374__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ net998 net977 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__nor2_2
X_07791_ datapath.rf.registers\[11\]\[11\] net774 net748 datapath.rf.registers\[10\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06742_ _01668_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__inv_2
X_09530_ _02433_ net685 net678 _02437_ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__A1 _03202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__B2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _02834_ _03320_ _02792_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a21o_1
X_06673_ _01584_ _01588_ _01598_ _01591_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_35_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10130__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08412_ _02260_ _02304_ _03337_ _02256_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__o31a_1
X_09392_ net371 _04317_ _04318_ net382 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ datapath.rf.registers\[4\]\[0\] net994 _01734_ vssd1 vssd1 vccd1 vccd1 _03270_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06562__C_N mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12338__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _03194_ _03196_ _03198_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__nor4_1
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07225_ datapath.rf.registers\[27\]\[24\] net871 net854 datapath.rf.registers\[5\]\[24\]
+ _02151_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__inv_2
X_07087_ _02002_ _02005_ _02006_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__or4_1
XFILLER_0_140_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1109 net1111 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout133 _05865_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12801__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout144 net148 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
XANTENNA__07365__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout166 _05574_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08562__A1 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 net178 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout942_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout199 _05537_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ datapath.rf.registers\[5\]\[7\] net782 net774 datapath.rf.registers\[11\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a22o_1
X_09728_ _02084_ _03362_ _03428_ _04631_ _03361_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a221o_1
XANTENNA__07117__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _01910_ _03437_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12670_ net1992 net291 net432 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XANTENNA__10672__A2 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11621_ screen.counter.ct\[13\] net1289 _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__and3_1
XANTENNA__08078__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12248__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ clknet_leaf_102_clk _01227_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07825__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ net1543 _05901_ _06018_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ net35 net36 _05346_ _05411_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__and4b_1
XFILLER_0_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11483_ net1511 _05953_ _05901_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14271_ clknet_leaf_38_clk _01158_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10434_ screen.register.currentXbus\[21\] screen.register.currentXbus\[20\] screen.register.currentXbus\[23\]
+ screen.register.currentXbus\[22\] vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or4_1
X_13222_ clknet_leaf_85_clk _00213_ net1231 vssd1 vssd1 vccd1 vccd1 screen.screenLogic.currentWrx
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_150_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09042__A2 _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ clknet_leaf_40_clk _00145_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10365_ screen.controlBus\[1\] _05279_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__or3_1
X_12104_ net324 _06370_ _06371_ net328 net1888 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__a32o_1
X_13084_ clknet_leaf_57_clk _00076_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10296_ _01625_ _03493_ _04658_ _05221_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o311a_1
X_12035_ _06311_ _06312_ _06310_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12711__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08553__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13986_ clknet_leaf_51_clk _00873_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07108__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06585__C_N mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ net280 net2022 net541 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__mux2_1
X_12868_ net292 datapath.rf.registers\[21\]\[3\] net550 vssd1 vssd1 vccd1 vccd1 _01293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ net701 _04819_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12799_ net180 net1978 net560 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14538_ net1325 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09018__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14469_ clknet_leaf_107_clk _01356_ net1110 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07010_ datapath.rf.registers\[7\]\[29\] net958 _01932_ _01934_ _01936_ vssd1 vssd1
+ vccd1 vccd1 _01937_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_113_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11915__A2 _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08241__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08961_ _03884_ _03887_ net381 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ datapath.rf.registers\[24\]\[8\] net907 net874 datapath.rf.registers\[25\]\[8\]
+ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a221o_1
XANTENNA__12621__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08892_ _03817_ _03818_ net391 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__a21o_1
XANTENNA__07347__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08544__A1 _03307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14185__RESET_B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ datapath.rf.registers\[10\]\[10\] net748 _02769_ net831 vssd1 vssd1 vccd1
+ vccd1 _02770_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06839__B _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _02679_ net517 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09513_ _02614_ _03411_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__xor2_1
X_06725_ datapath.ru.latched_instruction\[15\] _01461_ net1028 vssd1 vssd1 vccd1 vccd1
+ _01652_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11300__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1098_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06656_ datapath.ru.latched_instruction\[0\] net1042 net1009 _01585_ vssd1 vssd1
+ vccd1 vccd1 _01586_ sky130_fd_sc_hd__a22oi_2
X_09444_ _04368_ _04370_ net338 _03693_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06587_ datapath.ru.latched_instruction\[13\] _01516_ vssd1 vssd1 vccd1 vccd1 _01517_
+ sky130_fd_sc_hd__xnor2_1
X_09375_ net336 _03813_ _03821_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout523_A _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06574__B _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ datapath.rf.registers\[2\]\[0\] net973 _01741_ vssd1 vssd1 vccd1 vccd1 _03253_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07807__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08257_ datapath.rf.registers\[30\]\[1\] net909 net892 datapath.rf.registers\[14\]\[1\]
+ _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07208_ datapath.rf.registers\[5\]\[24\] net785 net716 datapath.rf.registers\[29\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a22o_1
XANTENNA__12159__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ datapath.rf.registers\[24\]\[3\] net758 net754 datapath.rf.registers\[22\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout892_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07139_ datapath.rf.registers\[16\]\[26\] net962 _02061_ _02063_ _02065_ vssd1 vssd1
+ vccd1 vccd1 _02066_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07586__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _04795_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or2_1
XANTENNA__10590__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ net206 _05007_ net1313 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12531__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09406__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_4_clk _00727_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ clknet_leaf_18_clk _00658_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10986__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ net211 net1798 net588 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ net217 net1948 net572 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__B2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ net226 net1815 net437 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11604_ _06067_ screen.csx _06063_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ net1759 net238 net446 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ clknet_leaf_48_clk _01210_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11535_ _05927_ _05993_ _05681_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_151_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12706__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire342 _02280_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_4
XFILLER_0_135_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14254_ clknet_leaf_1_clk _01141_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11466_ _05930_ _05931_ _05937_ _05917_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or4b_1
X_13205_ clknet_leaf_29_clk _00197_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10417_ datapath.multiplication_module.multiplier_i\[13\] datapath.multiplication_module.multiplier_i\[12\]
+ datapath.multiplication_module.multiplier_i\[15\] datapath.multiplication_module.multiplier_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14185_ clknet_leaf_105_clk _01072_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11397_ _02410_ net668 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__and2_1
XANTENNA__07577__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ clknet_leaf_1_clk _00128_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10348_ screen.counter.ct\[11\] screen.counter.ct\[10\] net1290 net1291 vssd1 vssd1
+ vccd1 vccd1 _05270_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_55_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__A1 _02831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ clknet_leaf_101_clk _00059_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10279_ _03913_ _05205_ net429 net675 vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__a211o_1
XANTENNA__08526__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ datapath.mulitply_result\[6\] net326 net322 _06299_ vssd1 vssd1 vccd1 vccd1
+ _00581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10896__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ clknet_leaf_9_clk _00856_ net1084 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_06510_ keypad.decode.q2 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__inv_2
X_07490_ datapath.rf.registers\[31\]\[18\] net949 net905 datapath.rf.registers\[24\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a22o_1
XANTENNA__06675__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10197__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09160_ net503 net619 net496 net515 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__a211o_1
XANTENNA__06825__D net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ datapath.rf.registers\[16\]\[4\] net961 _03023_ _03032_ _03037_ vssd1 vssd1
+ vccd1 vccd1 _03038_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_145_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07265__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ _03519_ _04017_ _04012_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12616__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ _02955_ _02956_ _02965_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold901 datapath.rf.registers\[24\]\[30\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 datapath.rf.registers\[27\]\[25\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold923 datapath.rf.registers\[8\]\[30\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 datapath.rf.registers\[13\]\[26\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 datapath.rf.registers\[18\]\[11\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 datapath.rf.registers\[9\]\[28\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 datapath.rf.registers\[11\]\[16\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 datapath.rf.registers\[20\]\[16\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10572__A1 _03285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold989 datapath.rf.registers\[16\]\[0\] vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _04916_ _04919_ datapath.PC\[23\] net1269 vssd1 vssd1 vccd1 vccd1 _04920_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12351__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ _03833_ _03870_ net673 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_4_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ net497 net494 net527 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout473_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07826_ datapath.rf.registers\[30\]\[10\] net908 net888 datapath.rf.registers\[12\]\[10\]
+ _02750_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a221o_1
XANTENNA__07740__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ datapath.rf.registers\[21\]\[12\] net936 net852 datapath.rf.registers\[5\]\[12\]
+ _02683_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout640_A _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout738_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ _01620_ _01635_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__or2_4
XANTENNA__11824__A1 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07688_ datapath.rf.registers\[25\]\[13\] net796 net789 datapath.rf.registers\[18\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ net639 _04347_ _04352_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_23_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06639_ mmio.memload_or_instruction\[30\] mmio.memload_or_instruction\[31\] mmio.memload_or_instruction\[27\]
+ mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_23_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ net364 _04141_ _04142_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ datapath.rf.registers\[3\]\[1\] net974 _01738_ vssd1 vssd1 vccd1 vccd1 _03236_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_35_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12526__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ net511 net352 _04215_ net388 vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10260__A0 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11320_ _05853_ net313 vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11251_ net1594 net143 net136 _02499_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08205__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net1051 _05126_ _05128_ net700 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a211o_1
X_11182_ net1493 _05828_ _05830_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11088__D _05737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ datapath.PC\[5\] _03571_ datapath.PC\[6\] vssd1 vssd1 vccd1 vccd1 _05060_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12261__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ datapath.PC\[19\] _03872_ net538 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07731__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_38_clk _00710_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11815__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ clknet_leaf_52_clk _00641_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10966_ net277 net2447 net586 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__mux2_1
X_12705_ net284 net2626 net569 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__mux2_1
X_13685_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[2\] net1228
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[2\] sky130_fd_sc_hd__dfrtp_1
X_10897_ net281 net2587 net594 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10448__C _02499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12636_ net297 net1793 net436 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12436__S net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ _05672_ net577 vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14306_ clknet_leaf_43_clk _01193_ net1181 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11518_ _05719_ _05810_ net975 vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10464__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12498_ net171 net2314 net458 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__mux2_1
Xhold208 datapath.rf.registers\[7\]\[7\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold219 datapath.rf.registers\[25\]\[2\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ clknet_leaf_32_clk _01124_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11449_ screen.register.currentXbus\[9\] net1016 net1014 screen.register.currentXbus\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a22o_1
XANTENNA__09074__A1_N net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10003__B1 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ clknet_leaf_42_clk _01055_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13119_ clknet_leaf_38_clk _00111_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07773__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14099_ clknet_leaf_48_clk _00986_ net1263 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ datapath.rf.registers\[26\]\[29\] net822 net819 datapath.rf.registers\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XANTENNA__07970__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1270 net1273 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09172__A1 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1281 screen.counter.ct\[19\] vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__clkbuf_2
X_08660_ datapath.PC\[25\] _03586_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__or2_1
Xfanout1292 screen.counter.ct\[9\] vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07722__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ datapath.rf.registers\[25\]\[15\] net797 net767 datapath.rf.registers\[3\]\[15\]
+ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a221o_1
X_08591_ net504 net622 _03517_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06930__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07542_ datapath.rf.registers\[10\]\[17\] net916 net896 datapath.rf.registers\[6\]\[17\]
+ _02468_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06836__C net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ datapath.rf.registers\[13\]\[18\] net793 net723 datapath.rf.registers\[27\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09212_ _04137_ _04138_ net370 vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09143_ _03848_ _03849_ net382 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12346__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09632__C1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06852__B _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07789__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ net636 _03986_ _03998_ net612 vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06997__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08025_ datapath.rf.registers\[0\]\[6\] net827 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1130_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 datapath.rf.registers\[6\]\[22\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 datapath.rf.registers\[24\]\[5\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 datapath.rf.registers\[24\]\[12\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 datapath.rf.registers\[23\]\[11\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold764 datapath.rf.registers\[27\]\[20\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 datapath.rf.registers\[29\]\[13\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 datapath.rf.registers\[8\]\[10\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08779__B _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 datapath.rf.registers\[26\]\[19\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07683__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ net705 _04900_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__or3_1
XANTENNA__07961__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net394 _03722_ _03723_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__a31o_1
X_08858_ net674 _03780_ _03784_ _03779_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__o22a_2
XANTENNA__07174__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07713__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ datapath.rf.registers\[4\]\[11\] net928 net872 datapath.rf.registers\[25\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a22o_1
X_08789_ _03711_ _03712_ net368 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__a21o_1
X_10820_ _01468_ net658 _05649_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_156_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10751_ net1278 datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _05591_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__10838__A2_N _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ clknet_leaf_84_clk _00423_ net1236 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ net1274 _05520_ datapath.PC\[25\] vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12421_ net1956 net244 net465 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
XANTENNA__12256__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08977__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ net1694 net247 net473 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__mux2_1
XANTENNA__06988__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ net25 net1047 net1036 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1
+ vccd1 _00317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12283_ net1817 net250 net480 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__mux2_1
XANTENNA__08729__A1 _02742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14022_ clknet_leaf_111_clk _00909_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11234_ datapath.ru.n_memwrite _05252_ _05256_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__nand3_4
X_11165_ _05761_ _05809_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07952__A2 _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _01424_ _04309_ net536 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__mux2_1
X_11096_ _05265_ net1022 vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ net841 _04662_ _04823_ _04973_ net702 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_42_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07165__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 net84 vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 screen.controlBus\[29\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
X_13806_ clknet_leaf_116_clk _00693_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12020__A datapath.mulitply_result\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11998_ _06276_ _06278_ _06275_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_133_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10459__B _02654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13737_ clknet_leaf_13_clk _00624_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10949_ net216 net2373 net592 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_70_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13668_ clknet_leaf_67_clk _00606_ net1262 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12619_ net1901 net242 net441 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13599_ clknet_leaf_87_clk net1395 net1221 vssd1 vssd1 vccd1 vccd1 datapath.ru.ack_mul_reg2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10775__A1 datapath.mulitply_result\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09378__D1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09830_ _04706_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__or2_1
Xfanout507 _03039_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
Xfanout518 _02654_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_111_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout529 _02167_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07943__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ net633 _04686_ datapath.PC\[17\] vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__o21a_1
X_06973_ datapath.rf.registers\[7\]\[30\] net957 net910 datapath.rf.registers\[30\]\[30\]
+ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a221o_1
X_08712_ _02172_ _03341_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__xor2_1
X_09692_ _03309_ _04618_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__nor2_1
X_08643_ net539 _03565_ _03566_ _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a31oi_1
XANTENNA__13671__D net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06847__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08574_ _01862_ net684 net679 _01864_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ datapath.rf.registers\[18\]\[17\] net792 net769 datapath.rf.registers\[3\]\[17\]
+ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_61_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07456_ datapath.rf.registers\[31\]\[19\] net949 net921 datapath.rf.registers\[2\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout603_A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ datapath.rf.registers\[8\]\[20\] net739 net724 datapath.rf.registers\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09126_ net419 _03836_ _04052_ net318 vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09057_ _03771_ _03983_ net382 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__mux2_1
XANTENNA__12804__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ datapath.rf.registers\[19\]\[6\] net944 net880 datapath.rf.registers\[17\]\[6\]
+ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a221o_1
Xhold550 datapath.rf.registers\[31\]\[1\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 datapath.rf.registers\[15\]\[4\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 datapath.rf.registers\[23\]\[4\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 datapath.rf.registers\[21\]\[21\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 datapath.rf.registers\[6\]\[17\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08302__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ net836 _04884_ _04885_ _04881_ net201 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_129_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ net277 net2063 net606 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__mux2_1
XANTENNA__07147__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 mmio.memload_or_instruction\[0\] vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 screen.counter.ct\[21\] vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ net153 _05873_ net128 net2615 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a22o_1
XANTENNA__09414__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1272 datapath.rf.registers\[18\]\[27\] vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 screen.register.currentXbus\[1\] vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _04664_ _05540_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_142_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ net1276 _05487_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__xor2_1
XANTENNA__10994__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11246__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14571_ net1341 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
X_11783_ net833 _04798_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08111__A2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ clknet_leaf_64_clk _00472_ net1271 vssd1 vssd1 vccd1 vccd1 datapath.PC\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_10734_ datapath.mulitply_result\[0\] net426 net658 vssd1 vssd1 vccd1 vccd1 _05578_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13453_ clknet_leaf_81_clk _00409_ net1238 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ _01485_ net710 _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_11_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12404_ net1687 net287 net467 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
X_13384_ clknet_leaf_92_clk net1382 net1202 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10596_ net1966 net513 net350 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[8\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10445__D net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12335_ net2031 net166 net479 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
XANTENNA__12714__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12266_ net164 net2204 net485 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__mux2_1
X_14005_ clknet_leaf_28_clk _00892_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11217_ net1408 net143 _05841_ vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__a21bo_1
X_12197_ _05850_ _06442_ _06426_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__a21bo_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XANTENNA__10461__C net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__07925__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
X_11148_ _05323_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_50_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11079_ net1022 _05719_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__nor2_1
XANTENNA__07138__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08350__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08638__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08102__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_07310_ datapath.rf.registers\[23\]\[22\] net934 net879 datapath.rf.registers\[29\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
X_08290_ datapath.rf.registers\[15\]\[1\] net995 _01746_ vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07310__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ net529 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07172_ datapath.rf.registers\[12\]\[25\] net736 net721 datapath.rf.registers\[28\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11945__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12624__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 net306 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_2
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
Xfanout326 net328 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
X_09813_ _04734_ _04739_ _04733_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o21bai_1
XANTENNA__07916__A2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout337 net340 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
Xfanout348 net351 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
Xfanout359 _03545_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
XANTENNA__10490__D_N net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _04669_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or2_1
X_06956_ _01877_ _01879_ _01882_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__or3_1
XANTENNA__07129__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _01717_ _04597_ _04600_ net492 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a31o_1
XANTENNA__08877__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ net999 net984 net978 _01803_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout553_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _01634_ _03552_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11228__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ _03445_ _03447_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout720_A _01782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout818_A _01747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07508_ _02434_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08488_ _03373_ _03375_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07301__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10827__B _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07439_ datapath.rf.registers\[27\]\[19\] net722 _02365_ net831 vssd1 vssd1 vccd1
+ vccd1 _02366_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12189__B1 _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09054__A0 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ _02783_ _02926_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__or3_1
XANTENNA__11936__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ _02678_ net517 net684 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ _05292_ screen.controlBus\[2\] screen.controlBus\[3\] _05301_ vssd1 vssd1
+ vccd1 vccd1 _05303_ sky130_fd_sc_hd__or4bb_1
X_12120_ _06377_ _06381_ _06384_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_107_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07080__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _06325_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__nand2_1
Xhold380 datapath.rf.registers\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07368__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 datapath.multiplication_module.multiplicand_i\[6\] vssd1 vssd1 vccd1 vccd1
+ net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ net268 net2288 net582 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
XANTENNA__10989__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 _01851_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout871 _01848_ vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_4
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_4
Xfanout893 net895 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_4
XANTENNA__11393__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ net217 net2583 net542 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
Xhold1080 datapath.rf.registers\[25\]\[16\] vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 datapath.rf.registers\[14\]\[27\] vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net1432 _05889_ net157 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12884_ net228 net2550 net551 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XANTENNA__07540__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _06233_ datapath.PC\[20\] net304 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12709__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06894__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
X_14554_ net1365 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11766_ _04663_ net304 vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__nor2_1
XANTENNA__10737__B _05208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ clknet_leaf_76_clk _00455_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_126_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10717_ datapath.PC\[30\] _05556_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__nand2_1
X_14485_ clknet_leaf_29_clk _01372_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11697_ screen.counter.currentCt\[20\] _06138_ net666 vssd1 vssd1 vccd1 vccd1 _06140_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ clknet_leaf_89_clk _00392_ net1213 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
X_10648_ datapath.PC\[20\] _05497_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_155_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11927__B1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13367_ clknet_leaf_72_clk _00352_ net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12444__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10579_ net1403 _02926_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[7\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ net1922 net250 net476 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XANTENNA__07071__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ clknet_leaf_110_clk _00288_ net1106 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12249_ net251 net2155 net484 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07359__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ _01731_ net973 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nand2_1
X_07790_ datapath.rf.registers\[5\]\[11\] net782 net726 datapath.rf.registers\[2\]\[11\]
+ _02705_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a221o_1
XANTENNA__12104__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06741_ mmio.memload_or_instruction\[8\] net1062 net1004 datapath.ru.latched_instruction\[8\]
+ net1038 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09460_ _02793_ _03403_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__xnor2_1
X_06672_ _01594_ _01600_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07531__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08411_ _02304_ _03337_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_106_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09391_ _04089_ _04090_ net374 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__a21o_1
XANTENNA__12619__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_08342_ datapath.rf.registers\[7\]\[0\] net994 _01739_ vssd1 vssd1 vccd1 vccd1 _03269_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09284__A0 _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06844__C _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ datapath.rf.registers\[19\]\[1\] net947 net855 datapath.rf.registers\[5\]\[1\]
+ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout134_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07224_ datapath.rf.registers\[31\]\[24\] net950 net695 _02150_ vssd1 vssd1 vccd1
+ vccd1 _02151_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09587__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12354__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09587__B2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _02060_ _02079_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07086_ _02008_ _02010_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11146__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
XANTENNA_fanout670_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
Xfanout156 net158 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout768_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout167 net170 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_2
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06588__A mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ datapath.rf.registers\[6\]\[7\] net813 net726 datapath.rf.registers\[2\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a22o_1
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _04652_ _04653_ _04633_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__o21a_1
XANTENNA__11449__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06939_ datapath.rf.registers\[26\]\[30\] net821 net771 datapath.rf.registers\[30\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10657__B1 _05510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ net221 _04562_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__and3_1
XANTENNA__07522__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ net982 _03121_ net617 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__mux2_1
X_09589_ _03556_ _04501_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12529__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ _01439_ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__nor2_1
XANTENNA__09275__A0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _05952_ _06012_ _06017_ net1017 _05902_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ net36 _05347_ _05411_ net35 vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_108_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14270_ clknet_leaf_52_clk _01157_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire535 _01929_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_4
X_11482_ _05811_ _05952_ _05951_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11909__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ clknet_leaf_77_clk _00212_ net1238 vssd1 vssd1 vccd1 vccd1 datapath.i_ack
+ sky130_fd_sc_hd__dfrtp_1
X_10433_ _05348_ _05349_ vssd1 vssd1 vccd1 vccd1 screen.register.controlFill sky130_fd_sc_hd__or2_1
XANTENNA__12264__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07053__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ clknet_leaf_47_clk _00144_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10364_ _01440_ _05284_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__or3_1
X_12103_ _06363_ _06369_ _06368_ _06367_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__o211ai_1
X_13083_ clknet_leaf_52_clk _00075_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ _01864_ _03438_ _03496_ _04629_ _01625_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__a2111o_1
X_12034_ _06310_ _06311_ _06312_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09750__A1 _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout690 _01829_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_6
XANTENNA__07761__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13985_ clknet_leaf_41_clk _00872_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ net283 net2393 net541 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__mux2_1
XANTENNA__07513__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ net298 net1637 net550 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__mux2_1
XANTENNA__12439__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06867__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11818_ net702 _03946_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__nand2_1
XANTENNA__08218__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12798_ net630 _06448_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14537_ net1324 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XANTENNA__06619__A2 _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ net1281 _06073_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14468_ clknet_leaf_16_clk _01355_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07292__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ clknet_leaf_89_clk _00375_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14399_ clknet_leaf_38_clk _01286_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11376__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07044__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ _03770_ _03886_ net374 vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12902__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07911_ datapath.rf.registers\[23\]\[8\] net935 net918 datapath.rf.registers\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a22o_1
X_08891_ net528 net357 _03814_ net389 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a211o_1
X_07842_ datapath.rf.registers\[22\]\[10\] net751 net744 datapath.rf.registers\[21\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07773_ _02679_ net517 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09512_ _01717_ _04438_ net492 vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a21o_1
X_06724_ datapath.ru.latched_instruction\[7\] net1038 _01649_ vssd1 vssd1 vccd1 vccd1
+ _01651_ sky130_fd_sc_hd__a21o_2
XFILLER_0_79_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11300__B2 mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net402 _04369_ net339 vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06655_ datapath.ru.latched_instruction\[0\] _01458_ net1029 vssd1 vssd1 vccd1 vccd1
+ _01585_ sky130_fd_sc_hd__mux2_1
XANTENNA__06858__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12349__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06855__B _01776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap1003_A _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09374_ net391 _04300_ _04298_ net399 vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__a211oi_1
X_06586_ net1305 net1303 mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1 vccd1
+ _01516_ sky130_fd_sc_hd__or3b_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ _03250_ _03251_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_145_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1160_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_A _02742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1258_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ datapath.rf.registers\[23\]\[1\] net932 net877 datapath.rf.registers\[29\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07207_ datapath.rf.registers\[20\]\[24\] net803 net798 datapath.rf.registers\[25\]\[24\]
+ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08187_ _03110_ _03111_ _03112_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ datapath.rf.registers\[24\]\[26\] net905 net873 datapath.rf.registers\[25\]\[26\]
+ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout885_A _01841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12812__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ _01994_ _01995_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__and2b_2
XANTENNA__07906__S net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ _04837_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or2_1
Xwire1024 _05690_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07743__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ clknet_leaf_10_clk _00657_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ net213 net1723 net588 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12721_ net223 net2427 net571 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__mux2_1
XANTENNA__12259__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net242 net1962 net437 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _05797_ _06053_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ net1652 net247 net445 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ clknet_leaf_35_clk _01209_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11534_ net1011 _06001_ _05969_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07274__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14253_ clknet_leaf_0_clk _01140_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11399__A _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11465_ _05932_ _05934_ _05936_ net1011 vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13204_ clknet_leaf_116_clk _00196_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07026__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ datapath.multiplication_module.multiplier_i\[9\] datapath.multiplication_module.multiplier_i\[8\]
+ datapath.multiplication_module.multiplier_i\[11\] datapath.multiplication_module.multiplier_i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14184_ clknet_leaf_13_clk _01071_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13443__SET_B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ screen.register.currentYbus\[17\] net130 _05883_ net159 vssd1 vssd1 vccd1
+ vccd1 _00375_ sky130_fd_sc_hd__a22o_1
X_13135_ clknet_leaf_5_clk _00127_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12722__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10347_ _05267_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ clknet_leaf_11_clk _00058_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ _03252_ _03309_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09492__A_N _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ _06297_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07734__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ clknet_leaf_0_clk _00855_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12919_ net2052 net224 net546 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
X_13899_ clknet_leaf_101_clk _00786_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08110_ net694 _03034_ _03036_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__or3_1
XANTENNA__07265__A2 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ net385 _04015_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08041_ datapath.rf.registers\[22\]\[6\] net751 _02959_ _02967_ vssd1 vssd1 vccd1
+ vccd1 _02968_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A1 _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold902 datapath.rf.registers\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 datapath.rf.registers\[9\]\[31\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07017__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 datapath.rf.registers\[3\]\[6\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 datapath.rf.registers\[21\]\[7\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold946 datapath.rf.registers\[28\]\[17\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 datapath.rf.registers\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 datapath.rf.registers\[23\]\[10\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ net201 _04918_ net1268 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__o21a_1
XANTENNA__12632__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold979 datapath.rf.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07973__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ net491 _03868_ _03869_ _03864_ _03866_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_4_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
X_08874_ net503 net619 net496 net528 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a211o_1
XANTENNA__06528__A1 mmio.memload_or_instruction\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ datapath.rf.registers\[11\]\[10\] net968 net956 datapath.rf.registers\[7\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout466_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ datapath.rf.registers\[4\]\[12\] net928 net864 datapath.rf.registers\[13\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a22o_1
X_06707_ net655 _01633_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nand2_1
X_07687_ _02611_ _02612_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__and2_2
XANTENNA__08150__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ net335 _03730_ _04350_ net640 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o211a_1
X_06638_ _01456_ _01464_ _01478_ _01501_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_23_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09357_ _04135_ _04136_ net366 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a21o_1
X_06569_ net1306 net1304 mmio.memload_or_instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ _01499_ sky130_fd_sc_hd__or3b_1
XFILLER_0_63_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12807__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08308_ datapath.rf.registers\[23\]\[1\] net991 _01739_ vssd1 vssd1 vccd1 vccd1 _03235_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09288_ net499 net620 net490 net509 vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__o211a_1
XANTENNA__10260__A1 _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08239_ datapath.rf.registers\[24\]\[2\] net758 _03151_ _03154_ _03155_ vssd1 vssd1
+ vccd1 vccd1 _03166_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_134_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11250_ net423 _05844_ net140 net1469 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07008__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10201_ _03574_ _05127_ net1051 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10012__A1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ mmio.key_data\[0\] net220 _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and3_1
XANTENNA__12542__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _01425_ _04191_ net536 vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10063_ _04473_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nand2_1
XANTENNA__07716__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10997__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ clknet_leaf_51_clk _00709_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11276__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13753_ clknet_leaf_60_clk _00640_ net1267 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10965_ net282 net2307 net586 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ net296 net2462 net570 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13684_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[1\] net1228
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07495__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10896_ net283 net2019 net595 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__mux2_1
X_12635_ net289 datapath.rf.registers\[14\]\[1\] net436 vssd1 vssd1 vccd1 vccd1 _01067_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12717__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07247__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ net165 net2458 net450 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10251__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14305_ clknet_leaf_41_clk _01192_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11517_ net1011 _05977_ _05985_ net1017 _05980_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12497_ net184 net2322 net457 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__mux2_1
XANTENNA__10464__C net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 datapath.rf.registers\[13\]\[4\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ clknet_leaf_53_clk _01123_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11448_ net1406 _05920_ _05901_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11200__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ clknet_leaf_44_clk _01054_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11379_ _02831_ net668 vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__and2_1
X_13118_ clknet_leaf_51_clk _00110_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14098_ clknet_leaf_36_clk _00985_ net1149 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13049_ clknet_leaf_47_clk _00041_ net1197 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07707__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
Xfanout1271 net1272 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__clkbuf_4
Xfanout1282 screen.counter.ct\[18\] vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1293 screen.counter.ct\[8\] vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_2
X_07610_ datapath.rf.registers\[15\]\[15\] net806 net752 datapath.rf.registers\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a22o_1
X_08590_ _01638_ net622 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__nand2_1
XANTENNA__10700__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ datapath.rf.registers\[4\]\[17\] net928 net904 datapath.rf.registers\[24\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__a22o_1
XANTENNA__11267__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11806__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06836__D _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ datapath.rf.registers\[6\]\[18\] net814 net810 datapath.rf.registers\[4\]\[18\]
+ _02398_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ _04133_ _04134_ net366 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12627__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ net378 _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nor2_1
XANTENNA__07238__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09073_ _03408_ _03979_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout214_A _05526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08024_ datapath.rf.registers\[0\]\[6\] net690 _02935_ _02950_ vssd1 vssd1 vccd1
+ vccd1 _02951_ sky130_fd_sc_hd__o22a_4
XFILLER_0_102_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold710 datapath.rf.registers\[22\]\[2\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold721 datapath.rf.registers\[2\]\[15\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 datapath.rf.registers\[6\]\[26\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 datapath.rf.registers\[7\]\[31\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12362__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold754 datapath.rf.registers\[11\]\[30\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold765 datapath.rf.registers\[28\]\[5\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 datapath.rf.registers\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 datapath.rf.registers\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _03589_ _04901_ net1053 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__a21oi_1
Xhold798 datapath.rf.registers\[8\]\[28\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_A _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ net384 _03525_ _03524_ net393 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__o211a_1
XANTENNA__07980__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ net615 _03754_ _03783_ _03782_ net676 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout750_A _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ datapath.rf.registers\[18\]\[11\] net912 net884 datapath.rf.registers\[9\]\[11\]
+ _02734_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a221o_1
X_08788_ _03713_ _03714_ net362 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11258__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ datapath.rf.registers\[25\]\[12\] net796 net718 datapath.rf.registers\[28\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a22o_1
X_10750_ net2291 net291 net605 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07477__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ _04333_ _04335_ net671 _04312_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12537__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ net1274 datapath.PC\[25\] _05520_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
X_12420_ net1946 net235 net464 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_1
XANTENNA__07229__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10233__B2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ net1788 net251 net473 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ net23 net1045 net1034 net2525 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__o22a_1
X_12282_ net2159 net254 net480 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ clknet_leaf_93_clk _00908_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11233_ datapath.ru.n_memwrite _05252_ _05256_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__and3_1
XANTENNA__12272__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09147__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ net1014 _05771_ _05812_ _05813_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__or4_1
XANTENNA__07401__A2 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10115_ _04310_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__or2_1
X_11095_ _05734_ _05738_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_147_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ _04784_ _04822_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__or2_1
Xhold70 screen.controlBus\[30\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 screen.controlBus\[22\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 net46 vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
X_13805_ clknet_leaf_119_clk _00692_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11997_ _06280_ _06281_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_67_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10459__C _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13736_ clknet_leaf_14_clk _00623_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07468__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ net217 net2421 net593 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12447__S net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ clknet_leaf_67_clk _00605_ net1259 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10879_ net219 net2548 net601 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12618_ net1865 net234 net440 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13598_ clknet_leaf_80_clk net1392 net1238 vssd1 vssd1 vccd1 vccd1 screen.register.cFill3
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10224__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12549_ net249 net2339 net448 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__mux2_1
XANTENNA__10775__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14219_ clknet_leaf_18_clk _01106_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout508 _03039_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_2
Xfanout519 _02608_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_111_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ datapath.PC\[17\] net633 _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__or3_1
XANTENNA__12910__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06972_ datapath.rf.registers\[27\]\[30\] net870 net849 datapath.rf.registers\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
X_08711_ _02172_ _03426_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__xnor2_1
X_09691_ _03288_ _03307_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__nor2_1
Xfanout1090 net1093 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
X_08642_ datapath.PC\[31\] net538 net1053 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__o21ai_1
X_08573_ net1003 _01632_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07524_ datapath.rf.registers\[31\]\[17\] net817 _02449_ _02450_ vssd1 vssd1 vccd1
+ vccd1 _02451_ sky130_fd_sc_hd__a211o_1
XANTENNA__07459__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07024__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07455_ datapath.rf.registers\[3\]\[19\] net965 net873 datapath.rf.registers\[25\]\[19\]
+ _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12357__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout429_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07386_ _02306_ _02308_ _02310_ _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__or4_1
XANTENNA__08136__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09125_ net419 _03840_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__nand2_1
XANTENNA_hold1279_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09056_ _03886_ _03982_ net374 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07631__A2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11497__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ datapath.rf.registers\[3\]\[6\] net964 net848 datapath.rf.registers\[1\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout798_A _01755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold540 datapath.rf.registers\[4\]\[20\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 datapath.rf.registers\[7\]\[19\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 datapath.rf.registers\[17\]\[14\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 datapath.mulitply_result\[30\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 datapath.rf.registers\[5\]\[26\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold595 datapath.rf.registers\[20\]\[21\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__C _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _01715_ _03637_ _04882_ net1052 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_129_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _03465_ _03469_ net413 vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09889_ _04760_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__xnor2_1
Xhold1240 screen.register.currentXbus\[31\] vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 screen.register.currentXbus\[11\] vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ net154 _05872_ net129 net2537 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a22o_1
Xhold1262 keypad.apps.app_c\[0\] vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 screen.register.currentXbus\[2\] vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__B1 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1284 screen.register.currentYbus\[2\] vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11851_ _04999_ net305 vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_142_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ net1615 net261 net602 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__mux2_1
X_14570_ net1340 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
X_11782_ net699 _04359_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__nand2_1
X_10733_ datapath.PC\[0\] _05234_ net839 vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13521_ clknet_leaf_64_clk _00471_ net1271 vssd1 vssd1 vccd1 vccd1 datapath.PC\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13452_ clknet_leaf_81_clk _00408_ net1238 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10664_ datapath.mulitply_result\[22\] net427 _05513_ _05517_ net660 vssd1 vssd1
+ vccd1 vccd1 _05518_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_11_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07870__A2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ net1567 net180 net464 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_90_clk _00357_ net1209 vssd1 vssd1 vccd1 vccd1 keypad.alpha sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10595_ net1757 net512 net350 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[7\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14438__RESET_B net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07083__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12334_ net1772 net167 net478 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07622__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ net168 net2161 net485 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ clknet_leaf_115_clk _00891_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11216_ _01404_ _05256_ _05838_ _05019_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a211o_1
X_12196_ columns.count\[9\] _01445_ _06433_ columns.count\[10\] vssd1 vssd1 vccd1
+ vccd1 _06442_ sky130_fd_sc_hd__a31o_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XANTENNA__08583__A0 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__10461__D net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
X_11147_ _05309_ net1017 vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__or2_1
XANTENNA__12730__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11078_ _05701_ _05718_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__or2_2
X_10029_ datapath.PC\[20\] _03831_ net538 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__mux2_1
XANTENNA__07689__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11890__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ clknet_leaf_88_clk datapath.multiplication_module.multiplier_i_n\[4\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10486__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07240_ datapath.rf.registers\[0\]\[24\] _01829_ _02152_ _02166_ vssd1 vssd1 vccd1
+ vccd1 _02167_ sky130_fd_sc_hd__o22a_2
XFILLER_0_144_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07171_ _02092_ _02093_ _02095_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12905__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09063__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10748__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07074__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08810__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07613__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_2
Xfanout316 _03549_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08574__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ datapath.PC\[0\] _03286_ _04738_ _04736_ vssd1 vssd1 vccd1 vccd1 _04739_
+ sky130_fd_sc_hd__a31oi_2
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
XANTENNA__12640__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout338 net340 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_1
Xfanout349 net351 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11764__B _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ net1274 net629 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nor2_1
X_06955_ _01867_ _01868_ _01875_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ net315 _04598_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__or2_1
X_06886_ net999 net983 net978 _01812_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__and4_1
X_08625_ _01593_ _01602_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__nor2_2
XANTENNA__06888__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1190_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ _03445_ _03447_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07507_ _02411_ _02431_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ _02523_ _03413_ _02524_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07438_ datapath.rf.registers\[19\]\[19\] net759 net718 datapath.rf.registers\[28\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07852__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09054__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07369_ datapath.rf.registers\[25\]\[21\] net873 net858 datapath.rf.registers\[15\]\[21\]
+ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a221o_1
XANTENNA__12815__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ net415 _03796_ _04034_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__o21ai_2
X_10380_ _05292_ screen.controlBus\[2\] screen.controlBus\[3\] _05301_ vssd1 vssd1
+ vccd1 vccd1 _05302_ sky130_fd_sc_hd__and4bb_1
XANTENNA__08801__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09039_ _03718_ _03965_ net381 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__mux2_1
X_12050_ datapath.mulitply_result\[12\] datapath.multiplication_module.multiplicand_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__or2_1
Xhold370 datapath.rf.registers\[24\]\[24\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 datapath.rf.registers\[10\]\[23\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net271 net2110 net584 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
Xhold392 datapath.rf.registers\[30\]\[15\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12550__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 _01851_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09109__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout872 net875 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
Xfanout883 _01843_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
X_12952_ net223 net2392 net543 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
XANTENNA__10124__B1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1070 datapath.rf.registers\[15\]\[6\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 datapath.rf.registers\[29\]\[7\] vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ _05888_ _06263_ net149 net1447 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__a22o_1
Xhold1092 datapath.rf.registers\[11\]\[31\] vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_47_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ net244 net2520 net551 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ net837 _03831_ _04664_ _05505_ _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553_ net1364 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
X_11765_ net699 _04789_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__or2_1
XANTENNA__08096__A2 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13504_ clknet_leaf_78_clk _00454_ net1247 vssd1 vssd1 vccd1 vccd1 datapath.PC\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_60_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ net174 net2287 net608 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14484_ clknet_leaf_115_clk _01371_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07843__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11696_ net666 _06137_ _06139_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13435_ clknet_leaf_89_clk _00391_ net1210 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
X_10647_ datapath.PC\[20\] _05497_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and2_1
XANTENNA__12725__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11927__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ clknet_leaf_96_clk _00351_ net1218 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ net1390 _02971_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[6\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09450__D1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ net2157 net254 net476 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__mux2_1
X_13297_ clknet_leaf_112_clk _00287_ net1094 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08223__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ net253 net2459 net484 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12179_ _05849_ _06426_ columns.count\[4\] vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__a21o_1
XANTENNA__08020__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12104__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ mmio.memload_or_instruction\[10\] net1061 net1006 datapath.ru.latched_instruction\[10\]
+ net1039 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__a32o_1
XFILLER_0_155_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06671_ _01584_ _01588_ _01598_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_35_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08410_ _02349_ _02390_ _03334_ _02345_ _02302_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_106_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09390_ net365 _04202_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a21o_1
X_14526__1317 vssd1 vssd1 vccd1 vccd1 _14526__1317/HI net1317 sky130_fd_sc_hd__conb_1
X_08341_ datapath.rf.registers\[31\]\[0\] net989 _01746_ vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08087__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09284__A1 _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08272_ datapath.rf.registers\[20\]\[1\] net903 net872 datapath.rf.registers\[25\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07295__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__A2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07223_ datapath.rf.registers\[23\]\[24\] net934 net915 datapath.rf.registers\[18\]\[24\]
+ _02149_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12635__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout127_A _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07047__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07154_ _02060_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__or2_2
XFILLER_0_14_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07085_ datapath.rf.registers\[6\]\[27\] net815 net806 datapath.rf.registers\[15\]\[27\]
+ _02011_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08011__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1203_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
Xfanout168 net170 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_2
X_07987_ datapath.rf.registers\[7\]\[7\] net824 net820 datapath.rf.registers\[26\]\[7\]
+ _02913_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a221o_1
Xfanout179 _06182_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09726_ _02259_ _03367_ _03422_ _04635_ _03366_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a221o_1
X_06938_ datapath.rf.registers\[20\]\[30\] net803 net731 datapath.rf.registers\[16\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a22o_1
XANTENNA__10657__A1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ net674 _04579_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a31oi_4
X_06869_ datapath.rf.registers\[4\]\[31\] net811 net742 datapath.rf.registers\[1\]\[31\]
+ _01768_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout928_A _01820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08608_ _01656_ _03120_ net617 vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__mux2_1
X_09588_ _04509_ _04514_ net615 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08539_ _03462_ _03465_ net414 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XANTENNA__08078__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A1 _02997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11550_ screen.register.currentXbus\[22\] net1015 net1013 screen.register.currentXbus\[30\]
+ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_42_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07825__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10501_ net36 _05346_ _05411_ net35 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__and4b_1
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12545__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ net975 _05813_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__or2_1
Xwire525 _02323_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_4
XANTENNA__10854__A _01650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13220_ clknet_leaf_90_clk net1497 net1209 vssd1 vssd1 vccd1 vccd1 keypad.decode.push
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10432_ screen.controlBus\[0\] _05284_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10042__C1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ clknet_leaf_38_clk _00143_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10363_ screen.controlBus\[2\] screen.controlBus\[3\] vssd1 vssd1 vccd1 vccd1 _05285_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07994__D1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ _06367_ _06368_ _06369_ _06363_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ clknet_leaf_23_clk _00074_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ _03310_ net686 _05213_ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_57_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12033_ datapath.mulitply_result\[9\] datapath.multiplication_module.multiplicand_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__and2_1
XANTENNA__12280__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _03499_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
Xfanout691 _01829_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12098__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ clknet_leaf_47_clk _00871_ net1195 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12935_ net295 net1938 net542 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__mux2_1
X_12866_ net290 net1646 net550 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11817_ _06218_ _06219_ _06220_ net303 datapath.PC\[15\] vssd1 vssd1 vccd1 vccd1
+ _00459_ sky130_fd_sc_hd__a32o_1
X_12797_ net163 net2254 net563 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07277__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536_ net1323 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_11748_ net1283 net664 _06169_ net713 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14467_ clknet_leaf_104_clk _01354_ net1120 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12455__S net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ screen.counter.currentCt\[14\] _06126_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13418_ clknet_leaf_88_clk _00374_ net1215 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14398_ clknet_leaf_52_clk _01285_ net1176 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11376__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10033__C1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08241__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ clknet_leaf_100_clk _00334_ net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07910_ datapath.rf.registers\[20\]\[8\] net902 net890 datapath.rf.registers\[12\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a22o_1
X_08890_ net526 net356 _03815_ net385 vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__a211o_1
X_07841_ datapath.rf.registers\[6\]\[10\] net813 net809 datapath.rf.registers\[4\]\[10\]
+ _02765_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07772_ _02678_ net517 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__nand2_1
X_06723_ datapath.ru.latched_instruction\[7\] net1037 _01649_ vssd1 vssd1 vccd1 vccd1
+ _01650_ sky130_fd_sc_hd__a21oi_4
X_09511_ net637 _04429_ _04436_ _04437_ net656 vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07504__A1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11300__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09442_ _04017_ _04300_ net397 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06654_ datapath.ru.latched_instruction\[6\] net1042 net1009 _01582_ vssd1 vssd1
+ vccd1 vccd1 _01584_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09373_ net385 _04164_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__o21ai_1
X_06585_ net1305 net1303 mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ _01515_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout244_A _05496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ net651 _03244_ _03245_ _03202_ _03204_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07268__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10811__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08255_ net505 net504 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__xor2_4
XANTENNA__12365__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1153_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A _02997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07206_ datapath.rf.registers\[6\]\[24\] net815 net807 datapath.rf.registers\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
X_08186_ datapath.rf.registers\[8\]\[3\] net737 _03094_ _03096_ _03098_ vssd1 vssd1
+ vccd1 vccd1 _03113_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_119_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07137_ datapath.rf.registers\[12\]\[26\] net889 net862 datapath.rf.registers\[28\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07068_ _01972_ _01991_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A _01844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08310__C _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _04634_ _03748_ _02349_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__or3b_1
X_10981_ net218 net1944 net588 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12720_ net233 net2631 net572 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ net235 net2396 net439 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _05295_ _06059_ _06062_ _05307_ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__o221a_1
XANTENNA__07259__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ net1849 net252 net444 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ clknet_leaf_8_clk _01208_ net1084 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11533_ screen.register.currentYbus\[21\] _05775_ _05997_ _05999_ _06000_ vssd1 vssd1
+ vccd1 vccd1 _06001_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12275__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire344 _01884_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_152_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11399__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ screen.register.currentYbus\[25\] _05777_ _05935_ vssd1 vssd1 vccd1 vccd1
+ _05936_ sky130_fd_sc_hd__a21o_1
X_14252_ clknet_leaf_31_clk _01139_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08759__A0 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10415_ datapath.multiplication_module.multiplier_i\[1\] datapath.multiplication_module.multiplier_i\[0\]
+ datapath.multiplication_module.multiplier_i\[3\] datapath.multiplication_module.multiplier_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13203_ clknet_leaf_61_clk _00195_ net1266 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11395_ _02456_ net668 vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__and2_1
X_14183_ clknet_leaf_25_clk _01070_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10346_ net1284 net1285 net1281 net1282 vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__or4_1
X_13134_ clknet_leaf_118_clk _00126_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525__1316 vssd1 vssd1 vccd1 vccd1 _14525__1316/HI net1316 sky130_fd_sc_hd__conb_1
XANTENNA__06785__A2 _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ clknet_leaf_105_clk _00057_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10277_ _05192_ _05195_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__and3b_1
X_12016_ _06290_ _06291_ _06292_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09184__B1 _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13967_ clknet_leaf_5_clk _00854_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07498__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ net2138 net232 net547 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__B2 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13898_ clknet_leaf_10_clk _00785_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09239__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ net234 net2388 net553 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14519_ net1308 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08040_ datapath.rf.registers\[13\]\[6\] net795 net755 datapath.rf.registers\[24\]\[6\]
+ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07670__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 datapath.rf.registers\[28\]\[11\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold914 datapath.rf.registers\[20\]\[11\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12913__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold925 datapath.rf.registers\[25\]\[3\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 datapath.rf.registers\[6\]\[0\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 datapath.rf.registers\[12\]\[6\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 datapath.rf.registers\[1\]\[14\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 datapath.rf.registers\[16\]\[10\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _04832_ _04917_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08942_ net642 _03868_ _03867_ _03356_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ net369 _03676_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07824_ datapath.rf.registers\[16\]\[10\] net960 net924 datapath.rf.registers\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a22o_1
X_07755_ datapath.rf.registers\[19\]\[12\] net944 net908 datapath.rf.registers\[30\]\[12\]
+ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a221o_1
X_06706_ _01633_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__inv_2
XANTENNA__07489__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__B2 mmio.memload_or_instruction\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__inv_2
XANTENNA__08139__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06637_ mmio.memload_or_instruction\[19\] mmio.memload_or_instruction\[21\] mmio.memload_or_instruction\[22\]
+ mmio.memload_or_instruction\[20\] vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__and4bb_1
X_09425_ _02932_ net680 _03736_ net320 _04351_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1270_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06568_ _01409_ _01456_ _01478_ _01408_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ _04237_ _04238_ net361 vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08989__B1 _03552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ datapath.rf.registers\[26\]\[1\] net823 net783 datapath.rf.registers\[5\]\[1\]
+ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ net386 _04211_ _04212_ net392 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o211a_1
X_06499_ datapath.PC\[21\] vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
X_08238_ datapath.rf.registers\[22\]\[2\] net754 net745 datapath.rf.registers\[21\]\[2\]
+ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07661__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout995_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ datapath.rf.registers\[3\]\[3\] net973 _01738_ vssd1 vssd1 vccd1 vccd1 _03096_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08205__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12823__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ datapath.PC\[8\] _03573_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__nand2_1
XANTENNA__07413__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11180_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08602__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__A2 _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ datapath.PC\[7\] net1245 _05054_ _05057_ vssd1 vssd1 vccd1 vccd1 _05058_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10062_ _03871_ _04472_ net704 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09433__A _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13821_ clknet_leaf_23_clk _00708_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13752_ clknet_leaf_42_clk _00639_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10964_ net283 net2438 net589 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__mux2_1
X_12703_ net293 net2523 net570 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[0\] net1224
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[0\] sky130_fd_sc_hd__dfrtp_1
X_10895_ net296 net1910 net595 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12634_ net182 net1526 net439 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12565_ net167 net2120 net449 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__mux2_1
XANTENNA__10787__B1 _05620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14304_ clknet_leaf_50_clk _01191_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11516_ screen.register.currentXbus\[12\] net1016 _05742_ screen.register.currentYbus\[28\]
+ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07652__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12496_ net190 net2125 net458 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ clknet_leaf_19_clk _01122_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10464__D net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12733__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11447_ _05903_ _05904_ _05911_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07404__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ screen.register.currentYbus\[8\] net131 _05874_ net160 vssd1 vssd1 vccd1
+ vccd1 _00366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14166_ clknet_leaf_26_clk _01053_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10329_ mmio.WEN _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__nand2b_1
X_13117_ clknet_leaf_24_clk _00109_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap424_A _02104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14097_ clknet_leaf_7_clk _00984_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08231__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ clknet_leaf_39_clk _00040_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_4
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
Xfanout1272 net1273 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__clkbuf_2
Xfanout1283 screen.counter.ct\[18\] vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_1
Xfanout1294 screen.counter.ct\[6\] vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__buf_2
XANTENNA__07183__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08380__B2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ datapath.rf.registers\[16\]\[17\] net960 net944 datapath.rf.registers\[19\]\[17\]
+ _02466_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07471_ datapath.rf.registers\[7\]\[18\] net825 net821 datapath.rf.registers\[26\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a22o_1
XANTENNA__09997__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12908__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08683__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ _04135_ _04136_ net361 vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07891__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ _03963_ _04067_ net374 vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09072_ net653 _03987_ _03997_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__or4_1
XANTENNA__07643__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08023_ datapath.rf.registers\[30\]\[6\] net908 _02937_ _02944_ _02949_ vssd1 vssd1
+ vccd1 vccd1 _02950_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06997__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold700 datapath.rf.registers\[24\]\[2\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12643__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold711 datapath.rf.registers\[7\]\[16\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold722 datapath.rf.registers\[11\]\[20\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold733 datapath.rf.registers\[4\]\[29\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11767__B net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold744 datapath.rf.registers\[30\]\[9\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 datapath.rf.registers\[27\]\[30\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 datapath.rf.registers\[18\]\[6\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 datapath.rf.registers\[29\]\[25\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 datapath.rf.registers\[11\]\[9\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 datapath.rf.registers\[30\]\[5\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ datapath.PC\[27\] _03588_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__nand2_1
XANTENNA__09148__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net637 _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout576_A _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11783__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__B _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ net634 _03773_ _03774_ net610 vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07174__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ datapath.rf.registers\[16\]\[11\] net960 net868 datapath.rf.registers\[27\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
X_08787_ net497 net494 net528 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11258__B2 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ datapath.rf.registers\[23\]\[12\] net786 net774 datapath.rf.registers\[11\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout910_A _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ datapath.rf.registers\[31\]\[14\] net948 net944 datapath.rf.registers\[19\]\[14\]
+ _02595_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a221o_1
XANTENNA__12818__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14524__1315 vssd1 vssd1 vccd1 vccd1 _14524__1315/HI net1315 sky130_fd_sc_hd__conb_1
XANTENNA__06685__A1 mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ net613 _04315_ _04334_ _04330_ net671 vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__o311a_1
X_10680_ net209 net1736 net608 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__mux2_1
XANTENNA__07882__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ _04258_ _04263_ net336 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ net1835 net255 net472 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__mux2_1
XANTENNA__07634__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__A2_N _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08831__C1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14539__1326 vssd1 vssd1 vccd1 vccd1 _14539__1326/HI net1326 sky130_fd_sc_hd__conb_1
X_11301_ net22 net1044 net1033 mmio.memload_or_instruction\[28\] vssd1 vssd1 vccd1
+ vccd1 _00315_ sky130_fd_sc_hd__o22a_1
X_12281_ net1909 net258 net480 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__mux2_1
XANTENNA__12553__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14020_ clknet_leaf_16_clk _00907_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09387__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ net1424 net146 _05840_ _04868_ vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__a22o_1
XANTENNA__09428__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ _05725_ _05806_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09139__A0 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _04232_ _04277_ _04309_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__a21oi_1
X_11094_ net1016 _05743_ net1014 _05741_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_147_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10045_ net834 _04969_ _04971_ _04967_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 keypad.apps.button\[4\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 net49 vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 keypad.decode.sticky\[4\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net71 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ clknet_leaf_30_clk _00691_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__B2 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11996_ datapath.mulitply_result\[3\] datapath.multiplication_module.multiplicand_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__nor2_1
XANTENNA__09311__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13735_ clknet_leaf_18_clk _00622_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10459__D _02742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12728__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10947_ net223 net2091 net592 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13666_ clknet_leaf_67_clk _00604_ net1262 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ net223 net2397 net600 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ net2532 net240 net442 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13597_ clknet_leaf_80_clk net1373 net1238 vssd1 vssd1 vccd1 vccd1 screen.register.cFill2
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07625__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ net254 net2568 net448 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12463__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _01749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net266 net2118 net456 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__mux2_1
XANTENNA__09378__B1 _04304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ clknet_leaf_10_clk _01105_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ clknet_leaf_94_clk _01036_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout509 _02997_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_111_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06971_ _01891_ _01893_ _01895_ _01897_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__or4_1
X_08710_ _03598_ _03636_ net673 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__mux2_2
X_09690_ _03068_ _04311_ _04614_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__and4_1
Xfanout1080 net1085 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_2
X_08641_ datapath.i_ack datapath.pc_module.i_ack2 vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__nand2b_1
Xfanout1091 net1093 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ net1003 _01632_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07523_ datapath.rf.registers\[30\]\[17\] net770 net748 datapath.rf.registers\[10\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
XANTENNA__12638__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ datapath.rf.registers\[6\]\[19\] net897 net860 datapath.rf.registers\[28\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07385_ datapath.rf.registers\[12\]\[20\] net736 net716 datapath.rf.registers\[29\]\[20\]
+ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09124_ _02787_ _03321_ _04048_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_98_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09055_ net367 _03981_ _03980_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a21o_1
XANTENNA__12373__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ datapath.rf.registers\[11\]\[6\] net968 net924 datapath.rf.registers\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a22o_1
Xhold530 datapath.rf.registers\[24\]\[3\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold541 datapath.rf.registers\[31\]\[10\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold552 datapath.rf.registers\[22\]\[24\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 datapath.rf.registers\[28\]\[12\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold574 datapath.rf.registers\[30\]\[13\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 datapath.rf.registers\[6\]\[2\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 datapath.rf.registers\[14\]\[18\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08592__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ _03637_ _04585_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout860_A _01851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ net421 _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_129_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__and2b_1
XANTENNA__07147__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1230 datapath.rf.registers\[31\]\[26\] vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 datapath.rf.registers\[0\]\[22\] vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 datapath.rf.registers\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ net368 _03711_ _03712_ _03765_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a31o_1
Xhold1263 screen.register.currentYbus\[30\] vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1274 screen.register.currentXbus\[22\] vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
X_11850_ net206 _04778_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _01518_ net709 _05632_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__o22a_2
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ datapath.PC\[6\] net302 _06191_ _06193_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__a22o_1
X_13520_ clknet_leaf_64_clk _00470_ net1271 vssd1 vssd1 vccd1 vccd1 datapath.PC\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_10732_ _05479_ net630 _05575_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13451_ clknet_leaf_81_clk _00407_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ net842 _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12402_ _05669_ _06445_ _06450_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__nor3_1
XANTENNA__07607__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ clknet_leaf_90_clk net1449 net1209 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10594_ net1558 net510 net350 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[6\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12333_ net2099 net171 net479 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XANTENNA__12283__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12264_ net173 net2370 net486 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14003_ clknet_leaf_49_clk _00890_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08032__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ net1433 net145 net138 _04987_ vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__a22o_1
X_12195_ _06436_ _06441_ _05851_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a21oi_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__08583__A1 _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_11146_ _05682_ _05745_ _05746_ _05795_ net1011 vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a32o_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__clkbuf_4
X_11077_ net1022 _05721_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__nor2_1
XANTENNA__07138__A2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _03831_ _04473_ net837 vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08099__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12458__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ datapath.multiplication_module.multiplier_i\[0\] datapath.multiplication_module.multiplicand_i\[0\]
+ datapath.mulitply_result\[0\] vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__a21oi_1
X_13718_ clknet_leaf_88_clk datapath.multiplication_module.multiplier_i_n\[3\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07846__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10486__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07310__A2 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13649_ clknet_leaf_100_clk _00587_ net1223 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__A0 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07170_ datapath.rf.registers\[14\]\[25\] net801 net761 datapath.rf.registers\[19\]\[25\]
+ _02096_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08810__A2 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09068__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12921__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 _06178_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_2
X_09811_ datapath.PC\[1\] _03208_ _03209_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__or3_1
Xfanout317 _03484_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
X_14523__1314 vssd1 vssd1 vccd1 vccd1 _14523__1314/HI net1314 sky130_fd_sc_hd__conb_1
Xfanout328 _06269_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
X_09742_ net1274 net629 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and2_1
X_06954_ datapath.rf.registers\[3\]\[30\] net767 net741 datapath.rf.registers\[1\]\[30\]
+ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a221o_1
XANTENNA__07129__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _03513_ _04598_ _04599_ net638 net656 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__o221a_1
X_06885_ _01672_ _01674_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__o22a_2
X_08624_ net637 _03548_ _03550_ _03503_ net657 vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__o2111a_1
X_14538__1325 vssd1 vssd1 vccd1 vccd1 _14538__1325/HI net1325 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_38_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07750__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__A _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _03478_ _03481_ net414 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout441_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12368__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _02411_ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__or2_1
X_08486_ _03376_ _03412_ _03377_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07301__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07437_ datapath.rf.registers\[10\]\[19\] net749 net731 datapath.rf.registers\[16\]\[19\]
+ _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout706_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ datapath.rf.registers\[7\]\[21\] net957 net862 datapath.rf.registers\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
X_09107_ net415 _03790_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__nand2_1
XANTENNA__08262__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07299_ datapath.rf.registers\[13\]\[22\] net794 _02225_ net832 vssd1 vssd1 vccd1
+ vccd1 _02226_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09038_ net372 _03963_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08313__C _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 datapath.rf.registers\[9\]\[0\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 datapath.rf.registers\[22\]\[16\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07368__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 datapath.rf.registers\[25\]\[0\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net275 net2238 net583 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__mux2_1
Xhold393 datapath.rf.registers\[12\]\[16\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08610__A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_2
Xfanout851 _01856_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout862 _01851_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout873 net874 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_4
Xfanout884 _01841_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08317__A1 datapath.rf.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 _01838_ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__buf_4
X_12951_ net232 net2625 net542 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
Xhold1060 datapath.rf.registers\[4\]\[28\] vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 datapath.rf.registers\[24\]\[20\] vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net1435 _05887_ net157 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
Xhold1082 datapath.rf.registers\[9\]\[22\] vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 datapath.rf.registers\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net234 net1931 net549 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
XANTENNA__07540__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07660__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ net208 _04783_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__nand2_1
XANTENNA__10587__A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14552_ net1363 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
X_11764_ net699 _04232_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ clknet_leaf_76_clk _00453_ net1248 vssd1 vssd1 vccd1 vccd1 datapath.PC\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10715_ _01487_ net661 _05560_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__o2bb2a_1
X_14483_ clknet_leaf_49_clk _01370_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11695_ _06138_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__inv_2
X_13434_ clknet_leaf_85_clk _00390_ net1254 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
X_10646_ net229 net2181 net607 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ clknet_leaf_100_clk _00350_ net1224 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10577_ datapath.multiplication_module.multiplier_i\[6\] _03017_ net347 vssd1 vssd1
+ vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[5\] sky130_fd_sc_hd__mux2_1
XANTENNA__09450__C1 _04376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net1974 net258 net476 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
X_13296_ clknet_leaf_92_clk _00286_ net1202 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08223__C _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ net258 net2517 net484 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__mux2_1
XANTENNA__12741__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07359__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ _05849_ _06426_ _06429_ net1908 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__o2bb2a_1
X_11129_ _05704_ _05772_ _05774_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06670_ _01583_ net847 vssd1 vssd1 vccd1 vccd1 datapath.MemWrite sky130_fd_sc_hd__and2_1
XANTENNA__07531__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06694__B _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ datapath.rf.registers\[18\]\[0\] _01741_ net972 vssd1 vssd1 vccd1 vccd1 _03267_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07819__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ datapath.rf.registers\[28\]\[1\] net861 _03197_ vssd1 vssd1 vccd1 vccd1 _03198_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12916__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ datapath.rf.registers\[24\]\[24\] net906 net887 datapath.rf.registers\[9\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07153_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08244__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11121__A _05705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ datapath.rf.registers\[14\]\[27\] net801 net794 datapath.rf.registers\[13\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12651__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1029_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _05843_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_4
Xfanout158 _05262_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_2
X_07986_ datapath.rf.registers\[15\]\[7\] net805 net722 datapath.rf.registers\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a22o_1
Xfanout169 net170 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_126_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ _04636_ _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__nor2_1
X_06937_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__nand2_2
XANTENNA__11303__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ net673 _04565_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06868_ datapath.rf.registers\[20\]\[31\] net802 net752 datapath.rf.registers\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07522__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ net997 _03062_ net617 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__mux2_1
X_09587_ net634 _04510_ _04512_ net612 vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o22a_1
X_06799_ _01602_ net839 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__nand2_2
X_08538_ _03463_ _03464_ net409 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08308__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _03066_ _03394_ _03392_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__a21o_1
XANTENNA__12826__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10500_ _05341_ _05342_ _05343_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ net1011 _05944_ _05950_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a21o_1
XANTENNA__08605__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11909__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08235__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ screen.controlBus\[1\] _05279_ _05285_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_137_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07589__A2 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ clknet_leaf_51_clk _00142_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10362_ _05280_ _05281_ _05282_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or4_2
XANTENNA__10593__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _06362_ _06364_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__nor2_1
X_10293_ _05218_ _05219_ _03506_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__a21o_1
XANTENNA__12561__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ clknet_leaf_60_clk _00073_ net1264 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12032_ datapath.mulitply_result\[9\] datapath.multiplication_module.multiplicand_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__nor2_1
XANTENNA__09735__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 datapath.rf.registers\[26\]\[1\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout670 net672 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07761__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout681 net682 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12098__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout692 net693 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_8
X_13983_ clknet_leaf_36_clk _00870_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12934_ net293 net1791 net541 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07513__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12865_ net183 net1878 net549 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__mux2_1
X_11816_ _04664_ _05651_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__or2_1
XANTENNA__10110__A _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12796_ net169 net2336 net564 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14535_ net1322 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
X_11747_ net1283 _06085_ _06073_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12736__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14466_ clknet_leaf_51_clk _01353_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11678_ net667 _06125_ _06127_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__and3_1
XANTENNA__09018__A2 _03940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ clknet_leaf_87_clk _00373_ net1219 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ datapath.PC\[11\] _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14397_ clknet_leaf_33_clk _01284_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13348_ clknet_leaf_99_clk _00333_ net1227 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10584__A1 _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14537__1324 vssd1 vssd1 vccd1 vccd1 _14537__1324/HI net1324 sky130_fd_sc_hd__conb_1
XANTENNA__12471__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ clknet_leaf_78_clk _00269_ net1246 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08250__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ datapath.rf.registers\[20\]\[10\] net804 net786 datapath.rf.registers\[23\]\[10\]
+ _02766_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07771_ datapath.rf.registers\[0\]\[12\] net690 _02685_ _02697_ vssd1 vssd1 vccd1
+ vccd1 _02698_ sky130_fd_sc_hd__o22a_4
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06960__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ net640 _04424_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__nand2_1
X_06722_ _01470_ net1028 net1004 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_56_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11836__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__B2 _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08701__A1 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09441_ net402 _03934_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__nor2_1
X_06653_ datapath.ru.latched_instruction\[6\] net1042 net1009 _01582_ vssd1 vssd1
+ vccd1 vccd1 _01583_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_121_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09372_ _02742_ net356 _04169_ net389 vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__a211o_1
X_06584_ mmio.memload_or_instruction\[9\] net1061 vssd1 vssd1 vccd1 vccd1 _01514_
+ sky130_fd_sc_hd__and2_1
X_08323_ _03202_ _03204_ _03244_ net647 _03211_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12646__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout237_A _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ net505 net504 vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_145_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07205_ datapath.rf.registers\[22\]\[24\] net753 net742 datapath.rf.registers\[1\]\[24\]
+ _02131_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08185_ datapath.rf.registers\[2\]\[3\] net726 _03099_ _03100_ _03102_ vssd1 vssd1
+ vccd1 vccd1 _03112_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_65_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07136_ datapath.rf.registers\[4\]\[26\] net930 net886 datapath.rf.registers\[9\]\[26\]
+ _02062_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a221o_1
XANTENNA__10575__A1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _01972_ _01991_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__nor2_1
XANTENNA__12381__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07991__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ datapath.rf.registers\[16\]\[7\] net960 net952 datapath.rf.registers\[22\]\[7\]
+ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_74_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06951__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__inv_2
X_10980_ net222 net2332 net587 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__mux2_1
X_09639_ net642 _04565_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__nand2_1
X_12650_ net239 net2466 net438 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _05297_ _06051_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12556__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ net1915 net253 net444 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ clknet_leaf_0_clk _01207_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ screen.register.currentXbus\[5\] _05704_ _05707_ screen.register.currentXbus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__a22o_1
Xwire301 _04040_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_83_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08208__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14251_ clknet_leaf_18_clk _01138_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11463_ screen.register.currentXbus\[17\] _05707_ _05709_ screen.register.currentXbus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08759__A1 _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13202_ clknet_leaf_34_clk _00194_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10414_ datapath.multiplication_module.multiplier_i\[5\] datapath.multiplication_module.multiplier_i\[4\]
+ datapath.multiplication_module.multiplier_i\[7\] datapath.multiplication_module.multiplier_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14182_ clknet_leaf_114_clk _01069_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11394_ screen.register.currentYbus\[16\] net131 _05882_ net160 vssd1 vssd1 vccd1
+ vccd1 _00374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13133_ clknet_leaf_119_clk _00125_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12291__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ net1279 net1280 screen.counter.ct\[22\] vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__or3_1
XANTENNA__10804__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ clknet_leaf_13_clk _00056_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _05201_ _05202_ _03506_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ _06295_ _06296_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nand2_1
XANTENNA__07195__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06942__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13966_ clknet_leaf_115_clk _00853_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12917_ net1877 net226 net546 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
X_13897_ clknet_leaf_2_clk _00784_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08229__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ net240 net2344 net555 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12466__S net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ net253 net2533 net561 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14518_ net1308 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ clknet_leaf_8_clk _01336_ net1084 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 datapath.rf.registers\[27\]\[3\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold915 datapath.rf.registers\[10\]\[2\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 datapath.rf.registers\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap645 _03195_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_1
Xhold937 datapath.rf.registers\[24\]\[27\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 datapath.rf.registers\[9\]\[29\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 datapath.multiplication_module.multiplicand_i\[1\] vssd1 vssd1 vccd1 vccd1
+ net2325 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _04782_ _04829_ _04831_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07973__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _03333_ _03832_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08872_ _03792_ _03794_ _03798_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__and3_1
XANTENNA__07186__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ datapath.rf.registers\[29\]\[10\] net876 net852 datapath.rf.registers\[5\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout187_A _05555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07754_ datapath.rf.registers\[3\]\[12\] net964 net932 datapath.rf.registers\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a22o_1
X_06705_ _01625_ _01632_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nor2_4
X_07685_ _02588_ _02609_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__nand2_1
XANTENNA__08150__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08139__B _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _02929_ net683 _03494_ _02928_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06636_ mmio.memload_or_instruction\[15\] mmio.memload_or_instruction\[16\] vssd1
+ vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09355_ _03067_ net680 _03797_ net320 _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a221o_1
X_06567_ datapath.ru.latched_instruction\[18\] _01496_ vssd1 vssd1 vccd1 vccd1 _01497_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12376__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08306_ datapath.rf.registers\[28\]\[1\] net990 _01776_ net974 _01731_ vssd1 vssd1
+ vccd1 vccd1 _03233_ sky130_fd_sc_hd__a32o_1
XANTENNA__08989__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ net386 _04211_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o21ai_1
X_06498_ datapath.PC\[17\] vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08237_ datapath.rf.registers\[1\]\[2\] net977 net973 net998 vssd1 vssd1 vccd1 vccd1
+ _03164_ sky130_fd_sc_hd__o211a_1
XANTENNA__07661__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08168_ datapath.rf.registers\[18\]\[3\] _01741_ net972 vssd1 vssd1 vccd1 vccd1 _03095_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ datapath.rf.registers\[25\]\[26\] net797 net771 datapath.rf.registers\[30\]\[26\]
+ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08099_ datapath.rf.registers\[9\]\[4\] net885 net869 datapath.rf.registers\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10130_ net203 _05056_ net1309 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a21o_1
XANTENNA__07964__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10061_ datapath.PC\[19\] net1269 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__or2_1
XANTENNA__07716__A2 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10181__C1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_54_clk _00707_ net1178 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09469__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13751_ clknet_leaf_44_clk _00638_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11276__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ net294 net1707 net587 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_82_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
X_14536__1323 vssd1 vssd1 vccd1 vccd1 _14536__1323/HI net1323 sky130_fd_sc_hd__conb_1
XANTENNA__08049__B net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ net298 net1663 net570 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__mux2_1
X_13682_ clknet_leaf_110_clk _00617_ net1103 vssd1 vssd1 vccd1 vccd1 columns.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894_ net292 net2270 net594 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__mux2_1
X_12633_ _05666_ _05671_ net577 vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__or3_1
XFILLER_0_156_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12286__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ net174 net2034 net450 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07101__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14303_ clknet_leaf_37_clk _01190_ net1150 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11515_ screen.register.currentXbus\[20\] net1015 _05981_ _05983_ vssd1 vssd1 vccd1
+ vccd1 _05984_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12495_ net192 net2474 net457 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__mux2_1
X_14234_ clknet_leaf_23_clk _01121_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11446_ _05294_ net1014 _05916_ net1012 _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14165_ clknet_leaf_28_clk _01052_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11377_ _02875_ net714 vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13116_ clknet_leaf_53_clk _00108_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ datapath.i_ack mmio.WEN2 _01583_ _01599_ vssd1 vssd1 vccd1 vccd1 _05254_
+ sky130_fd_sc_hd__and4bb_1
X_14096_ clknet_leaf_4_clk _00983_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08231__C _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13047_ clknet_leaf_44_clk _00039_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ net508 net360 _04203_ net361 vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__o211a_1
XANTENNA__07168__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A2 _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
Xfanout1251 net1252 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__clkbuf_4
Xfanout1262 net1273 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__clkbuf_2
Xfanout1273 _00004_ vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06915__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1284 screen.counter.ct\[17\] vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__clkbuf_2
Xfanout1295 screen.counter.ct\[5\] vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_2
XANTENNA__09343__B _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13949_ clknet_leaf_33_clk _00836_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_73_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
X_07470_ datapath.rf.registers\[22\]\[18\] net752 net746 datapath.rf.registers\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
XANTENNA__07340__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _03981_ _04066_ net367 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09071_ _03988_ _03994_ _03505_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__o21a_1
XANTENNA__12924__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ net696 _02946_ _02948_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_116_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold701 datapath.rf.registers\[18\]\[17\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 screen.controlBus\[3\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold723 datapath.rf.registers\[5\]\[20\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold734 datapath.rf.registers\[14\]\[7\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 datapath.rf.registers\[21\]\[5\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 datapath.rf.registers\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 datapath.rf.registers\[28\]\[7\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 net40 vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _01715_ _04558_ _04560_ _04899_ net1053 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o311a_1
Xhold789 datapath.rf.registers\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09148__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ net330 _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__nand2_1
XANTENNA__07159__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _03776_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout569_A _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ datapath.rf.registers\[22\]\[11\] net952 net936 datapath.rf.registers\[21\]\[11\]
+ _02724_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08371__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08786_ net529 net359 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__or2_1
XANTENNA__11258__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ datapath.rf.registers\[14\]\[12\] net799 net722 datapath.rf.registers\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout736_A _01777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07668_ datapath.rf.registers\[26\]\[14\] net940 net904 datapath.rf.registers\[24\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09407_ net634 _04321_ _04331_ net612 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06619_ _01420_ _01512_ _01520_ _01526_ _01548_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__a2111o_1
X_07599_ _02522_ _02524_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__nor2_2
X_09338_ net397 _04171_ _04264_ net402 vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a211o_1
XANTENNA__10769__A1 _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12834__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _03122_ _03494_ net680 _03127_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ net21 net1045 net1034 mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1
+ vccd1 _00314_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ net2600 net263 net480 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11231_ net1427 net146 _05840_ _04878_ vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__a22o_1
XANTENNA__07398__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _05808_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__or2_1
XANTENNA__09139__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _05039_ net200 _04792_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__or3b_1
X_11093_ _05722_ net1013 _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__or3_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _03581_ _04970_ net1054 vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__a21o_1
Xhold50 datapath.multiplication_module.multiplier_i\[2\] vssd1 vssd1 vccd1 vccd1 net1416
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 net63 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 screen.controlBus\[25\] vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 keypad.decode.sticky_n\[4\] vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 screen.controlBus\[24\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ clknet_leaf_17_clk _00690_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11995_ datapath.mulitply_result\[3\] datapath.multiplication_module.multiplicand_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_55_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
X_13734_ clknet_leaf_111_clk _00621_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10946_ net232 net2578 net592 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_11_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07322__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13665_ clknet_leaf_57_clk _00603_ net1258 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10877_ net233 net2371 net600 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ net1629 net246 net441 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ clknet_leaf_80_clk screen.register.controlFill net1233 vssd1 vssd1 vccd1
+ vccd1 screen.register.cFill1 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08226__C _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12547_ net258 net2403 net448 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__mux2_1
XANTENNA__12744__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ net272 net1997 net457 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _01845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09378__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ clknet_leaf_2_clk _01104_ net1075 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11429_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_20_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07389__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07928__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ clknet_leaf_14_clk _01035_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06970_ datapath.rf.registers\[3\]\[30\] net965 net933 datapath.rf.registers\[23\]\[30\]
+ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a221o_1
X_14079_ clknet_leaf_38_clk _00966_ net1151 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06978__A _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1076 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_2
X_08640_ datapath.i_ack datapath.pc_module.i_ack2 vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__and2b_1
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07561__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ net1003 _03496_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__or2_1
XANTENNA__12919__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07522_ datapath.rf.registers\[11\]\[17\] net774 net734 datapath.rf.registers\[12\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a22o_1
XANTENNA__07313__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ datapath.rf.registers\[11\]\[19\] net970 net938 datapath.rf.registers\[21\]\[19\]
+ _02371_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07384_ datapath.rf.registers\[23\]\[20\] net788 net721 datapath.rf.registers\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09123_ _02787_ _03321_ _04048_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08813__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12654__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ net519 net518 _03545_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__mux2_1
XANTENNA__11778__B _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08005_ _02928_ _02929_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nor2_2
XANTENNA__09369__A1 _02997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 datapath.rf.registers\[20\]\[24\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 datapath.rf.registers\[19\]\[13\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 columns.count\[3\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07919__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14535__1322 vssd1 vssd1 vccd1 vccd1 _14535__1322/HI net1322 sky130_fd_sc_hd__conb_1
Xhold553 datapath.rf.registers\[16\]\[13\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 datapath.rf.registers\[14\]\[14\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 datapath.rf.registers\[26\]\[10\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 datapath.rf.registers\[14\]\[24\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 datapath.rf.registers\[14\]\[20\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10902__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _04849_ _04854_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__or2_1
XANTENNA__07483__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ _03462_ _03481_ net411 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__mux2_1
X_09887_ _04812_ _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 screen.register.currentYbus\[6\] vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 datapath.rf.registers\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 mmio.memload_or_instruction\[7\] vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ net362 _03707_ _03708_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1253 datapath.rf.registers\[30\]\[16\] vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 screen.register.currentYbus\[24\] vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 screen.register.currentXbus\[30\] vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ _01717_ _03695_ net493 vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a21o_1
XANTENNA__12829__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_10800_ datapath.mulitply_result\[11\] net426 net658 vssd1 vssd1 vccd1 vccd1 _05633_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _05604_ net175 _06192_ net177 vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10731_ _01651_ _01668_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__nand2_2
XFILLER_0_137_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ clknet_leaf_81_clk _00406_ net1240 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10662_ _05514_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ net164 net2362 net469 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ clknet_leaf_90_clk keypad.decode.sticky_n\[3\] net1210 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12564__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ net1411 net509 net350 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[5\]
+ sky130_fd_sc_hd__mux2_1
X_12332_ net2426 net184 net478 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XANTENNA__07083__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ net186 net2478 net485 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__mux2_1
X_14002_ clknet_leaf_34_clk _00889_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11214_ net1458 net145 net138 _05145_ vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__a22o_1
X_12194_ columns.count\[9\] _06438_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__xnor2_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_11145_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__inv_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__07791__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ net1023 _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nor2_1
XANTENNA__10127__C1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _04946_ _04953_ _04944_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__a21o_1
XANTENNA__07543__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11890__A2 _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11978_ net165 net2246 net580 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
XANTENNA__08518__A _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[2\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[2\] sky130_fd_sc_hd__dfrtp_1
X_10929_ net291 net2460 net591 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10486__C net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ clknet_leaf_100_clk _00586_ net1224 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13579_ clknet_leaf_89_clk _00529_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12474__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07074__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout307 _05860_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
X_09810_ datapath.PC\[1\] _03210_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__nand2_1
Xfanout318 net320 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
Xfanout329 net331 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
XANTENNA__07782__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09084__A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ datapath.PC\[26\] net628 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__xnor2_1
X_06953_ datapath.rf.registers\[7\]\[30\] net825 net806 datapath.rf.registers\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a22o_1
XANTENNA__06532__C_N mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ net331 _04425_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__nand2_1
X_06884_ datapath.rf.registers\[7\]\[31\] net957 net953 datapath.rf.registers\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a22o_1
XANTENNA__07534__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ net337 _03528_ net316 vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06888__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12649__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout267_A _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _03479_ _03480_ net409 vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ _02613_ _03409_ _03410_ _02611_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout434_A _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1176_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ datapath.rf.registers\[18\]\[19\] net790 net746 datapath.rf.registers\[21\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12384__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A _05668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ datapath.rf.registers\[16\]\[21\] net962 net910 datapath.rf.registers\[30\]\[21\]
+ _02293_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08798__C1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ net329 _04031_ _04032_ net380 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07298_ datapath.rf.registers\[31\]\[22\] net819 net761 datapath.rf.registers\[19\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09037_ net367 _03847_ _03846_ net374 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold350 datapath.rf.registers\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 datapath.rf.registers\[5\]\[8\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold372 datapath.rf.registers\[6\]\[9\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 datapath.rf.registers\[15\]\[20\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 datapath.rf.registers\[8\]\[24\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08610__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 _01737_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
Xfanout841 _01720_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_4
Xfanout852 net855 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_4
X_09939_ net206 _04864_ _04865_ net1312 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_144_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout863 _01851_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
Xfanout885 _01841_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_2
XANTENNA__08317__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
Xfanout896 net899 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_4
X_12950_ net229 net2390 net543 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__mux2_1
XANTENNA__07525__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11321__A1 _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 datapath.rf.registers\[13\]\[22\] vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 datapath.rf.registers\[16\]\[21\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net1439 _05886_ net157 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
Xhold1072 datapath.rf.registers\[29\]\[5\] vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 datapath.rf.registers\[18\]\[1\] vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ net238 net1668 net552 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
Xhold1094 datapath.rf.registers\[28\]\[3\] vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12559__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ datapath.PC\[19\] net304 _06229_ _06231_ vssd1 vssd1 vccd1 vccd1 _00463_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__B _05333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ net1362 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_11763_ _06179_ net1278 net302 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13502_ clknet_leaf_78_clk _00452_ net1246 vssd1 vssd1 vccd1 vccd1 datapath.PC\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_10714_ datapath.mulitply_result\[29\] net427 net661 vssd1 vssd1 vccd1 vccd1 _05561_
+ sky130_fd_sc_hd__a21o_1
X_14482_ clknet_leaf_35_clk _01369_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ screen.counter.currentCt\[19\] screen.counter.currentCt\[18\] _06134_ vssd1
+ vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13433_ clknet_leaf_79_clk _00389_ net1235 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ _01494_ net662 _05500_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12294__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10807__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__B2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ clknet_leaf_71_clk _00349_ net1230 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_10576_ net1388 _03060_ net347 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12315_ net1583 net263 net476 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
X_13295_ clknet_leaf_77_clk _00285_ net1247 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ net262 net2576 net484 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12177_ _06429_ _06430_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__nor2_1
XANTENNA__07764__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _05700_ _05775_ _05776_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__or4_1
XANTENNA__07417__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11059_ net1022 _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nor2_4
XANTENNA__07516__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12469__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09269__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14534__1321 vssd1 vssd1 vccd1 vccd1 _14534__1321/HI net1321 sky130_fd_sc_hd__conb_1
XFILLER_0_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ datapath.rf.registers\[26\]\[1\] net943 net913 datapath.rf.registers\[18\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07295__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07221_ net648 net530 net626 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07047__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ datapath.rf.registers\[0\]\[26\] net692 _02066_ _02078_ vssd1 vssd1 vccd1
+ vccd1 _02079_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_95_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09992__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12932__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ datapath.rf.registers\[9\]\[27\] net780 net768 datapath.rf.registers\[3\]\[27\]
+ _02009_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_8_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout126 _06265_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
XANTENNA__07755__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__B _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 net138 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 _05839_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_4
Xfanout159 _05261_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_07985_ datapath.rf.registers\[20\]\[7\] net804 net786 datapath.rf.registers\[23\]\[7\]
+ _02909_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a221o_1
X_09724_ _04649_ _04650_ _04639_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_126_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06936_ _01800_ _01860_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__nand2_1
XANTENNA__11303__B2 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ net614 _04574_ _04581_ _04580_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__o31a_1
XANTENNA__12379__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06867_ datapath.rf.registers\[6\]\[31\] net814 net806 datapath.rf.registers\[15\]\[31\]
+ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout551_A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08606_ net992 _03061_ net617 vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09586_ _04504_ _04509_ _04511_ _04512_ net657 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o41a_1
X_06798_ datapath.MemWrite _01723_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__or2_1
X_08537_ net514 net513 net407 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08468_ _03126_ _03389_ _03394_ _03124_ _03065_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_147_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ _02324_ net524 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__nor2_1
X_08399_ _02656_ _03325_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__or2_1
XANTENNA__11312__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _05344_ _00003_ vssd1 vssd1 vccd1 vccd1 keypad.decode.d1 sky130_fd_sc_hd__and2_1
XFILLER_0_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09432__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10042__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ screen.controlBus\[29\] screen.controlBus\[28\] screen.controlBus\[31\] screen.controlBus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12842__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12100_ datapath.mulitply_result\[20\] datapath.multiplication_module.multiplicand_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ clknet_leaf_39_clk _00072_ net1153 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10292_ net398 _04369_ _05217_ net339 vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12031_ _06306_ _06307_ _06305_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_57_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold180 datapath.rf.registers\[12\]\[1\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 datapath.rf.registers\[4\]\[24\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08340__B _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout660 net662 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11982__A datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout671 net672 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout682 net683 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout693 _01829_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_8
X_13982_ clknet_leaf_52_clk _00869_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09452__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ net298 net1572 net541 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__mux2_1
XANTENNA__12289__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06721__A1 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12864_ net630 _05575_ _06450_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__or3_4
X_11815_ net833 _03977_ net303 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_96_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12795_ net173 net2103 net564 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__mux2_1
XANTENNA__10110__B _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11746_ _06085_ _06168_ _06167_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__o21ai_1
X_14534_ net1321 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XANTENNA__07277__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13603__RESET_B net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10281__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11677_ _06126_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__inv_2
X_14465_ clknet_leaf_45_clk _01352_ net1186 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07029__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13416_ clknet_leaf_87_clk _00372_ net1220 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10628_ net1277 datapath.PC\[10\] _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__and3_1
X_14396_ clknet_leaf_57_clk _01283_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13347_ clknet_leaf_99_clk _00332_ net1227 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11230__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10559_ _05418_ _05460_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__nand2_1
XANTENNA__12752__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13278_ clknet_leaf_92_clk _00268_ net1204 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12229_ net191 net1986 net576 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__mux2_1
XANTENNA__07737__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06689__C _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07770_ net696 _02687_ _02696_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_108_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06721_ mmio.memload_or_instruction\[24\] net1059 net1005 datapath.ru.latched_instruction\[24\]
+ net1038 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09440_ _03684_ _04366_ net331 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__mux2_1
X_06652_ _01457_ net1029 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_88_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ _04296_ _04297_ net391 vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a21oi_1
X_06583_ net1307 net1303 mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ _01513_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12927__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _03203_ _03205_ _03244_ net651 _03245_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a221o_1
XANTENNA__07268__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08253_ net504 net505 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout132_A _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07204_ datapath.rf.registers\[19\]\[24\] net761 net728 datapath.rf.registers\[2\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08184_ datapath.rf.registers\[5\]\[3\] net783 _03093_ _03095_ _03101_ vssd1 vssd1
+ vccd1 vccd1 _03111_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11221__B1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07135_ datapath.rf.registers\[30\]\[26\] net910 net865 datapath.rf.registers\[13\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a22o_1
XANTENNA__12662__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07976__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09537__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__B _04383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ net533 _01972_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11259__A1_N net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A _05668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ datapath.rf.registers\[23\]\[7\] net932 net884 datapath.rf.registers\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__a22o_1
XANTENNA__10910__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09707_ _02258_ _02259_ _03704_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__or3_1
X_06919_ _01837_ _01840_ _01842_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__or4_1
XANTENNA__11827__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout933_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07899_ datapath.rf.registers\[23\]\[9\] net787 _02820_ _02825_ vssd1 vssd1 vccd1
+ vccd1 _02826_ sky130_fd_sc_hd__a211o_1
XANTENNA__08153__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _01996_ _03433_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__xnor2_1
X_09569_ _04477_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__nor2_1
XANTENNA__12837__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _05722_ _05791_ _05682_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ net1679 net257 net444 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__mux2_1
XANTENNA__07259__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09653__B1 _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__A _01682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ screen.register.currentXbus\[29\] _05700_ _05998_ vssd1 vssd1 vccd1 vccd1
+ _05999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08335__B _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14250_ clknet_leaf_11_clk _01137_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11462_ screen.register.currentYbus\[17\] _05775_ _05933_ vssd1 vssd1 vccd1 vccd1
+ _05934_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ clknet_leaf_8_clk _00193_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10015__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ datapath.multiplication_module.mul_prev _01636_ vssd1 vssd1 vccd1 vccd1 _05333_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11212__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ clknet_leaf_108_clk _01068_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11393_ _02499_ net668 vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and2_1
XANTENNA__12572__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07967__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ clknet_leaf_30_clk _00124_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10344_ net1296 net1295 vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_72_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ clknet_leaf_20_clk _00055_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10275_ net400 _04101_ _05200_ net340 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a211o_1
X_14533__1320 vssd1 vssd1 vccd1 vccd1 _14533__1320/HI net1320 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_72_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ datapath.mulitply_result\[6\] datapath.multiplication_module.multiplicand_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__or2_1
Xfanout490 _03625_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11279__B1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ clknet_leaf_0_clk _00852_ net1066 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08144__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ net1654 net244 net546 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XANTENNA__07498__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_13_clk _00783_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08229__C net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12747__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ net246 net1983 net554 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12778_ net259 net2227 net561 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14517_ net1308 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11729_ _06077_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14448_ clknet_leaf_4_clk _01335_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07670__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11203__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12482__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold905 datapath.rf.registers\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ clknet_leaf_56_clk _01266_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold916 datapath.rf.registers\[7\]\[21\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold927 datapath.rf.registers\[21\]\[6\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 datapath.rf.registers\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 datapath.rf.registers\[3\]\[20\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
X_08940_ net642 _03833_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08871_ _03448_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07822_ datapath.rf.registers\[4\]\[10\] net928 net864 datapath.rf.registers\[13\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10730__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ datapath.rf.registers\[22\]\[12\] net952 net856 datapath.rf.registers\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
X_06704_ _01627_ _01631_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__nand2_2
X_07684_ _02588_ _02609_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__or2_1
XANTENNA__07489__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09423_ net403 _03954_ _04349_ net336 vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__o211ai_2
X_06635_ mmio.memload_or_instruction\[8\] mmio.memload_or_instruction\[10\] mmio.memload_or_instruction\[9\]
+ mmio.memload_or_instruction\[7\] vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__and4bb_1
XANTENNA__12657__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ _03063_ _03494_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a21o_1
X_06566_ net1306 net1302 mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ _01496_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_23_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06655__S net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ datapath.rf.registers\[4\]\[1\] net812 _03229_ _03230_ _03231_ vssd1 vssd1
+ vccd1 vccd1 _03232_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ _02763_ net354 _04097_ net390 vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06497_ datapath.PC\[16\] vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout514_A _02812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ _03160_ _03161_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07661__A2 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08167_ datapath.rf.registers\[20\]\[3\] net987 _01734_ vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12392__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ datapath.rf.registers\[15\]\[26\] net806 net800 datapath.rf.registers\[14\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__a22o_1
XANTENNA__07413__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ datapath.rf.registers\[19\]\[4\] net945 net849 datapath.rf.registers\[1\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a22o_1
X_07049_ datapath.rf.registers\[8\]\[28\] net926 net901 datapath.rf.registers\[20\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_54_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__inv_2
XANTENNA__08374__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09433__C _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _05590_ net1592 net589 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__mux2_1
X_13750_ clknet_leaf_25_clk _00637_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ net290 net1631 net570 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__mux2_1
X_10893_ net297 net1844 net595 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__mux2_1
X_13681_ clknet_leaf_110_clk _00616_ net1104 vssd1 vssd1 vccd1 vccd1 columns.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12632_ net2212 net164 net441 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11433__B1 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12563_ net184 net1926 net449 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__mux2_1
XANTENNA__10787__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11514_ screen.register.currentXbus\[28\] net1013 _05982_ vssd1 vssd1 vccd1 vccd1
+ _05983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14302_ clknet_leaf_50_clk _01189_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07652__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12494_ net199 net2229 net458 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11445_ _05681_ _05741_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06860__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14233_ clknet_leaf_47_clk _01120_ net1265 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14164_ clknet_leaf_116_clk _01051_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11376_ screen.register.currentYbus\[7\] net132 _05873_ net161 vssd1 vssd1 vccd1
+ vccd1 _00365_ sky130_fd_sc_hd__a22o_1
XANTENNA__07404__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__A3 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ _01434_ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or2_1
XANTENNA__06612__B1 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13115_ clknet_leaf_55_clk _00107_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14095_ clknet_leaf_6_clk _00982_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13046_ clknet_leaf_26_clk _00038_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10258_ _03252_ _03386_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08365__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1230 net1255 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_2
X_10189_ net1276 _04047_ net540 vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__mux2_1
Xfanout1263 net1267 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_4
Xfanout1274 datapath.PC\[24\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_2
Xfanout1285 screen.counter.ct\[16\] vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__clkbuf_2
Xfanout1296 screen.counter.ct\[4\] vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_2
XANTENNA__08117__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10489__C net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ clknet_leaf_56_clk _00835_ net1256 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ clknet_leaf_44_clk _00766_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07891__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09070_ _02657_ net687 _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07643__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08021_ datapath.rf.registers\[22\]\[6\] net952 net896 datapath.rf.registers\[6\]\[6\]
+ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold702 datapath.rf.registers\[15\]\[17\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold713 datapath.rf.registers\[18\]\[9\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold724 datapath.rf.registers\[16\]\[23\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 datapath.rf.registers\[19\]\[17\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 datapath.rf.registers\[28\]\[14\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06603__B1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold757 datapath.rf.registers\[31\]\[8\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 net82 vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ datapath.PC\[27\] net539 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__or2_1
XANTENNA__12940__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold779 datapath.rf.registers\[10\]\[31\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08923_ net382 _03848_ _03849_ _03845_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08854_ net706 _03780_ net623 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10163__B1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ datapath.rf.registers\[31\]\[11\] net948 net908 datapath.rf.registers\[30\]\[11\]
+ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a221o_1
X_08785_ net497 net494 net531 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__a21o_1
XANTENNA__08108__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout464_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ datapath.rf.registers\[22\]\[12\] net751 net744 datapath.rf.registers\[21\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XANTENNA__09550__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12387__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ datapath.rf.registers\[27\]\[14\] net868 net848 datapath.rf.registers\[1\]\[14\]
+ _02589_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06618_ datapath.ru.latched_instruction\[24\] _01473_ _01496_ datapath.ru.latched_instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__a22o_1
X_09406_ net653 _04315_ _04329_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__or4_1
X_07598_ _02524_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__inv_2
XANTENNA__07882__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06549_ mmio.memload_or_instruction\[17\] net1058 vssd1 vssd1 vccd1 vccd1 _01479_
+ sky130_fd_sc_hd__and2_1
X_09337_ net387 _04014_ _04161_ net392 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10769__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07095__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ net506 _03121_ net684 vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__o21a_1
XANTENNA__07634__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ datapath.rf.registers\[0\]\[2\] net690 _03133_ _03145_ vssd1 vssd1 vccd1
+ vccd1 _03146_ sky130_fd_sc_hd__o22a_4
X_09199_ _02974_ net686 _04124_ net317 _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11230_ net1418 net146 net139 _04888_ vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09387__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08332__C _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _05705_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__nor2_1
XANTENNA__12850__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _04790_ _04791_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__nor2_1
X_11092_ _05731_ net1021 vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__nor2_4
X_10043_ net1275 _03580_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nand2_1
XANTENNA__08898__A1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 net113 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 datapath.multiplication_module.multiplier_i\[11\] vssd1 vssd1 vccd1 vccd1
+ net1417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 net59 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 screen.controlBus\[20\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 net52 vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 net50 vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_11_clk _00689_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11994_ net2277 net326 net322 _06279_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13733_ clknet_leaf_94_clk _00620_ net1206 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12297__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ net227 net1964 net590 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13664_ clknet_leaf_57_clk _00602_ net1261 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10876_ net228 net2163 net598 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__mux2_1
XANTENNA__07873__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12615_ net1717 net249 net440 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ clknet_leaf_81_clk net1385 net1238 vssd1 vssd1 vccd1 vccd1 screen.register.xFill3
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ net262 net2018 net448 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07625__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12477_ net273 net1903 net459 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
XANTENNA_4 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output93_A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ clknet_leaf_15_clk _01103_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09378__A2 _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11428_ net1011 _05712_ _05898_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08586__B1 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ clknet_leaf_106_clk _01034_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11359_ keypad.alpha _05864_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12760__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ clknet_leaf_51_clk _00965_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13029_ clknet_leaf_93_clk _00021_ net1203 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10145__B1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 _01455_ vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1084 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1125 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_2
X_08570_ net1003 _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__nor2_2
X_07521_ _02441_ _02443_ _02445_ _02447_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__or4_1
XANTENNA__11405__A _02234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07452_ datapath.rf.registers\[8\]\[19\] net926 net893 datapath.rf.registers\[14\]\[19\]
+ _02378_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07383_ datapath.rf.registers\[15\]\[20\] net807 net764 datapath.rf.registers\[17\]\[20\]
+ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a221o_1
XANTENNA__12935__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09122_ _03404_ _04048_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07077__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09053_ net363 _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout212_A _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08004_ net512 _02927_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XANTENNA__08433__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold510 datapath.rf.registers\[18\]\[10\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 datapath.rf.registers\[31\]\[11\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 datapath.rf.registers\[16\]\[8\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold543 datapath.rf.registers\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 datapath.rf.registers\[14\]\[11\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12670__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold565 datapath.rf.registers\[21\]\[17\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1121_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 datapath.rf.registers\[6\]\[24\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 datapath.rf.registers\[8\]\[11\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11794__B _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 datapath.rf.registers\[28\]\[19\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ datapath.PC\[29\] _01715_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout581_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ _03418_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__xnor2_1
X_09886_ _04700_ _04759_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__xor2_1
Xhold1210 datapath.rf.registers\[2\]\[11\] vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 datapath.rf.registers\[27\]\[6\] vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 datapath.rf.registers\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 datapath.rf.registers\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net381 _03623_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nor2_1
Xhold1254 screen.register.currentYbus\[14\] vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 datapath.rf.registers\[16\]\[20\] vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 datapath.rf.registers\[8\]\[0\] vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ _03669_ _03685_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_49_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _02640_ _02641_ _02645_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_49_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ net499 net620 net488 vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10730_ net163 net2547 net607 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__mux2_1
XANTENNA__08327__C _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ datapath.PC\[21\] _05503_ datapath.PC\[22\] vssd1 vssd1 vccd1 vccd1 _05515_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__12845__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ net167 net2569 net470 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_149_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13380_ clknet_leaf_90_clk keypad.decode.sticky_n\[2\] net1210 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10592_ net1562 net507 net350 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[4\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07607__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ net1769 net188 net478 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XANTENNA__08343__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12262_ net188 net2477 net486 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__mux2_1
XANTENNA__13699__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ net1431 net144 net138 _05165_ vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__a22o_1
X_14001_ clknet_leaf_27_clk _00888_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08032__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ _05851_ _06440_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__nor2_1
XANTENNA__12580__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_120_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11144_ _05738_ _05793_ _05739_ _05790_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or4b_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11075_ net1298 _05718_ net1297 vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__or3b_2
X_10026_ net201 _04952_ net1312 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11875__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__B net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08099__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11977_ net167 net2247 net580 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ clknet_leaf_96_clk datapath.multiplication_module.multiplier_i_n\[1\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[1\] sky130_fd_sc_hd__dfrtp_1
X_10928_ net299 net2360 net591 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__mux2_1
XANTENNA__07846__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12755__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ clknet_leaf_69_clk _00585_ net1224 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09048__A1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10859_ net300 net2484 net599 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__mux2_1
XANTENNA__09048__B2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07059__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13578_ clknet_leaf_89_clk _00528_ net1213 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10602__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ net2245 net188 net453 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__mux2_1
XANTENNA__08271__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08559__A0 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12490__S net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold33_A datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 _05860_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
X_09740_ _03637_ _04585_ _04608_ _04610_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a31o_1
X_06952_ datapath.rf.registers\[13\]\[30\] net793 net739 datapath.rf.registers\[8\]\[30\]
+ _01878_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a221o_1
.ends

