* NGSPICE file created from team_05.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt team_05 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
X_05903_ net489 _02538_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__or2_1
X_06883_ top.compVal\[12\] top.findLeastValue.val1\[12\] net154 vssd1 vssd1 vccd1
+ vccd1 _03647_ sky130_fd_sc_hd__mux2_1
X_09671_ net754 net589 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__and2_1
X_08622_ top.cb_syn.end_cnt\[3\] _04841_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__or2_1
XANTENNA__05545__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05834_ top.hTree.state\[2\] _02841_ _02853_ _02854_ vssd1 vssd1 vccd1 vccd1 _02856_
+ sky130_fd_sc_hd__and4_1
X_08553_ net1327 top.cb_syn.char_path_n\[6\] net238 vssd1 vssd1 vccd1 vccd1 _01489_
+ sky130_fd_sc_hd__mux2_1
X_05765_ top.compVal\[43\] net162 _02806_ top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XANTENNA__09304__S top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ net1367 top.cb_syn.char_path_n\[75\] net244 vssd1 vssd1 vccd1 vccd1 _01558_
+ sky130_fd_sc_hd__mux2_1
X_07504_ _02989_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_85_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout162_A _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05696_ top.cb_syn.char_path\[5\] net549 net541 top.cb_syn.char_path\[69\] vssd1
+ vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a22o_1
XANTENNA__06987__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07435_ net344 top.dut.bits_in_buf_next\[2\] vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout427_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07366_ _03814_ _03850_ _03812_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06317_ net406 _03089_ _03185_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__nand3_1
X_09105_ net481 _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__nor2_1
X_07297_ _03743_ _03747_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__nand3_1
X_06248_ net482 net406 _03090_ _02503_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a211o_1
X_09036_ top.WB.CPU_DAT_O\[14\] net1286 net315 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout796_A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold340 top.cb_syn.char_path\[58\] vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 top.cb_syn.char_path\[99\] vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ net445 _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__nand2_1
Xhold362 top.hTree.tree_reg\[34\] vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 top.cb_syn.char_path\[33\] vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 top.hTree.nulls\[55\] vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 top.histogram.sram_out\[3\] vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
X_09938_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__and2_1
XANTENNA__08970__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout842 net843 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07773__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout820 net826 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_2
Xfanout831 net834 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_2
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_2
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_2
X_09869_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__and2_1
XANTENNA__06130__C net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ net931 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
X_11831_ clknet_leaf_67_clk _02364_ _01203_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07289__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ clknet_leaf_74_clk net1276 vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10713_ clknet_leaf_45_clk _01344_ _00103_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_11693_ clknet_leaf_103_clk _02243_ _01083_ vssd1 vssd1 vccd1 vccd1 top.compVal\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_10644_ clknet_leaf_75_clk _01275_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10575_ net785 net620 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__and2_1
XANTENNA__08636__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ clknet_leaf_62_clk _01692_ _00517_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[73\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07764__B2 top.findLeastValue.sum\[45\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__A0 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05775__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ clknet_leaf_47_clk _01623_ _00448_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10009_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05550_ net1796 net166 _02631_ net213 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05481_ net29 net415 net364 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 _02377_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08229__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07220_ top.findLeastValue.val2\[40\] top.findLeastValue.val1\[40\] vssd1 vssd1 vccd1
+ vccd1 _03896_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07151_ top.findLeastValue.val2\[1\] top.findLeastValue.val1\[1\] vssd1 vssd1 vccd1
+ vccd1 _03827_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_30_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06102_ top.cb_syn.count\[4\] _03000_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07082_ _03743_ _03747_ _03744_ _03742_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__a211oi_1
X_06033_ _02928_ _02937_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__nor2_1
XANTENNA__07755__A1 top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout127 _03611_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_4
Xfanout116 _03661_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08952__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05766__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07984_ net436 net1538 net250 top.findLeastValue.sum\[1\] _04513_ vssd1 vssd1 vccd1
+ vccd1 _01790_ sky130_fd_sc_hd__a221o_1
X_09723_ net867 net702 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__and2_1
X_06935_ top.findLeastValue.val1\[22\] net139 net116 net1784 vssd1 vssd1 vccd1 vccd1
+ _01983_ sky130_fd_sc_hd__o22a_1
X_09654_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout377_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ top.findLeastValue.val2\[21\] net132 net117 _03638_ vssd1 vssd1 vccd1 vccd1
+ _02029_ sky130_fd_sc_hd__o22a_1
X_08605_ _02541_ _04820_ _04822_ _04824_ top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1
+ vccd1 _04825_ sky130_fd_sc_hd__o221a_1
X_05817_ net442 net431 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09585_ net745 net580 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__and2_1
X_06797_ _02421_ top.findLeastValue.val2\[31\] _03572_ vssd1 vssd1 vccd1 vccd1 _03595_
+ sky130_fd_sc_hd__a21oi_1
X_08536_ net1056 top.cb_syn.char_path_n\[23\] net236 vssd1 vssd1 vccd1 vccd1 _01506_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05748_ top.findLeastValue.histo_index\[7\] _02789_ _02791_ _02500_ vssd1 vssd1 vccd1
+ vccd1 _02792_ sky130_fd_sc_hd__o211a_1
X_08467_ net1082 top.cb_syn.char_path_n\[92\] net236 vssd1 vssd1 vccd1 vccd1 _01575_
+ sky130_fd_sc_hd__mux2_1
X_05679_ top.cb_syn.char_path\[40\] net529 net312 top.cb_syn.char_path\[104\] vssd1
+ vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ top.cb_syn.char_path_n\[5\] net197 _04761_ vssd1 vssd1 vccd1 vccd1 _01624_
+ sky130_fd_sc_hd__o21a_1
X_07418_ _02521_ net125 net123 _04039_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07349_ _03859_ _03995_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10360_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__and2_1
XANTENNA__09717__B net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ net829 net664 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__and2_1
X_09019_ top.WB.CPU_DAT_O\[31\] net1306 net314 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
XANTENNA__07994__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 top.cb_syn.char_path\[51\] vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05737__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 top.cb_syn.char_path\[90\] vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 top.findLeastValue.histo_index\[1\] vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_2
Xfanout683 net689 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_2
Xfanout694 net700 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_1
Xfanout672 net680 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_1
Xfanout661 net670 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ clknet_leaf_82_clk _02347_ _01186_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
X_11745_ clknet_leaf_11_clk _02295_ _01135_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.zero_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07700__B _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11676_ clknet_leaf_87_clk _02226_ _01066_ vssd1 vssd1 vccd1 vccd1 top.compVal\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08226__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10627_ clknet_leaf_82_clk _01258_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10558_ net860 net695 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05996__A0 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__A1 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ net785 net620 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06720_ _02414_ top.findLeastValue.val2\[33\] vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06651_ _03447_ _03448_ _03446_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__or3b_1
X_05602_ top.histogram.sram_out\[21\] net359 net410 top.hTree.node_reg\[21\] vssd1
+ vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06582_ top.header_synthesis.count\[3\] _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _03382_
+ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_82_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09370_ top.hTree.nulls\[49\] net398 net228 vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08321_ top.cb_syn.char_path_n\[44\] net381 net338 top.cb_syn.char_path_n\[42\] net184
+ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__a221o_1
X_05533_ _02615_ _02617_ top.WB.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__or3b_1
X_08252_ top.cb_syn.char_path_n\[78\] net203 _04688_ vssd1 vssd1 vccd1 vccd1 _01697_
+ sky130_fd_sc_hd__o21a_1
X_05464_ net16 net414 net363 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 _02394_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07203_ _02462_ _02487_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08217__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ top.cb_syn.char_path_n\[113\] net378 net334 top.cb_syn.char_path_n\[111\]
+ net181 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_05395_ top.cw2\[0\] vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout125_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07425__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07134_ _03807_ _03809_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07520__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05987__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ top.findLeastValue.val2\[30\] top.findLeastValue.val1\[30\] vssd1 vssd1 vccd1
+ vccd1 _03741_ sky130_fd_sc_hd__xor2_1
X_06016_ top.sram_interface.init_counter\[5\] top.sram_interface.init_counter\[4\]
+ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout661_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ net477 _04498_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__or2_1
X_09706_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout759_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06918_ top.findLeastValue.val1\[39\] net137 net112 net1764 vssd1 vssd1 vccd1 vccd1
+ _02000_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07898_ net421 _04443_ _04444_ net263 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o211a_1
XANTENNA__09350__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__and2_1
X_06849_ top.compVal\[29\] top.findLeastValue.val1\[29\] net151 vssd1 vssd1 vccd1
+ vccd1 _03630_ sky130_fd_sc_hd__mux2_1
X_09568_ net773 net608 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__and2_1
X_08519_ net1319 top.cb_syn.char_path_n\[40\] net240 vssd1 vssd1 vccd1 vccd1 _01523_
+ sky130_fd_sc_hd__mux2_1
X_11530_ clknet_leaf_81_clk net1465 _00920_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09499_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_102_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ clknet_leaf_79_clk _02026_ _00851_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[18\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__05690__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11392_ clknet_leaf_13_clk _01957_ _00782_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10412_ net739 net574 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__and2_1
XANTENNA__06851__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05978__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__and2_1
XANTENNA__08392__A1 top.cb_syn.char_path_n\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout491 top.cb_syn.char_found vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_2
XANTENNA__06942__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout480 top.hTree.state\[0\] vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09341__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10402__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ clknet_leaf_46_clk _02278_ _01118_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ clknet_leaf_117_clk _02209_ _01049_ vssd1 vssd1 vccd1 vccd1 top.path\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05681__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07958__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08870_ top.translation.totalEn _05049_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__and2_1
X_07821_ top.hTree.tree_reg\[33\] top.findLeastValue.sum\[33\] net266 vssd1 vssd1
+ vccd1 vccd1 _04383_ sky130_fd_sc_hd__mux2_1
XANTENNA__07569__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ net472 _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nand2_1
XANTENNA__09332__B1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ top.hTree.tree_reg\[59\] top.findLeastValue.least1\[4\] net280 vssd1 vssd1
+ vccd1 vccd1 _04271_ sky130_fd_sc_hd__mux2_1
X_06703_ _03479_ _03500_ _03482_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06001__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ net966 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07894__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06634_ _02443_ top.findLeastValue.val1\[3\] top.findLeastValue.val1\[2\] _02444_
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__o22a_1
X_09353_ net1475 net225 net215 _04363_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ net1697 net197 _04714_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06565_ top.dut.out\[7\] top.dut.out\[6\] top.dut.out\[5\] top.dut.out\[4\] vssd1
+ vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__or4b_1
X_05516_ top.findLeastValue.wipe_the_char_1 _02576_ vssd1 vssd1 vccd1 vccd1 _02601_
+ sky130_fd_sc_hd__and2_1
X_06496_ top.histogram.total\[6\] _03325_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_
+ sky130_fd_sc_hd__and3_1
X_09284_ top.histogram.total\[20\] top.histogram.total\[21\] top.histogram.total\[22\]
+ top.histogram.total\[23\] net508 net506 vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__mux4_1
X_08235_ top.cb_syn.char_path_n\[87\] net377 net334 top.cb_syn.char_path_n\[85\] net180
+ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__a221o_1
X_05447_ top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__inv_2
XANTENNA__05672__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08166_ top.cb_syn.char_path_n\[121\] net194 _04645_ vssd1 vssd1 vccd1 vccd1 _01740_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09399__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05378_ top.findLeastValue.val1\[13\] vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__inv_2
X_07117_ top.findLeastValue.val2\[15\] top.findLeastValue.val1\[15\] vssd1 vssd1 vccd1
+ vccd1 _03793_ sky130_fd_sc_hd__nand2_1
X_08097_ top.cb_syn.num_lefts\[7\] _04589_ _04590_ _04598_ vssd1 vssd1 vccd1 vccd1
+ _01762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07048_ _03722_ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ top.WB.CPU_DAT_O\[21\] net1168 net365 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XANTENNA__06924__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ clknet_leaf_61_clk _01526_ _00351_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06137__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ clknet_leaf_31_clk _01464_ _00282_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11513_ clknet_leaf_117_clk _02078_ _00903_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05663__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ clknet_leaf_90_clk _02009_ _00834_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_11375_ clknet_leaf_13_clk _01940_ _00765_ vssd1 vssd1 vccd1 vccd1 top.cw1\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ net728 net563 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__and2_1
X_10257_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__and2_1
X_10188_ net800 net635 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__and2_1
XANTENNA__06915__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06350_ top.cb_syn.char_index\[0\] _02605_ _03217_ top.controller.state_reg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06300__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06281_ top.cb_syn.char_index\[3\] _03034_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__xnor2_1
X_05301_ top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__inv_2
XANTENNA__05654__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08020_ _02783_ _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 top.compVal\[45\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 top.hTree.node_reg\[47\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold725 top.findLeastValue.sum\[27\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 top.compVal\[8\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 top.cb_syn.char_path_n\[83\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold758 top.findLeastValue.sum\[17\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 top.compVal\[3\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net750 net585 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08922_ top.cb_syn.max_index\[5\] _05060_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout192_A _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _02550_ _02812_ _05037_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__a21oi_1
X_07804_ net435 net1594 net249 top.findLeastValue.sum\[37\] _04369_ vssd1 vssd1 vccd1
+ vccd1 _01826_ sky130_fd_sc_hd__a221o_1
X_08784_ top.path\[10\] top.path\[11\] net510 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__mux2_1
X_05996_ top.WB.CPU_DAT_O\[5\] net1052 net347 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
X_07735_ net473 _04310_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__or2_1
X_09405_ net999 _05283_ net229 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
X_07666_ top.hTree.tree_reg\[63\] net471 net282 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or3_1
XANTENNA__07351__A _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ net412 _02896_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06617_ top.findLeastValue.val1\[18\] top.compVal\[18\] vssd1 vssd1 vccd1 vccd1 _03415_
+ sky130_fd_sc_hd__and2b_1
X_09336_ net998 net221 net219 _04431_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__a22o_1
XANTENNA__09084__A2 top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06548_ _03325_ _03328_ _03330_ top.histogram.total\[8\] vssd1 vssd1 vccd1 vccd1
+ _03358_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09267_ net1684 _04046_ top.dut.bits_in_buf_next\[0\] _04098_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf_next\[0\] sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_23_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08218_ top.cb_syn.char_path_n\[95\] net190 _04671_ vssd1 vssd1 vccd1 vccd1 _01714_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06479_ net1155 net297 _03316_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ _05180_ _05181_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__nor2_1
X_08149_ top.cb_syn.cb_length\[0\] net172 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__xnor2_1
X_11160_ clknet_leaf_60_clk _01725_ _00550_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[106\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08910__A top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11091_ clknet_leaf_63_clk _01656_ _00481_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[37\]
+ sky130_fd_sc_hd__dfrtp_2
X_10111_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10042_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__and2_1
Xhold30 top.sram_interface.check vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 top.hTree.node_reg\[4\] vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 top.hTree.node_reg\[8\] vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 top.hTree.node_reg\[40\] vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 top.hTree.node_reg\[14\] vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 net57 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 top.sram_interface.word_cnt\[4\] vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10944_ clknet_leaf_36_clk _01509_ _00334_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10875_ clknet_leaf_23_clk _01460_ _00265_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05636__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_5 DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ clknet_leaf_100_clk _01992_ _00817_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[31\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11358_ clknet_leaf_94_clk _01923_ _00748_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_10309_ net839 net674 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__and2_1
X_11289_ clknet_leaf_24_clk _01854_ _00679_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05850_ net1761 _02869_ _02870_ _02871_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07870__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ top.cb_syn.char_path_n\[126\] top.cb_syn.char_path_n\[125\] top.cb_syn.curr_path\[127\]
+ top.cb_syn.char_path_n\[127\] net394 net292 vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__mux4_1
XANTENNA__05572__B2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05781_ net505 net402 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__nor2_1
XANTENNA__07849__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07451_ top.dut.out\[7\] net343 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__and2_1
X_06402_ top.hist_data_o\[16\] _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07382_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__nand2b_1
X_06333_ net458 _03190_ _03198_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__a211o_1
X_09121_ top.histogram.init_edge _02416_ _03244_ _05080_ vssd1 vssd1 vccd1 vccd1 _05133_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_20_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09052_ net412 _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05627__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06264_ _02605_ _03046_ _03135_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or3_1
Xhold511 net76 vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 _01833_ vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
X_08003_ top.findLeastValue.least2\[4\] top.findLeastValue.least1\[4\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
X_06195_ _02590_ _03052_ _03067_ _03068_ _02607_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout205_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold533 net86 vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 top.hTree.tree_reg\[28\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 net73 vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold588 top.cb_syn.char_path\[76\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 top.histogram.wr_r_en\[1\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 top.hist_data_o\[5\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 top.histogram.total\[27\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net771 net606 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__and2_1
Xhold599 top.cb_syn.curr_index\[5\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
X_09885_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__and2_1
X_08905_ net470 _02851_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nor2_1
X_08836_ _05024_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout839_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05979_ top.WB.CPU_DAT_O\[22\] net1296 net345 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
X_08767_ net425 _04954_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout741_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08698_ top.header_synthesis.count\[2\] top.header_synthesis.count\[1\] _04896_ vssd1
+ vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__and3_1
X_07718_ net449 net1066 _04257_ _04299_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__o22a_1
XANTENNA__07304__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ top.cb_syn.h_element\[55\] top.cb_syn.h_element\[46\] _04176_ vssd1 vssd1
+ vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ clknet_leaf_67_clk _01291_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_09319_ net992 net224 net216 _04499_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_114_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10591_ net799 net634 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__and2_1
XANTENNA__05618__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11212_ clknet_leaf_107_clk _01777_ _00602_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11143_ clknet_leaf_36_clk _01708_ _00533_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[89\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__clkbuf_4
X_11074_ clknet_leaf_53_clk _01639_ _00464_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
X_10025_ net833 net668 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__and2_1
XANTENNA__05554__B2 top.hTree.node_reg\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ clknet_leaf_61_clk _01492_ _00317_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10858_ clknet_leaf_10_clk _01452_ _00248_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.TRN_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_105_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10789_ clknet_leaf_117_clk _01395_ _00179_ vssd1 vssd1 vccd1 vccd1 top.path\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05609__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08559__A1 top.cb_syn.char_path_n\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07865__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout309 net312 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_4
X_06951_ top.findLeastValue.val1\[6\] net136 net113 net1793 vssd1 vssd1 vccd1 vccd1
+ _01967_ sky130_fd_sc_hd__o22a_1
X_05902_ _02882_ _02883_ top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 _02884_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__06990__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ net733 net568 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ _04839_ _04840_ net497 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__mux2_1
X_06882_ top.findLeastValue.val2\[13\] net130 net120 _03646_ vssd1 vssd1 vccd1 vccd1
+ _02021_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05833_ top.sram_interface.counter_HTREE\[1\] top.sram_interface.counter_HTREE\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__nand2_1
X_08552_ net1284 top.cb_syn.char_path_n\[7\] net240 vssd1 vssd1 vccd1 vccd1 _01490_
+ sky130_fd_sc_hd__mux2_1
X_05764_ top.compVal\[44\] net163 _02806_ top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 _02329_ sky130_fd_sc_hd__a22o_1
XANTENNA__09287__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ net1539 top.cb_syn.char_path_n\[76\] net245 vssd1 vssd1 vccd1 vccd1 _01559_
+ sky130_fd_sc_hd__mux2_1
X_07503_ _02990_ _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_85_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08590__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05695_ net1392 net170 _02752_ net209 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout155_A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07434_ _04044_ vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf_next\[2\] sky130_fd_sc_hd__inv_2
XFILLER_0_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07365_ top.findLeastValue.sum\[12\] net279 net272 _04007_ vssd1 vssd1 vccd1 vccd1
+ _01899_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout322_A _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06316_ net486 _03088_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__nand2_1
X_09104_ top.histogram.init_edge _05080_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__or2_2
XFILLER_0_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07296_ _03762_ _03957_ _03749_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a21o_1
XANTENNA__08798__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06247_ _03081_ _03118_ _02600_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__and3b_1
X_09035_ top.WB.CPU_DAT_O\[15\] net1134 net315 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold352 top.cb_syn.char_path\[124\] vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 top.cb_syn.char_path\[93\] vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ top.TRN_char_index\[1\] top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 _03053_
+ sky130_fd_sc_hd__or2_1
Xhold330 top.sram_interface.write_counter_FLV\[1\] vssd1 vssd1 vccd1 vccd1 net1281
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold385 top.cb_syn.char_path\[57\] vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 top.cb_syn.char_path\[71\] vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 net95 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 top.dut.out\[5\] vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
X_09937_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__and2_1
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
Xfanout832 net833 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout821 net822 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_2
Xfanout810 net812 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__buf_1
Xfanout854 net877 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_2
Xfanout865 net876 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_2
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_2
X_09868_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__and2_1
XANTENNA__06130__D net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09291__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__and2_1
X_08819_ net505 _05004_ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a21oi_1
X_11830_ clknet_leaf_67_clk _02363_ _01202_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11761_ clknet_leaf_45_clk _02300_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07289__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ clknet_leaf_46_clk _01343_ _00102_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_11692_ clknet_leaf_103_clk _02242_ _01082_ vssd1 vssd1 vccd1 vccd1 top.compVal\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_10643_ clknet_leaf_74_clk _01274_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10574_ net838 net673 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08636__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ clknet_leaf_61_clk _01691_ _00516_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[72\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05775__B2 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ clknet_leaf_48_clk _01622_ _00447_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09405__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ net840 net675 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05480_ net30 net413 net362 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 _02378_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08229__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06101_ _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__inv_2
X_07081_ _03753_ _03754_ _03755_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__or3_1
X_06032_ _02924_ _02926_ net1702 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout117 net122 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout128 net131 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_4
X_09722_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__and2_1
Xfanout139 _03508_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
XANTENNA__05766__B2 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ net419 _04511_ _04512_ net261 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o211a_1
XANTENNA__06963__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ top.findLeastValue.val1\[23\] net138 net115 net1776 vssd1 vssd1 vccd1 vccd1
+ _01984_ sky130_fd_sc_hd__o22a_1
X_09653_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__and2_1
X_06865_ top.compVal\[21\] top.findLeastValue.val1\[21\] net156 vssd1 vssd1 vccd1
+ vccd1 _03638_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ net496 _04823_ top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__a21o_1
X_05816_ top.hTree.write_HT_fin net417 _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__or3b_1
X_09584_ net797 net632 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ net1230 top.cb_syn.char_path_n\[24\] net235 vssd1 vssd1 vccd1 vccd1 _01507_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06796_ top.compVal\[16\] _02471_ _03561_ _03562_ vssd1 vssd1 vccd1 vccd1 _03594_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout537_A top.sram_interface.word_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05747_ _02789_ _02790_ _02785_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__o21a_1
X_08466_ net1292 top.cb_syn.char_path_n\[93\] net230 vssd1 vssd1 vccd1 vccd1 _01576_
+ sky130_fd_sc_hd__mux2_1
X_05678_ top.cb_syn.char_path\[8\] net547 net540 top.cb_syn.char_path\[72\] vssd1
+ vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout704_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ top.cb_syn.char_path_n\[6\] net375 net332 top.cb_syn.char_path_n\[4\] net178
+ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ top.findLeastValue.histo_index\[0\] top.findLeastValue.least1\[0\] net148
+ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _03859_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08640__B1 top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07279_ _03874_ _03888_ _03886_ _03883_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ net829 net664 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__and2_1
XANTENNA__09286__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ top.sram_interface.TRN_counter\[2\] _02914_ top.sram_interface.TRN_counter\[1\]
+ top.sram_interface.TRN_counter\[0\] vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__or4b_1
Xhold171 _01534_ vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 top.cb_syn.char_path\[35\] vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 top.cb_syn.char_path\[115\] vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05319__A top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 top.path\[112\] vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout651 net712 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_2
Xfanout640 net643 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_1
Xfanout684 net689 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_1
Xfanout673 net680 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06849__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 net670 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_2
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07903__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ clknet_leaf_65_clk _02346_ _01185_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11744_ clknet_leaf_6_clk _02294_ _01134_ vssd1 vssd1 vccd1 vccd1 top.histogram.init_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11675_ clknet_leaf_87_clk _02225_ _01065_ vssd1 vssd1 vccd1 vccd1 top.compVal\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_10626_ clknet_leaf_67_clk _01257_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05501__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ net860 net695 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10488_ net785 net620 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__and2_1
XANTENNA__07709__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05748__A1 top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06945__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ clknet_leaf_49_clk _01674_ _00499_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_06650_ _02436_ top.findLeastValue.val1\[10\] top.findLeastValue.val1\[9\] _02437_
+ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a22o_1
X_05601_ _02672_ _02673_ net467 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07370__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06581_ _02544_ _03380_ _03379_ _03375_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08320_ top.cb_syn.char_path_n\[44\] net202 _04722_ vssd1 vssd1 vccd1 vccd1 _01663_
+ sky130_fd_sc_hd__o21a_1
X_05532_ _02599_ _02614_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__nor2_1
X_08251_ top.cb_syn.char_path_n\[79\] net384 net339 top.cb_syn.char_path_n\[77\] net186
+ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05463_ net17 net414 net363 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 _02395_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_15_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05684__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ top.findLeastValue.val2\[35\] top.findLeastValue.val1\[35\] vssd1 vssd1 vccd1
+ vccd1 _03878_ sky130_fd_sc_hd__nor2_1
X_08182_ net1755 net199 _04653_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__o21a_1
X_05394_ top.cw2\[1\] vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07133_ top.findLeastValue.val2\[11\] top.findLeastValue.val1\[11\] vssd1 vssd1 vccd1
+ vccd1 _03809_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07520__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07064_ top.findLeastValue.val2\[31\] top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1
+ vccd1 _03740_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout118_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06015_ _02924_ _02927_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06936__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ top.findLeastValue.sum\[4\] _04498_ net391 vssd1 vssd1 vccd1 vccd1 _04499_
+ sky130_fd_sc_hd__mux2_1
X_09705_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__and2_1
X_06917_ top.findLeastValue.val1\[40\] net137 net112 top.compVal\[40\] vssd1 vssd1
+ vccd1 vccd1 _02001_ sky130_fd_sc_hd__o22a_1
X_09636_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07897_ net478 _04442_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout654_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06164__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06848_ top.findLeastValue.val2\[30\] net127 net118 _03629_ vssd1 vssd1 vccd1 vccd1
+ _02038_ sky130_fd_sc_hd__o22a_1
X_09567_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__and2_1
X_06779_ top.findLeastValue.val2\[23\] top.compVal\[23\] vssd1 vssd1 vccd1 vccd1 _03577_
+ sky130_fd_sc_hd__nand2b_1
X_08518_ net1357 top.cb_syn.char_path_n\[41\] net240 vssd1 vssd1 vccd1 vccd1 _01524_
+ sky130_fd_sc_hd__mux2_1
X_09498_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__and2_1
X_08449_ net1063 top.cb_syn.char_path_n\[110\] net244 vssd1 vssd1 vccd1 vccd1 _01593_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08861__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05675__B1 _02735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11460_ clknet_leaf_101_clk _02025_ _00850_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_11391_ clknet_leaf_13_clk _01956_ _00781_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_10411_ net741 net576 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10342_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10273_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__and2_1
XANTENNA__06927__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout492 top.cb_syn.end_cnt\[2\] vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
Xfanout481 top.histogram.init vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_2
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_2
XANTENNA__10402__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08794__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06155__B2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ clknet_leaf_45_clk _02277_ _01117_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05666__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ clknet_leaf_114_clk _02208_ _01048_ vssd1 vssd1 vccd1 vccd1 top.path\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_11589_ clknet_leaf_30_clk _02154_ _00979_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08604__B1 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ net797 net632 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ top.hTree.tree_reg\[33\] top.findLeastValue.sum\[33\] net283 vssd1 vssd1
+ vccd1 vccd1 _04382_ sky130_fd_sc_hd__mux2_1
X_07751_ _02520_ net387 _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__o21a_1
XANTENNA__07569__S1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ _03492_ _03499_ _03491_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__o21a_1
X_07682_ top.hTree.tree_reg\[59\] _04248_ net389 vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ net959 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07902__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06633_ _02441_ top.findLeastValue.val1\[5\] top.findLeastValue.val1\[4\] _02442_
+ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_32_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ net1288 net225 net215 _04367_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__a22o_1
XANTENNA__09096__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06564_ net453 _03364_ top.controller.fin_HG vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__a21bo_1
X_08303_ top.cb_syn.char_path_n\[53\] net376 net332 top.cb_syn.char_path_n\[51\] net179
+ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a221o_1
XANTENNA__07646__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05515_ net440 top.findLeastValue.wipe_the_char_2 net527 vssd1 vssd1 vccd1 vccd1
+ _02600_ sky130_fd_sc_hd__and3_2
XANTENNA__05657__B1 _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout235_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07646__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06495_ top.histogram.total\[5\] top.histogram.total\[4\] top.histogram.total\[3\]
+ top.histogram.total\[2\] vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__and4_1
X_09283_ top.translation.totalEn _05023_ _05024_ top.translation.writeEn vssd1 vssd1
+ vccd1 vccd1 _05227_ sky130_fd_sc_hd__and4b_1
X_08234_ top.cb_syn.char_path_n\[87\] net198 _04679_ vssd1 vssd1 vccd1 vccd1 _01706_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05446_ net535 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08165_ top.cb_syn.char_path_n\[122\] net373 net327 top.cb_syn.char_path_n\[120\]
+ net176 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout402_A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05377_ top.findLeastValue.val1\[14\] vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__inv_2
X_07116_ _03790_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_41_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08096_ top.cb_syn.num_lefts\[7\] _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08359__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ top.findLeastValue.val2\[38\] top.findLeastValue.val1\[38\] vssd1 vssd1 vccd1
+ vccd1 _03723_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout771_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ top.WB.CPU_DAT_O\[22\] net1212 net366 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
X_07949_ net437 net1564 net251 top.findLeastValue.sum\[8\] _04485_ vssd1 vssd1 vccd1
+ vccd1 _01797_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_67_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_50_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10960_ clknet_leaf_61_clk net1361 _00350_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ net770 net605 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__and2_1
X_10891_ clknet_leaf_33_clk net1483 _00281_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cond
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07812__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936__899 vssd1 vssd1 vccd1 vccd1 _11936__899/HI net899 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05648__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ clknet_leaf_118_clk _02077_ _00902_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11443_ clknet_leaf_90_clk _02008_ _00833_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06163__A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11374_ clknet_leaf_16_clk _01939_ _00764_ vssd1 vssd1 vccd1 vccd1 top.cw1\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08789__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10325_ net728 net563 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__and2_1
X_10256_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__and2_1
XANTENNA__07706__B _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__A0 _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ net802 net637 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_58_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06280_ _03022_ _03150_ _03018_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__o21ai_1
X_05300_ net454 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 top.cb_syn.i\[1\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 top.cb_syn.zero_count\[7\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold704 top.hTree.nullSumIndex\[3\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 top.hTree.state\[4\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold759 top.cb_syn.char_path_n\[117\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__A1 top.findLeastValue.sum\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold748 top.hTree.wait_cnt vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09002__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ _05066_ top.cb_syn.max_index\[6\] _05059_ vssd1 vssd1 vccd1 vccd1 _01406_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08356__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ _02813_ _05038_ _05039_ _05036_ top.translation.index\[6\] vssd1 vssd1 vccd1
+ vccd1 _01448_ sky130_fd_sc_hd__o32a_1
X_07803_ net418 _04367_ _04368_ net260 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout185_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
X_08783_ top.path\[12\] net404 net324 top.path\[13\] top.translation.index\[2\] vssd1
+ vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__o221a_1
X_05995_ top.WB.CPU_DAT_O\[6\] net1142 net347 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
X_07734_ net473 _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nand2_1
XANTENNA__07316__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05590__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ net449 _04255_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__nand2_4
XANTENNA__08728__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ top.hTree.nulls\[61\] _04263_ net401 vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06616_ top.compVal\[21\] _02492_ _02493_ top.compVal\[20\] vssd1 vssd1 vccd1 vccd1
+ _03414_ sky130_fd_sc_hd__a22o_1
XANTENNA__07351__B _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07596_ net412 _02884_ _02886_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07619__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07619__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ net1415 net223 net214 _04435_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__a22o_1
X_06547_ net1593 _03331_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ net1666 _05223_ _05224_ _05207_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06478_ top.hist_data_o\[4\] _03246_ _03315_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_23_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08217_ top.cb_syn.char_path_n\[96\] net370 net326 top.cb_syn.char_path_n\[94\] net172
+ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05429_ top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06842__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ top.controller.fin_reg\[5\] top.controller.fin_reg\[6\] top.controller.fin_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__nand3_1
X_08148_ top.cb_syn.cb_length\[1\] _04636_ net190 vssd1 vssd1 vccd1 vccd1 _01749_
+ sky130_fd_sc_hd__mux2_1
X_08079_ _04566_ _04576_ _02533_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__mux2_1
X_11090_ clknet_leaf_63_clk _01655_ _00480_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07807__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__and2_1
X_10041_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__and2_1
Xhold20 top.sram_interface.init_counter\[20\] vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 top.hTree.node_reg\[44\] vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10233__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold64 top.hTree.node_reg\[42\] vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 top.hTree.node_reg\[9\] vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top.hTree.state\[10\] vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 top.cb_syn.check_right vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net110 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net48 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06857__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05581__A2 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ clknet_leaf_37_clk _01508_ _00333_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07858__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10874_ clknet_leaf_23_clk _01459_ _00264_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_6 _01191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ clknet_leaf_99_clk _01991_ _00816_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[30\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11357_ clknet_leaf_100_clk _01922_ _00747_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_10308_ net839 net674 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__and2_1
XANTENNA__07794__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11288_ clknet_leaf_14_clk _01853_ _00678_ vssd1 vssd1 vccd1 vccd1 top.hTree.closing
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__and2_1
X_05780_ net506 net508 vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or2_2
XANTENNA__05572__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07450_ top.dut.bit_buf\[13\] top.dut.bit_buf\[6\] net713 vssd1 vssd1 vccd1 vccd1
+ _04058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06401_ top.hist_data_o\[15\] top.hist_data_o\[14\] _03255_ vssd1 vssd1 vccd1 vccd1
+ _03266_ sky130_fd_sc_hd__and3_1
X_07381_ _03845_ _04018_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__nand2_1
X_06332_ _02927_ _03019_ _03020_ _03200_ net454 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__o311a_1
X_09120_ _05126_ _05132_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__and2_1
X_09051_ _02552_ _02882_ _02883_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_20_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ _04525_ net1670 _04522_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__mux2_1
X_06263_ top.cb_syn.char_index\[4\] _03044_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__nor2_1
XANTENNA__06824__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold501 net82 vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
X_06194_ top.cb_syn.char_index\[6\] _03036_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold512 top.cb_syn.count\[2\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 top.cb_syn.h_element\[53\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 top.path\[105\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 top.hTree.tree_reg\[2\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 top.hist_data_o\[29\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 top.sram_interface.init_counter\[10\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _03346_ vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 _01559_ vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net771 net606 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__and2_1
X_09884_ net867 net702 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__and2_1
X_08904_ _02418_ net422 _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__nor3_1
X_08835_ top.translation.write_fin top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 _05024_
+ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout567_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ top.path\[88\] net402 net323 top.path\[89\] net429 vssd1 vssd1 vccd1 vccd1
+ _04955_ sky130_fd_sc_hd__o221a_1
XANTENNA__05563__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ _04297_ _04298_ net474 vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__mux2_1
X_05978_ top.WB.CPU_DAT_O\[23\] net1227 net345 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ top.header_synthesis.count\[1\] _04896_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ net1070 _04242_ _04212_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07579_ net516 net521 vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__or2_2
XFILLER_0_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ net1027 net224 net216 _04503_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10590_ net737 net572 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__and2_1
X_09249_ _05207_ _05211_ _05212_ _05208_ net1605 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[2\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__08017__A1 _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ clknet_leaf_107_clk _01776_ _00601_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_11142_ clknet_leaf_52_clk _01707_ _00532_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[88\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
X_11073_ clknet_leaf_53_clk _01638_ _00463_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
X_10024_ net829 net664 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__and2_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05554__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951__914 vssd1 vssd1 vccd1 vccd1 _11951__914/HI net914 sky130_fd_sc_hd__conb_1
X_10926_ clknet_leaf_61_clk _01491_ _00316_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10857_ clknet_leaf_11_clk _01451_ _00247_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.TRN_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ clknet_leaf_117_clk _01394_ _00178_ vssd1 vssd1 vccd1 vccd1 top.path\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_11409_ clknet_leaf_86_clk _01974_ _00799_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[13\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09300__S0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06950_ top.findLeastValue.val1\[7\] net135 net113 net1693 vssd1 vssd1 vccd1 vccd1
+ _01968_ sky130_fd_sc_hd__o22a_1
X_05901_ top.cb_syn.h_element\[52\] top.cb_syn.h_element\[51\] top.cb_syn.h_element\[50\]
+ top.cb_syn.h_element\[53\] vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__or4b_1
XANTENNA__07881__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ top.compVal\[13\] top.findLeastValue.val1\[13\] net154 vssd1 vssd1 vccd1
+ vccd1 _03646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08620_ top.cb_syn.char_path_n\[3\] top.cb_syn.char_path_n\[4\] top.cb_syn.char_path_n\[7\]
+ top.cb_syn.char_path_n\[8\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__mux4_1
X_05832_ top.sram_interface.counter_HTREE\[1\] top.sram_interface.counter_HTREE\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05545__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08551_ net1323 top.cb_syn.char_path_n\[8\] net240 vssd1 vssd1 vccd1 vccd1 _01491_
+ sky130_fd_sc_hd__mux2_1
X_05763_ net1802 net163 net147 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 _02330_
+ sky130_fd_sc_hd__a22o_1
X_08482_ net1163 top.cb_syn.char_path_n\[77\] net245 vssd1 vssd1 vccd1 vccd1 _01560_
+ sky130_fd_sc_hd__mux2_1
X_07502_ _02975_ _04101_ _02974_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_85_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05694_ top.histogram.sram_out\[6\] net358 net408 top.hTree.node_reg\[6\] _02751_
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a221o_1
XANTENNA__09141__C1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07433_ top.dut.bits_in_buf\[2\] _04043_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__xor2_4
XFILLER_0_92_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11887__919 vssd1 vssd1 vccd1 vccd1 net919 _11887__919/LO sky130_fd_sc_hd__conb_1
XANTENNA__05430__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07364_ _03799_ _03852_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_33_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09103_ net1004 net1604 net254 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__mux2_1
X_06315_ _03071_ _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nand2_1
X_07295_ _03789_ _03864_ _03870_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08798__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout315_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06246_ top.cw2\[6\] _03080_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__or2_1
X_09034_ top.WB.CPU_DAT_O\[16\] net1144 net313 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__mux2_1
Xhold320 top.cb_syn.char_path\[37\] vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05481__B2 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 top.cb_syn.char_path\[22\] vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _01576_ vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ top.TRN_char_index\[6\] _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__nand2_1
Xhold331 net102 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout684_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout800 net803 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_1
Xhold386 top.path\[25\] vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 top.path\[21\] vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 top.path\[102\] vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
X_09936_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__and2_1
Xhold397 _01554_ vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_2
Xfanout822 net825 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_2
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_2
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_2
Xfanout855 net859 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_2
Xfanout844 net845 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07791__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout851_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__and2_1
Xfanout877 net34 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
X_09798_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__and2_1
X_08818_ net427 _05005_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__o21a_1
X_08749_ net425 _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__or2_1
X_11760_ clknet_leaf_46_clk _02299_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10711_ clknet_leaf_74_clk _01342_ _00101_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08581__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ clknet_leaf_102_clk _02241_ _01081_ vssd1 vssd1 vccd1 vccd1 top.compVal\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_11911__942 vssd1 vssd1 vccd1 vccd1 net942 _11911__942/LO sky130_fd_sc_hd__conb_1
X_10642_ clknet_leaf_74_clk _01273_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10573_ net833 net668 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__and2_1
XANTENNA__07966__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05472__B2 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ clknet_leaf_62_clk _01690_ _00515_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[71\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08797__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ clknet_leaf_48_clk _01621_ _00446_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_79_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05775__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__and2_1
XANTENNA__05515__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11875__878 vssd1 vssd1 vccd1 vccd1 _11875__878/HI net878 sky130_fd_sc_hd__conb_1
XFILLER_0_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11889_ net920 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ clknet_leaf_3_clk top.controller.fin_TRN _00299_ vssd1 vssd1 vccd1 vccd1
+ top.controller.fin_reg\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08229__B2 top.cb_syn.char_path_n\[88\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06100_ _02450_ _02999_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__nor2_1
XANTENNA__07876__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07080_ _03754_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__nor2_1
X_06031_ net1626 _02928_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_10_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05463__B2 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__B2 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout129 net130 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_4
Xfanout118 net122 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
X_07982_ net477 _04510_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or2_1
X_09721_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__and2_1
X_06933_ top.findLeastValue.val1\[24\] net134 net115 net1127 vssd1 vssd1 vccd1 vccd1
+ _01985_ sky130_fd_sc_hd__o22a_1
X_09652_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__and2_1
X_06864_ top.findLeastValue.val2\[22\] net132 net117 _03637_ vssd1 vssd1 vccd1 vccd1
+ _02030_ sky130_fd_sc_hd__o22a_1
X_08603_ top.cb_syn.char_path_n\[115\] top.cb_syn.char_path_n\[116\] top.cb_syn.char_path_n\[119\]
+ top.cb_syn.char_path_n\[120\] net499 net493 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__mux4_1
X_05815_ _02832_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or2_2
X_09583_ net797 net632 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__and2_1
X_06795_ _03570_ _03571_ _03592_ _03587_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_38_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ net1342 top.cb_syn.char_path_n\[25\] net234 vssd1 vssd1 vccd1 vccd1 _01508_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout265_A _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05746_ top.findLeastValue.alternator_timer\[2\] _02784_ top.findLeastValue.alternator_timer\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__o21a_1
X_08465_ net1074 net1805 net230 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05677_ net1469 net168 _02737_ net209 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08396_ top.cb_syn.char_path_n\[6\] net196 _04760_ vssd1 vssd1 vccd1 vccd1 _01625_
+ sky130_fd_sc_hd__o21a_1
X_07416_ _02520_ net126 net124 _04038_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a2bb2o_1
X_07347_ _03772_ _03977_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_98_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07786__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ net1740 _05081_ _05082_ top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 _01326_
+ sky130_fd_sc_hd__a22o_1
X_07278_ _03874_ _03888_ _03886_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__o21ai_1
X_06229_ _02418_ _02524_ net533 top.sram_interface.word_cnt\[5\] vssd1 vssd1 vccd1
+ vccd1 _03102_ sky130_fd_sc_hd__a31o_2
Xhold161 top.cb_syn.char_path\[80\] vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 top.sram_interface.init_counter\[11\] vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 top.cb_syn.char_path\[13\] vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 top.histogram.sram_out\[21\] vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 top.path\[111\] vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_2
Xfanout641 net643 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_2
X_09919_ net871 net706 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__and2_1
Xfanout685 net689 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_2
Xfanout674 net680 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_2
Xfanout663 net670 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_1
Xfanout652 net661 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_2
Xfanout696 net700 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_107_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ clknet_leaf_82_clk _02345_ _01184_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06865__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11743_ clknet_leaf_10_clk _02293_ _01133_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.write_counter_FLV\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11674_ clknet_leaf_93_clk _02224_ _01064_ vssd1 vssd1 vccd1 vccd1 top.compVal\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10625_ clknet_leaf_65_clk _01256_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06890__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05693__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10556_ net834 net669 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10487_ net838 net673 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__and2_1
XANTENNA__10416__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11108_ clknet_leaf_49_clk _01673_ _00498_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_11039_ clknet_leaf_37_clk _01604_ _00429_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10151__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05600_ top.cb_syn.char_path\[53\] net530 net311 top.cb_syn.char_path\[117\] vssd1
+ vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07370__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07370__B2 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06580_ top.cb_syn.num_lefts\[7\] top.cb_syn.num_lefts\[5\] top.cb_syn.num_lefts\[3\]
+ top.cb_syn.num_lefts\[1\] top.header_synthesis.count\[1\] top.header_synthesis.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_96_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05531_ top.WB.curr_state\[0\] _02572_ _02615_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__and3_1
X_08250_ top.cb_syn.char_path_n\[79\] net205 _04687_ vssd1 vssd1 vccd1 vccd1 _01698_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08990__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05462_ net18 net415 net364 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 _02396_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08181_ top.cb_syn.char_path_n\[114\] net378 net335 top.cb_syn.char_path_n\[112\]
+ net181 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07201_ _03875_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05393_ top.cw2\[2\] vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__inv_2
X_07132_ top.findLeastValue.val2\[11\] top.findLeastValue.val1\[11\] vssd1 vssd1 vccd1
+ vccd1 _03808_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07063_ top.findLeastValue.val2\[25\] top.findLeastValue.val1\[25\] _03738_ vssd1
+ vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06014_ top.sram_interface.init_counter\[3\] _02926_ vssd1 vssd1 vccd1 vccd1 _02927_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_93_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout382_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ top.hTree.tree_reg\[4\] top.findLeastValue.sum\[4\] net284 vssd1 vssd1 vccd1
+ vccd1 _04498_ sky130_fd_sc_hd__mux2_1
X_09704_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__and2_1
X_06916_ top.findLeastValue.val1\[41\] net137 net112 top.compVal\[41\] vssd1 vssd1
+ vccd1 vccd1 _02002_ sky130_fd_sc_hd__o22a_1
X_09635_ net760 net595 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__and2_1
X_07896_ top.hTree.tree_reg\[18\] top.findLeastValue.sum\[18\] net267 vssd1 vssd1
+ vccd1 vccd1 _04443_ sky130_fd_sc_hd__mux2_1
XANTENNA__09350__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06164__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ top.compVal\[30\] top.findLeastValue.val1\[30\] net151 vssd1 vssd1 vccd1
+ vccd1 _03629_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout647_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__and2_1
X_06778_ top.compVal\[23\] top.findLeastValue.val2\[23\] vssd1 vssd1 vccd1 vccd1 _03576_
+ sky130_fd_sc_hd__nand2b_1
X_08517_ net1360 top.cb_syn.char_path_n\[42\] net241 vssd1 vssd1 vccd1 vccd1 _01525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout814_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05729_ top.hTree.node_reg\[32\] net308 _02780_ net469 vssd1 vssd1 vccd1 vccd1 _02781_
+ sky130_fd_sc_hd__a22o_1
X_09497_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__and2_1
X_08448_ net1097 top.cb_syn.char_path_n\[111\] net242 vssd1 vssd1 vccd1 vccd1 _01594_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08861__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05675__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06872__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08379_ top.cb_syn.char_path_n\[15\] net384 net340 top.cb_syn.char_path_n\[13\] net187
+ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a221o_1
X_10410_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__and2_1
X_11390_ clknet_leaf_14_clk _01955_ _00780_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10341_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__and2_1
X_10272_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout493 top.cb_syn.end_cnt\[2\] vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_2
Xfanout482 top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_2
Xfanout460 net462 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 net480 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07888__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11726_ clknet_leaf_47_clk _02276_ _01116_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__B2 top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ clknet_leaf_114_clk _02207_ _01047_ vssd1 vssd1 vccd1 vccd1 top.path\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_11588_ clknet_leaf_31_clk _02153_ _00978_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10608_ net745 net580 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10539_ net728 net563 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__and2_1
XANTENNA__09935__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07750_ net387 _04325_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__nand2_1
XANTENNA__09332__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06701_ _03478_ _03483_ _02413_ top.findLeastValue.val1\[34\] vssd1 vssd1 vccd1 vccd1
+ _03499_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07681_ net257 _04268_ _04269_ net1131 net433 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a32o_1
X_09420_ net963 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06632_ _02439_ top.findLeastValue.val1\[7\] vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__and2_1
X_09351_ net1020 net225 net215 _04371_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__a22o_1
X_06563_ _02454_ top.histogram.state\[0\] vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__and2_1
X_08302_ net1692 net197 _04713_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__o21a_1
X_05514_ net457 _02579_ _02598_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a21oi_1
X_09282_ net343 _04058_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[13\] sky130_fd_sc_hd__and2_1
X_08233_ top.cb_syn.char_path_n\[88\] net377 net330 top.cb_syn.char_path_n\[86\] net180
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a221o_1
XANTENNA__06303__C1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06494_ top.histogram.total\[4\] _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__and2_1
XANTENNA__05657__B2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout130_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06854__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05445_ net455 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_105_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ top.cb_syn.char_path_n\[122\] net191 _04644_ vssd1 vssd1 vccd1 vccd1 _01741_
+ sky130_fd_sc_hd__o21a_1
X_05376_ top.findLeastValue.val1\[20\] vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__inv_2
X_08095_ top.cb_syn.num_lefts\[6\] _04595_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__nand2_1
XANTENNA__07803__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07115_ top.findLeastValue.val2\[14\] top.findLeastValue.val1\[14\] vssd1 vssd1 vccd1
+ vccd1 _03791_ sky130_fd_sc_hd__or2_1
XANTENNA__11797__D net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07046_ top.findLeastValue.val2\[38\] top.findLeastValue.val1\[38\] vssd1 vssd1 vccd1
+ vccd1 _03722_ sky130_fd_sc_hd__nand2_1
XANTENNA__08359__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ top.WB.CPU_DAT_O\[23\] net1335 net365 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
XANTENNA__05593__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ net420 _04483_ _04484_ net262 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__o211a_1
XANTENNA__09323__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ net438 net1557 net248 net1807 _04429_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a221o_1
X_09618_ net769 net604 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__and2_1
X_10890_ clknet_leaf_32_clk _01462_ _00280_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.pulse_first
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ net723 net558 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__and2_1
XANTENNA__05896__A1 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08834__A1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ clknet_leaf_117_clk _02076_ _00901_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ clknet_leaf_106_clk _02007_ _00832_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[46\]
+ sky130_fd_sc_hd__dfstp_2
X_11373_ clknet_leaf_15_clk _01938_ _00763_ vssd1 vssd1 vccd1 vccd1 top.cw1\[5\] sky130_fd_sc_hd__dfrtp_1
X_10324_ net731 net566 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__and2_1
X_10186_ net802 net637 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__and2_1
Xfanout290 _04111_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_2
XANTENNA__05584__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05887__A1 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05639__A1 top.hTree.node_reg\[47\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ clknet_leaf_80_clk _02259_ _01099_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06836__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold716 top.compVal\[25\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold705 top.findLeastValue.sum\[29\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 top.sram_interface.TRN_counter\[1\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold738 top.hist_data_o\[16\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 top.compVal\[0\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08920_ _04217_ _05065_ _04255_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__mux2_1
X_08851_ _02550_ _05036_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__nand2_1
X_07802_ net476 _04366_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__or2_1
XANTENNA__05575__B1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ net426 _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__or2_1
X_05994_ top.WB.CPU_DAT_O\[7\] net1076 net347 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
X_07733_ _02517_ net388 _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__o21a_1
X_07664_ net433 _04254_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__nor2_2
XANTENNA__08728__B net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09403_ net1029 net221 _05281_ _05282_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a22o_1
XANTENNA__05878__A1 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06615_ _02429_ top.findLeastValue.val1\[23\] vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__and2_1
X_07595_ net519 _02884_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08277__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ net1363 net223 net214 _04439_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__a22o_1
X_06546_ _03356_ _03357_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__nor2_1
X_09265_ top.cb_syn.zero_count\[7\] _05222_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__nor2_1
X_06477_ top.hist_data_o\[4\] _03246_ net297 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_23_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08216_ top.cb_syn.char_path_n\[96\] net192 _04670_ vssd1 vssd1 vccd1 vccd1 _01715_
+ sky130_fd_sc_hd__o21a_1
X_05428_ top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__inv_2
X_09196_ top.controller.fin_reg\[1\] top.controller.fin_reg\[4\] top.controller.fin_reg\[3\]
+ top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08147_ _04632_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__nor2_1
X_05359_ top.findLeastValue.val2\[8\] vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__inv_2
X_08078_ _03386_ _04567_ _04576_ _04566_ net1717 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a32o_1
X_07029_ top.findLeastValue.val1\[6\] top.findLeastValue.val1\[5\] top.findLeastValue.val1\[4\]
+ top.findLeastValue.val1\[3\] vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__and4_1
X_10040_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__and2_1
Xhold10 top.sram_interface.init_counter\[23\] vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 top.sram_interface.init_counter\[17\] vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 top.hTree.node_reg\[25\] vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 top.hTree.tree_reg\[50\] vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05566__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 top.hTree.node_reg\[34\] vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _01786_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 top.hTree.node_reg\[50\] vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 top.hTree.node_reg\[5\] vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 top.hTree.node_reg\[3\] vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
X_10942_ clknet_leaf_52_clk _01507_ _00332_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05869__A1 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ clknet_leaf_27_clk _01458_ _00263_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06873__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06818__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ clknet_leaf_99_clk _01990_ _00815_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[29\]
+ sky130_fd_sc_hd__dfstp_2
X_11356_ clknet_leaf_100_clk _01921_ _00746_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08991__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ net840 net675 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__and2_1
XANTENNA__07794__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06597__A2 _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__B2 top.findLeastValue.sum\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ clknet_leaf_104_clk _01852_ _00677_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__and2_1
XANTENNA__05557__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10169_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06400_ top.hist_data_o\[30\] _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ _03842_ _03845_ _03847_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__nand3_1
X_06331_ top.hist_addr\[3\] top.hist_addr\[2\] top.hist_addr\[1\] top.hist_addr\[0\]
+ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a41o_1
XFILLER_0_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06262_ top.cb_syn.max_index\[6\] _03102_ _03104_ top.hTree.nullSumIndex\[5\] vssd1
+ vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ top.WB.CPU_DAT_O\[0\] net1533 net316 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ top.findLeastValue.least2\[5\] top.findLeastValue.least1\[5\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06193_ top.TRN_char_index\[6\] _03051_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__or2_1
Xhold502 top.path\[73\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 top.hTree.nulls\[51\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 top.hTree.node_reg\[38\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 top.histogram.sram_out\[5\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__and2_1
Xhold557 top.header_synthesis.count\[4\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08982__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold579 net77 vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 top.hTree.tree_reg\[43\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 top.histogram.total\[11\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _02522_ _02831_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05428__A top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05548__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08834_ top.translation.index\[4\] _04962_ _04969_ _05017_ _05022_ vssd1 vssd1 vccd1
+ vccd1 _05023_ sky130_fd_sc_hd__a32o_1
X_08765_ top.path\[90\] top.path\[91\] net508 vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__mux2_1
X_07716_ top.findLeastValue.least2\[7\] _04297_ net389 vssd1 vssd1 vccd1 vccd1 _04298_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout462_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05977_ top.WB.CPU_DAT_O\[24\] net1154 net345 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ top.header_synthesis.count\[4\] top.header_synthesis.count\[3\] top.header_synthesis.count\[2\]
+ top.header_synthesis.count\[1\] vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_0_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07647_ top.cb_syn.max_index\[2\] _04181_ _04238_ _04241_ vssd1 vssd1 vccd1 vccd1
+ _04242_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07578_ net519 net524 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__or2_2
XANTENNA__05720__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06529_ top.histogram.total\[19\] _03335_ net1520 vssd1 vssd1 vccd1 vccd1 _03351_
+ sky130_fd_sc_hd__a21oi_1
X_09317_ net1109 net224 net215 _04507_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__a22o_1
X_09248_ _02558_ _05209_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_09179_ net1592 top.controller.fin_reg\[7\] _05172_ vssd1 vssd1 vccd1 vccd1 _00013_
+ sky130_fd_sc_hd__and3_1
X_11210_ clknet_leaf_107_clk _01775_ _00600_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11141_ clknet_leaf_53_clk _01706_ _00531_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[87\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_112_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
X_11072_ clknet_leaf_54_clk _01637_ _00462_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__05539__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ net855 net690 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__and2_1
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925_ clknet_leaf_65_clk _01490_ _00315_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05711__B1 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ clknet_leaf_11_clk _01450_ _00246_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.TRN_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10787_ clknet_leaf_117_clk _01393_ _00177_ vssd1 vssd1 vccd1 vccd1 top.path\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09199__B top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10419__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05536__A_N net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11408_ clknet_leaf_86_clk _01973_ _00798_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09300__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__A0 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ clknet_leaf_77_clk _01904_ _00729_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05900_ top.cb_syn.h_element\[49\] top.cb_syn.h_element\[48\] top.cb_syn.h_element\[47\]
+ top.cb_syn.h_element\[46\] vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__or4_1
XANTENNA__06990__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06880_ top.findLeastValue.val2\[14\] net130 net122 _03645_ vssd1 vssd1 vccd1 vccd1
+ _02022_ sky130_fd_sc_hd__o22a_1
X_05831_ _02514_ _02522_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nor2_1
XANTENNA__08811__S0 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ net1368 top.cb_syn.char_path_n\[9\] net240 vssd1 vssd1 vccd1 vccd1 _01492_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08993__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05762_ _02564_ net162 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__nor2_2
X_08481_ net1513 top.cb_syn.char_path_n\[78\] net245 vssd1 vssd1 vccd1 vccd1 _01561_
+ sky130_fd_sc_hd__mux2_1
X_07501_ _02980_ _02984_ _02982_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_85_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05693_ top.hTree.node_reg\[38\] net307 _02750_ net469 vssd1 vssd1 vccd1 vccd1 _02751_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05702__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07432_ _02405_ top.dut.bits_in_buf\[1\] top.dut.bits_in_buf\[0\] vssd1 vssd1 vccd1
+ vccd1 _04043_ sky130_fd_sc_hd__or3_2
XANTENNA__07402__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ top.hTree.wait_cnt net1522 net254 _05091_ net1542 vssd1 vssd1 vccd1 vccd1
+ _00027_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_33_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07363_ net273 _04005_ _04006_ net279 net1559 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a32o_1
X_06314_ top.cw1\[3\] _03070_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__nand2_1
X_07294_ _03865_ _03869_ _03739_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__o21ai_1
X_06245_ top.cw1\[6\] _03072_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__nor2_1
X_09033_ top.WB.CPU_DAT_O\[17\] net1263 net313 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout210_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold310 net66 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
X_06176_ top.TRN_char_index\[5\] top.TRN_char_index\[4\] _03050_ vssd1 vssd1 vccd1
+ vccd1 _03051_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout308_A _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 top.cb_syn.char_path\[117\] vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__A0 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold332 top.path\[58\] vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 top.path\[120\] vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 net78 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 top.cb_syn.char_path\[6\] vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 top.histogram.sram_out\[17\] vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05769__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 top.dut.out\[4\] vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ net794 net629 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__and2_1
Xhold398 top.cb_syn.char_path\[39\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout823 net825 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_2
Xfanout801 net802 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_2
Xfanout812 net816 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_2
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_2
Xfanout867 net876 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_2
X_09866_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__and2_1
Xfanout856 net858 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_2
Xfanout845 net877 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ top.path\[104\] net405 net325 top.path\[105\] net430 vssd1 vssd1 vccd1 vccd1
+ _05006_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_116_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09797_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout844_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07930__A1 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ top.path\[26\] top.path\[27\] net509 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__mux2_1
XANTENNA__05941__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ _04879_ _04883_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nor2_1
X_10710_ clknet_leaf_104_clk _01341_ _00100_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ clknet_leaf_76_clk _02240_ _01080_ vssd1 vssd1 vccd1 vccd1 top.compVal\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ clknet_leaf_76_clk _01272_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10572_ net860 net695 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08651__B _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ clknet_leaf_56_clk _01689_ _00514_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[70\]
+ sky130_fd_sc_hd__dfrtp_2
X_11055_ clknet_leaf_39_clk _01620_ _00445_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[1\]
+ sky130_fd_sc_hd__dfstp_2
X_10006_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__and2_1
XANTENNA__07921__A1 top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05932__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ clknet_leaf_33_clk _01480_ _00298_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_check
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11888_ net884 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08229__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839_ clknet_leaf_116_clk _01433_ _00229_ vssd1 vssd1 vccd1 vccd1 top.path\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08634__C1 _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07532__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05999__A0 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06030_ _02929_ _02936_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__nor2_1
XANTENNA__05463__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout119 net121 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
X_07981_ top.hTree.tree_reg\[1\] top.findLeastValue.sum\[1\] net267 vssd1 vssd1 vccd1
+ vccd1 _04511_ sky130_fd_sc_hd__mux2_1
X_09720_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__and2_1
X_06932_ top.findLeastValue.val1\[25\] net134 net115 net1667 vssd1 vssd1 vccd1 vccd1
+ _01986_ sky130_fd_sc_hd__o22a_1
XANTENNA__10612__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__and2_1
X_11893__924 vssd1 vssd1 vccd1 vccd1 net924 _11893__924/LO sky130_fd_sc_hd__conb_1
X_06863_ top.compVal\[22\] top.findLeastValue.val1\[22\] net156 vssd1 vssd1 vccd1
+ vccd1 _03637_ sky130_fd_sc_hd__mux2_1
X_08602_ _02542_ _04821_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__and2_1
X_05814_ top.findLeastValue.least2\[8\] _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nand2_1
X_09582_ net748 net583 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__and2_1
X_06794_ _03567_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__nand2_1
X_08533_ net1128 top.cb_syn.char_path_n\[26\] net236 vssd1 vssd1 vccd1 vccd1 _01509_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05745_ _02783_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout160_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ net1329 top.cb_syn.char_path_n\[95\] net233 vssd1 vssd1 vccd1 vccd1 _01578_
+ sky130_fd_sc_hd__mux2_1
X_05676_ top.histogram.sram_out\[9\] net357 net408 top.hTree.node_reg\[9\] _02736_
+ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_18_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ top.cb_syn.char_path_n\[7\] net375 net332 top.cb_syn.char_path_n\[5\] net178
+ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a221o_1
X_07415_ net487 top.findLeastValue.least1\[1\] net149 vssd1 vssd1 vccd1 vccd1 _04038_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout425_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ net1706 net274 net269 _03994_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XANTENNA__07523__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07979__B2 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ net1797 _05081_ _05082_ top.TRN_char_index\[1\] vssd1 vssd1 vccd1 vccd1 _01327_
+ sky130_fd_sc_hd__a22o_1
X_07277_ net270 _03933_ _03943_ net276 top.findLeastValue.sum\[36\] vssd1 vssd1 vccd1
+ vccd1 _01923_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06228_ _03019_ _03096_ _03100_ net454 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold162 _01563_ vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _02169_ vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
X_06159_ top.cb_syn.char_index\[2\] top.cb_syn.char_index\[1\] vssd1 vssd1 vccd1 vccd1
+ _03034_ sky130_fd_sc_hd__nand2_1
Xhold140 top.path\[6\] vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 top.path\[72\] vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 top.path\[83\] vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 top.path\[126\] vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__and2_1
Xfanout620 net621 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06954__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout631 net44 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_2
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_1
Xfanout675 net679 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09353__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 net661 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_1
Xfanout664 net665 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_2
Xfanout686 net689 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlymetal6s2s_1
X_09849_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__and2_1
Xfanout697 net700 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_107_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ clknet_leaf_82_clk _02344_ _01183_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
X_11742_ clknet_leaf_4_clk _02292_ _01132_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.write_counter_FLV\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11673_ clknet_leaf_93_clk _02223_ _01063_ vssd1 vssd1 vccd1 vccd1 top.compVal\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10624_ clknet_leaf_82_clk _01255_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06881__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05693__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07514__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10555_ net834 net669 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10486_ net839 net674 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08395__A1 top.cb_syn.char_path_n\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881__883 vssd1 vssd1 vccd1 vccd1 _11881__883/HI net883 sky130_fd_sc_hd__conb_1
X_11107_ clknet_leaf_48_clk _01672_ _00497_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[53\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06910__A _03394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09344__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ clknet_leaf_50_clk _01603_ _00428_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10151__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05526__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09940__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11918__949 vssd1 vssd1 vccd1 vccd1 net949 _11918__949/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05530_ _02599_ _02614_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05461_ net19 net414 net363 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 _02397_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_15_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05684__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ net1737 net199 _04652_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__o21a_1
X_05392_ top.cw2\[3\] vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ top.findLeastValue.val2\[34\] top.findLeastValue.val1\[34\] vssd1 vssd1 vccd1
+ vccd1 _03876_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07131_ top.findLeastValue.val2\[11\] top.findLeastValue.val1\[11\] vssd1 vssd1 vccd1
+ vccd1 _03807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07062_ top.findLeastValue.val2\[25\] top.findLeastValue.val1\[25\] top.findLeastValue.val1\[24\]
+ top.findLeastValue.val2\[24\] vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__a22o_1
X_06013_ top.sram_interface.init_counter\[2\] top.sram_interface.init_counter\[1\]
+ top.sram_interface.init_counter\[0\] vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_93_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06936__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ net436 net1579 net249 top.findLeastValue.sum\[5\] _04497_ vssd1 vssd1 vccd1
+ vccd1 _01794_ sky130_fd_sc_hd__a221o_1
X_09703_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__and2_1
X_07895_ top.hTree.tree_reg\[18\] top.findLeastValue.sum\[18\] net286 vssd1 vssd1
+ vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
XANTENNA__09335__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ top.findLeastValue.val1\[42\] net137 net112 net1636 vssd1 vssd1 vccd1 vccd1
+ _02003_ sky130_fd_sc_hd__o22a_1
X_09634_ net760 net595 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06846_ top.findLeastValue.val2\[31\] net127 net118 _03628_ vssd1 vssd1 vccd1 vccd1
+ _02039_ sky130_fd_sc_hd__o22a_1
XANTENNA__05870__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ net780 net615 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__and2_1
X_06777_ top.compVal\[22\] top.findLeastValue.val2\[22\] vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__xnor2_1
X_08516_ net1402 top.cb_syn.char_path_n\[43\] net244 vssd1 vssd1 vccd1 vccd1 _01526_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05728_ _02778_ _02779_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__or2_2
X_09496_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ net1061 top.cb_syn.char_path_n\[112\] net242 vssd1 vssd1 vccd1 vccd1 _01595_
+ sky130_fd_sc_hd__mux2_1
X_05659_ net1462 net168 _02722_ net210 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout807_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05675__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ top.cb_syn.char_path_n\[15\] net205 _04751_ vssd1 vssd1 vccd1 vccd1 _01634_
+ sky130_fd_sc_hd__o21a_1
X_07329_ _03763_ _03981_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__nand2_1
X_10340_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__and2_1
X_10271_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__and2_1
XANTENNA__06927__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 top.sram_interface.write_HT_fin_n vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_1
Xfanout472 net474 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_2
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_2
Xfanout483 top.findLeastValue.histo_index\[5\] vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11725_ clknet_leaf_45_clk _02275_ _01115_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05666__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ clknet_leaf_115_clk _02206_ _01046_ vssd1 vssd1 vccd1 vccd1 top.path\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_11587_ clknet_leaf_30_clk _02152_ _00977_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10607_ net743 net578 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ net717 net552 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09935__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ net829 net664 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06918__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ _03495_ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__nor2_1
X_07680_ net472 _04266_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__or2_1
XANTENNA__07879__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06631_ top.findLeastValue.val1\[12\] top.compVal\[12\] vssd1 vssd1 vccd1 vccd1 _03429_
+ sky130_fd_sc_hd__and2b_1
X_09350_ net976 net225 net215 _04375_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__a22o_1
XANTENNA__08828__C1 top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06562_ net1578 _03324_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__xor2_1
X_08301_ top.cb_syn.char_path_n\[54\] net376 net329 top.cb_syn.char_path_n\[52\] net179
+ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05513_ _02584_ _02592_ _02597_ _02595_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__or4b_1
X_09281_ net343 _04062_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[12\] sky130_fd_sc_hd__and2_1
X_08232_ top.cb_syn.char_path_n\[88\] net194 _04678_ vssd1 vssd1 vccd1 vccd1 _01707_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05657__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06493_ top.histogram.total\[3\] top.histogram.total\[2\] _03325_ vssd1 vssd1 vccd1
+ vccd1 _03326_ sky130_fd_sc_hd__and3_1
XANTENNA__06815__A _03394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05444_ top.dut.out_valid vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__inv_2
X_08163_ top.cb_syn.char_path_n\[123\] net369 net326 top.cb_syn.char_path_n\[121\]
+ net173 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a221o_1
X_05375_ top.findLeastValue.val1\[21\] vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__inv_2
X_08094_ _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__inv_2
X_07114_ top.findLeastValue.val2\[14\] top.findLeastValue.val1\[14\] vssd1 vssd1 vccd1
+ vccd1 _03790_ sky130_fd_sc_hd__nand2_1
X_07045_ top.findLeastValue.val2\[39\] top.findLeastValue.val1\[39\] vssd1 vssd1 vccd1
+ vccd1 _03721_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11899__930 vssd1 vssd1 vccd1 vccd1 net930 _11899__930/LO sky130_fd_sc_hd__conb_1
X_08996_ top.WB.CPU_DAT_O\[24\] net1340 net366 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07947_ net478 _04482_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout757_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ net417 _04427_ _04428_ net263 vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06829_ top.compVal\[39\] top.findLeastValue.val1\[39\] net152 vssd1 vssd1 vccd1
+ vccd1 _03620_ sky130_fd_sc_hd__mux2_1
X_09617_ net733 net568 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09548_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09479_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__and2_1
X_11510_ clknet_leaf_119_clk _02075_ _00900_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05648__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08416__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11441_ clknet_leaf_94_clk _02006_ _00831_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[45\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06444__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ clknet_leaf_15_clk _01937_ _00762_ vssd1 vssd1 vccd1 vccd1 top.cw1\[4\] sky130_fd_sc_hd__dfrtp_2
X_10323_ net730 net565 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__and2_1
X_10185_ net802 net637 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__and2_1
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_66_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08825__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ clknet_leaf_80_clk _02258_ _01098_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11639_ clknet_leaf_98_clk _02189_ _01029_ vssd1 vssd1 vccd1 vccd1 top.path\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold706 top.hTree.nullSumIndex\[1\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 top.histogram.total\[4\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 top.controller.fin_reg\[5\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold739 top.sram_interface.counter_HTREE\[1\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08850_ top.translation.index\[5\] _02812_ top.translation.index\[6\] vssd1 vssd1
+ vccd1 vccd1 _05038_ sky130_fd_sc_hd__o21a_1
XANTENNA__08996__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ top.hTree.tree_reg\[37\] top.findLeastValue.sum\[37\] net266 vssd1 vssd1
+ vccd1 vccd1 _04367_ sky130_fd_sc_hd__mux2_1
X_08781_ top.path\[14\] top.path\[15\] net510 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__mux2_1
X_05993_ top.WB.CPU_DAT_O\[8\] net1201 net347 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
X_07732_ net388 _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand2_1
XANTENNA__07316__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ top.hTree.write_HT_fin _02837_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or2_4
X_09402_ top.hTree.nulls\[60\] net401 net229 vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o21a_1
X_06614_ top.controller.fin_FLV _02500_ net456 _03411_ vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__and4b_2
X_07594_ net550 _04189_ _04190_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a21oi_1
X_09333_ net1252 net226 net218 _04443_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout240_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06545_ top.histogram.total\[9\] _03331_ net1632 vssd1 vssd1 vccd1 vccd1 _03357_
+ sky130_fd_sc_hd__a21oi_1
X_09264_ _05207_ _05222_ _05208_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a21o_1
X_06476_ net1464 net297 _03313_ _03314_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _04541_ _04548_ _05179_ _02543_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__o22ai_1
X_05427_ top.header_synthesis.count\[0\] vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__inv_2
X_08215_ top.cb_syn.char_path_n\[97\] net370 net328 top.cb_syn.char_path_n\[95\] net174
+ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08146_ _04630_ _04631_ _04611_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout505_A top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05358_ top.findLeastValue.val2\[9\] vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__inv_2
X_08077_ _04568_ _04576_ _04582_ _04566_ net1703 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05289_ top.compVal\[45\] vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07028_ top.findLeastValue.val1\[14\] top.findLeastValue.val1\[13\] top.findLeastValue.val1\[12\]
+ top.findLeastValue.val1\[11\] vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07004__B2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 top.sram_interface.init_counter\[16\] vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 top.hTree.node_reg\[32\] vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ top.WB.CPU_DAT_O\[22\] top.cb_syn.h_element\[54\] net368 vssd1 vssd1 vccd1
+ vccd1 _01359_ sky130_fd_sc_hd__mux2_1
Xhold33 top.hTree.node_reg\[43\] vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 top.hTree.node_reg\[23\] vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 top.hTree.node_reg\[10\] vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 top.cb_syn.char_index\[7\] vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 top.hTree.node_reg\[16\] vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 top.hTree.node_reg\[11\] vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 top.hTree.tree_reg\[61\] vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ clknet_leaf_51_clk _01506_ _00331_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ clknet_leaf_27_clk _01457_ _00262_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11424_ clknet_leaf_99_clk _01989_ _00814_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[28\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_8 _03182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11355_ clknet_leaf_100_clk _01920_ _00745_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[33\]
+ sky130_fd_sc_hd__dfrtp_2
X_10306_ net840 net675 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__and2_1
X_11286_ clknet_leaf_14_clk _01851_ _00676_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_10237_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__and2_1
XANTENNA__08743__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10168_ net820 net655 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__and2_1
X_10099_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08259__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ _02416_ _03098_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06261_ top.TRN_char_index\[4\] _03050_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_20_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07482__A1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08000_ _04524_ net1728 _04522_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__mux2_1
X_06192_ top.TRN_char_index\[6\] _03057_ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__o21a_1
Xhold514 _02095_ vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 top.histogram.sram_out\[0\] vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 top.FLV_done vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 top.histogram.total\[26\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11926__889 vssd1 vssd1 vccd1 vccd1 _11926__889/HI net889 sky130_fd_sc_hd__conb_1
X_09951_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__and2_1
Xhold558 top.hist_data_o\[26\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06812__B _03609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold547 top.histogram.sram_out\[2\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 top.histogram.total\[20\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06993__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ net1239 top.WB.CPU_DAT_O\[0\] net305 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__mux2_1
X_09882_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout190_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05548__B2 top.hTree.node_reg\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__inv_2
X_05976_ top.WB.CPU_DAT_O\[25\] net1172 net345 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
X_08764_ top.path\[92\] net402 _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__o21a_1
X_07715_ top.findLeastValue.least2\[7\] top.hTree.tree_reg\[53\] _04248_ vssd1 vssd1
+ vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _02544_ _03389_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__A2_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout455_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ net521 _04237_ _04240_ net516 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout622_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ top.cb_syn.h_element\[61\] top.cb_syn.h_element\[52\] _04176_ vssd1 vssd1
+ vccd1 vccd1 _04177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ net1096 net224 net215 _04511_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__a22o_1
X_06528_ _03337_ _03350_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ _02558_ _05209_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nand2_1
XANTENNA__06276__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06459_ net1366 _03303_ net300 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ top.controller.fin_reg\[1\] top.controller.fin_reg\[2\] top.controller.fin_reg\[3\]
+ top.controller.fin_reg\[5\] vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__nor4_1
X_08129_ top.cb_syn.cb_length\[5\] _04611_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nand2_1
X_11140_ clknet_leaf_53_clk _01705_ _00530_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__clkbuf_4
X_11071_ clknet_leaf_57_clk _01636_ _00461_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[17\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10022_ net830 net665 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__and2_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10924_ clknet_leaf_71_clk _01489_ _00314_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10855_ clknet_leaf_2_clk _01449_ _00245_ vssd1 vssd1 vccd1 vccd1 top.translation.writeEn
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05711__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ clknet_leaf_114_clk _01392_ _00176_ vssd1 vssd1 vccd1 vccd1 top.path\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ clknet_leaf_87_clk _01972_ _00797_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[11\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_74_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11338_ clknet_leaf_77_clk _01903_ _00728_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11269_ clknet_leaf_69_clk _01834_ _00659_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05830_ net443 _02849_ net401 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__or3_1
XANTENNA__08811__S1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05950__B2 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ net1628 top.dut.out_valid_next _04061_ _04083_ _04100_ vssd1 vssd1 vccd1
+ vccd1 _01861_ sky130_fd_sc_hd__o221a_1
X_05761_ net442 net536 _02564_ _02804_ _02803_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a221o_2
X_08480_ net1197 top.cb_syn.char_path_n\[79\] net243 vssd1 vssd1 vccd1 vccd1 _01562_
+ sky130_fd_sc_hd__mux2_1
X_05692_ _02748_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_85_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07431_ net344 vssd1 vssd1 vccd1 vccd1 top.dut.out_valid_next sky130_fd_sc_hd__inv_2
X_07362_ _03801_ _03802_ _03999_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nand3_1
X_06313_ net68 net165 _03182_ net208 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a22o_1
X_09101_ top.hTree.wait_cnt net255 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07293_ _03865_ _03868_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06244_ net1379 net164 _03116_ net207 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
X_09032_ top.WB.CPU_DAT_O\[18\] net1300 net313 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
Xhold311 top.cb_syn.char_path\[87\] vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 top.histogram.sram_out\[30\] vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ top.TRN_char_index\[3\] net445 top.TRN_char_index\[1\] vssd1 vssd1 vccd1
+ vccd1 _03050_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout203_A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 _01600_ vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 top.cb_syn.char_path\[61\] vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 top.cb_syn.char_path\[7\] vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 top.cb_syn.char_path\[121\] vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05769__B2 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 top.path\[125\] vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 top.path\[127\] vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09853__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__and2_1
XANTENNA__06430__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold399 top.hTree.tree_reg\[19\] vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 net816 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_2
Xfanout824 net825 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_1
Xfanout802 net803 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_2
Xhold388 top.path\[33\] vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
X_09865_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__and2_1
Xfanout846 net854 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05873__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net858 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_2
Xfanout835 net877 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 net876 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_2
X_08816_ top.path\[106\] top.path\[107\] net510 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__mux2_1
X_09796_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__and2_1
XANTENNA__07391__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05959_ net1804 net160 net143 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 _02219_
+ sky130_fd_sc_hd__a22o_1
X_08747_ top.path\[112\] top.path\[113\] top.path\[114\] top.path\[115\] net508 net506
+ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__mux4_1
XANTENNA__05941__B2 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ _04887_ _04885_ net1649 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07629_ net517 top.cb_syn.h_element\[49\] net525 top.cb_syn.h_element\[58\] _04180_
+ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__a221o_1
X_10640_ clknet_leaf_73_clk _01271_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ net860 net695 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08424__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07997__A2 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06452__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ clknet_leaf_70_clk _01688_ _00513_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[69\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06879__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ clknet_leaf_32_clk _01619_ _00444_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.state8
+ sky130_fd_sc_hd__dfrtp_1
X_10005_ net841 net676 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05515__C net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05932__B2 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ clknet_leaf_32_clk _01479_ _00297_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.check_right
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05696__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ net919 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_73_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ clknet_leaf_115_clk _01432_ _00228_ vssd1 vssd1 vccd1 vccd1 top.path\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10769_ clknet_leaf_111_clk _01375_ _00159_ vssd1 vssd1 vccd1 vccd1 top.path\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07532__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09954__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ top.hTree.tree_reg\[1\] top.findLeastValue.sum\[1\] net284 vssd1 vssd1 vccd1
+ vccd1 _04510_ sky130_fd_sc_hd__mux2_1
XANTENNA__05620__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06931_ top.findLeastValue.val1\[26\] net134 net115 top.compVal\[26\] vssd1 vssd1
+ vccd1 vccd1 _01987_ sky130_fd_sc_hd__o22a_1
XANTENNA__08165__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08601_ top.cb_syn.char_path_n\[113\] top.cb_syn.char_path_n\[114\] top.cb_syn.char_path_n\[117\]
+ top.cb_syn.char_path_n\[118\] net499 net493 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__mux4_1
X_06862_ top.findLeastValue.val2\[23\] net132 net117 _03636_ vssd1 vssd1 vccd1 vccd1
+ _02031_ sky130_fd_sc_hd__o22a_1
X_05813_ _02833_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__nor2_1
X_09581_ net745 net580 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06793_ _03577_ _03589_ _03590_ top.findLeastValue.val2\[24\] _02428_ vssd1 vssd1
+ vccd1 vccd1 _03591_ sky130_fd_sc_hd__a32o_1
X_08532_ net1384 top.cb_syn.char_path_n\[27\] net234 vssd1 vssd1 vccd1 vccd1 _01510_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05744_ top.findLeastValue.alternator_timer\[3\] top.findLeastValue.alternator_timer\[2\]
+ net406 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09114__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ net1158 top.cb_syn.char_path_n\[96\] net232 vssd1 vssd1 vccd1 vccd1 _01579_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07413__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ _02519_ net126 net124 _04037_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a2bb2o_1
X_05675_ top.hTree.node_reg\[41\] net308 _02735_ net469 vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout153_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05687__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08394_ top.cb_syn.char_path_n\[7\] net197 _04759_ vssd1 vssd1 vccd1 vccd1 _01626_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07428__A1 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ _03768_ _03990_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_30_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07523__S1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05868__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ _03732_ _03890_ _03893_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout418_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06227_ top.hist_addr\[6\] _03099_ net481 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a21o_1
X_09015_ top.hist_addr\[2\] _05081_ _05082_ net445 vssd1 vssd1 vccd1 vccd1 _01328_
+ sky130_fd_sc_hd__a22o_1
X_11941__904 vssd1 vssd1 vccd1 vccd1 _11941__904/HI net904 sky130_fd_sc_hd__conb_1
Xhold130 top.header_synthesis.header\[1\] vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 top.hTree.tree_reg\[58\] vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ _02610_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__nor2_1
Xhold152 top.translation.writeEn vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__A0 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06089_ _02535_ top.cb_syn.i\[3\] vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__and2_1
Xhold185 top.cb_syn.char_path\[52\] vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 top.histogram.sram_out\[15\] vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 top.path\[27\] vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05611__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_2
X_09917_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__and2_1
Xhold196 top.header_synthesis.header\[2\] vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout621 net630 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout632 net638 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08156__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net679 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_1
Xfanout665 net670 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_97_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout643 net651 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_2
Xfanout654 net661 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_2
Xfanout687 net688 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_2
X_09848_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__and2_1
Xfanout698 net700 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_1
X_09779_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ clknet_leaf_82_clk _02343_ _01182_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
X_11741_ clknet_leaf_4_clk _02291_ _01131_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.write_counter_FLV\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05678__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ clknet_leaf_93_clk _02222_ _01062_ vssd1 vssd1 vccd1 vccd1 top.compVal\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10623_ clknet_leaf_81_clk _01254_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06890__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07514__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ net862 net697 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_21_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10485_ net839 net674 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09041__A0 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ clknet_leaf_48_clk _01671_ _00496_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[52\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05602__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
X_11037_ clknet_leaf_51_clk _01602_ _00427_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05526__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11939_ net902 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_82_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05669__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05460_ net20 net416 _02570_ top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 _02398_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05391_ top.cw2\[4\] vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_12_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07130_ _03804_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__nor2_1
X_07061_ top.findLeastValue.val2\[24\] top.findLeastValue.val1\[24\] vssd1 vssd1 vccd1
+ vccd1 _03737_ sky130_fd_sc_hd__nand2_1
XANTENNA__09684__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06012_ top.sram_interface.init_counter\[1\] top.sram_interface.init_counter\[0\]
+ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__and3_1
XANTENNA__05841__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901__932 vssd1 vssd1 vccd1 vccd1 net932 _11901__932/LO sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_79_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
X_07963_ net419 _04495_ _04496_ net261 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__o211a_1
X_09702_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__and2_1
X_07894_ net438 net1350 net252 top.findLeastValue.sum\[19\] _04441_ vssd1 vssd1 vccd1
+ vccd1 _01808_ sky130_fd_sc_hd__a221o_1
X_06914_ top.findLeastValue.val1\[43\] net135 net113 net1730 vssd1 vssd1 vccd1 vccd1
+ _02004_ sky130_fd_sc_hd__o22a_1
X_09633_ net760 net595 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__and2_1
X_06845_ top.compVal\[31\] top.findLeastValue.val1\[31\] net151 vssd1 vssd1 vccd1
+ vccd1 _03628_ sky130_fd_sc_hd__mux2_1
X_09564_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout270_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ net1322 top.cb_syn.char_path_n\[44\] net244 vssd1 vssd1 vccd1 vccd1 _01527_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05452__A top.WB.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06776_ top.compVal\[29\] _02465_ _03572_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_
+ sky130_fd_sc_hd__o211a_1
X_05727_ top.cb_syn.char_path\[32\] net528 net309 top.cb_syn.char_path\[96\] vssd1
+ vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a22o_1
X_09495_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__and2_1
X_08446_ net1149 top.cb_syn.char_path_n\[113\] net243 vssd1 vssd1 vccd1 vccd1 _01596_
+ sky130_fd_sc_hd__mux2_1
X_05658_ top.histogram.sram_out\[12\] net358 net409 top.hTree.node_reg\[12\] _02721_
+ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a221o_1
X_08377_ top.cb_syn.char_path_n\[16\] net385 net340 top.cb_syn.char_path_n\[14\] net188
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_102_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06872__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05589_ _02662_ _02663_ net467 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__o21a_1
X_07328_ _03763_ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07259_ _03901_ _03929_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nand2_1
XANTENNA__07821__A1 top.findLeastValue.sum\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ net723 net558 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__and2_1
XANTENNA__09594__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _02404_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_2
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_2
Xfanout462 net466 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_4
Xfanout495 top.cb_syn.end_cnt\[2\] vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11724_ clknet_leaf_74_clk _02274_ _01114_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ clknet_leaf_114_clk _02205_ _01045_ vssd1 vssd1 vccd1 vccd1 top.path\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11586_ clknet_leaf_30_clk _02151_ _00976_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10606_ net743 net578 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10537_ net819 net654 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__and2_1
X_10468_ net829 net664 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10399_ net801 net636 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07879__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06000__A0 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ _02434_ top.findLeastValue.val1\[15\] _02494_ top.compVal\[14\] vssd1 vssd1
+ vccd1 vccd1 _03428_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_48_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06561_ _03325_ _03363_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and2b_1
X_08300_ top.cb_syn.char_path_n\[54\] net193 _04712_ vssd1 vssd1 vccd1 vccd1 _01673_
+ sky130_fd_sc_hd__o21a_1
X_05512_ net447 net526 _02596_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a21o_1
X_09280_ net343 _04063_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[11\] sky130_fd_sc_hd__and2_1
X_06492_ _02454_ _03321_ _03323_ top.histogram.total\[0\] top.histogram.total\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__o2111a_2
X_08231_ top.cb_syn.char_path_n\[89\] net373 net327 top.cb_syn.char_path_n\[87\] net176
+ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a221o_1
X_05443_ net470 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06854__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08162_ top.cb_syn.char_path_n\[123\] net191 _04643_ vssd1 vssd1 vccd1 vccd1 _01742_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05374_ top.findLeastValue.val1\[26\] vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__inv_2
X_08093_ top.cb_syn.num_lefts\[5\] top.cb_syn.num_lefts\[4\] top.cb_syn.num_lefts\[3\]
+ _04592_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__and4_1
XANTENNA__07803__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07113_ top.findLeastValue.val2\[23\] top.findLeastValue.val1\[23\] _03787_ _03788_
+ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a211o_1
XANTENNA__07927__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09005__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_A _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ _02455_ _02480_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__nor2_1
XANTENNA__08359__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Left_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08995_ top.WB.CPU_DAT_O\[25\] net1344 net365 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XANTENNA__05447__A top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ top.hTree.tree_reg\[8\] top.findLeastValue.sum\[8\] net267 vssd1 vssd1 vccd1
+ vccd1 _04483_ sky130_fd_sc_hd__mux2_1
XANTENNA__05593__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__A top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ net475 _04426_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout652_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06828_ top.findLeastValue.val2\[40\] net129 net119 _03619_ vssd1 vssd1 vccd1 vccd1
+ _02048_ sky130_fd_sc_hd__o22a_1
X_09616_ net750 net585 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09547_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__and2_1
X_06759_ _02434_ top.findLeastValue.val2\[15\] top.findLeastValue.val2\[14\] vssd1
+ vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__a21oi_1
X_09478_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08429_ top.cb_syn.h_element\[55\] top.cb_syn.h_element\[46\] net517 vssd1 vssd1
+ vccd1 vccd1 _04780_ sky130_fd_sc_hd__mux2_1
X_11947__910 vssd1 vssd1 vccd1 vccd1 _11947__910/HI net910 sky130_fd_sc_hd__conb_1
X_11440_ clknet_leaf_93_clk _02005_ _00830_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_11371_ clknet_leaf_16_clk _01936_ _00761_ vssd1 vssd1 vccd1 vccd1 top.cw1\[3\] sky130_fd_sc_hd__dfrtp_1
X_10322_ net730 net565 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__and2_1
X_10184_ net801 net636 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__and2_1
XANTENNA__09771__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout292 net295 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05584__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06887__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 net273 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ clknet_leaf_80_clk _02257_ _01097_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06836__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11638_ clknet_leaf_100_clk _02188_ _01028_ vssd1 vssd1 vccd1 vccd1 top.path\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ clknet_leaf_23_clk _02134_ _00959_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
Xhold718 top.findLeastValue.sum\[25\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold707 top.histogram.state\[3\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold729 top.findLeastValue.sum\[21\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08746__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ top.hTree.tree_reg\[37\] top.findLeastValue.sum\[37\] net283 vssd1 vssd1
+ vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
X_08780_ _02546_ _04963_ _04966_ _04968_ top.translation.index\[6\] vssd1 vssd1 vccd1
+ vccd1 _04969_ sky130_fd_sc_hd__a311o_1
XANTENNA__05575__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ top.hTree.tree_reg\[50\] top.findLeastValue.least2\[4\] net280 vssd1 vssd1
+ vccd1 vccd1 _04310_ sky130_fd_sc_hd__mux2_1
X_05992_ top.WB.CPU_DAT_O\[9\] net1332 net347 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07662_ top.hTree.write_HT_fin _02837_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__nor2_2
X_07593_ net550 _04175_ _04189_ _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_88_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ net401 _04267_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nand2_1
X_06613_ _03403_ _03405_ _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__or3_2
X_09332_ net974 net226 net218 _04447_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06544_ net1519 _03356_ _03332_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08517__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ _05207_ _05221_ _05222_ _05208_ net1708 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[6\]
+ sky130_fd_sc_hd__a32o_1
X_06475_ net297 _03248_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__nor2_1
X_09194_ top.cb_syn.char_path_n\[1\] _04201_ _04563_ net463 vssd1 vssd1 vccd1 vccd1
+ _05179_ sky130_fd_sc_hd__o211a_1
X_08214_ top.cb_syn.char_path_n\[97\] net195 _04669_ vssd1 vssd1 vccd1 vccd1 _01716_
+ sky130_fd_sc_hd__o21a_1
X_05426_ net516 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__inv_2
X_08145_ net172 _04633_ _04634_ _04628_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05357_ top.findLeastValue.val2\[10\] vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__inv_2
XANTENNA__05876__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ _02531_ _04567_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05288_ net715 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ top.findLeastValue.val1\[10\] top.findLeastValue.val1\[9\] top.findLeastValue.val1\[8\]
+ top.findLeastValue.val1\[7\] vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold12 top.sram_interface.init_counter\[14\] vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 top.hTree.node_reg\[17\] vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__B net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08978_ top.WB.CPU_DAT_O\[23\] top.cb_syn.h_element\[55\] net368 vssd1 vssd1 vccd1
+ vccd1 _01360_ sky130_fd_sc_hd__mux2_1
Xhold34 top.hTree.tree_reg\[51\] vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05566__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold56 top.hTree.node_reg\[39\] vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 top.hTree.node_reg\[7\] vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 top.hTree.node_reg\[60\] vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ net437 net1433 net252 top.findLeastValue.sum\[12\] _04469_ vssd1 vssd1 vccd1
+ vccd1 _01801_ sky130_fd_sc_hd__a221o_1
Xhold89 top.sram_interface.word_cnt\[11\] vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 net60 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ clknet_leaf_52_clk _01505_ _00330_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07712__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ clknet_leaf_27_clk _01456_ _00261_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_42_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06455__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06818__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09217__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11423_ clknet_leaf_103_clk _01988_ _00813_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[27\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_9 _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ clknet_leaf_100_clk _01919_ _00744_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_10305_ net841 net676 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__and2_1
X_11285_ clknet_leaf_44_clk _01850_ _00675_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_10236_ net799 net634 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__and2_1
XANTENNA__05557__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10167_ net820 net655 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__and2_1
X_10098_ net830 net665 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06260_ top.TRN_char_index\[4\] _03050_ _02591_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06191_ top.TRN_char_index\[6\] _03057_ _02585_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a21oi_1
Xhold504 top.cb_syn.curr_index\[3\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 net85 vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 net58 vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__and2_1
Xhold537 top.hTree.node_reg\[46\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 top.hTree.tree_reg\[46\] vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 top.cb_syn.curr_index\[7\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
X_08901_ net1240 top.WB.CPU_DAT_O\[1\] net306 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ net858 net693 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__and2_1
XANTENNA__08800__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05548__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ top.translation.index\[6\] _05019_ _05020_ top.translation.index\[4\] vssd1
+ vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a31o_1
X_05975_ top.WB.CPU_DAT_O\[26\] net1283 net345 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
X_08763_ top.path\[93\] net323 _04951_ net425 net504 vssd1 vssd1 vccd1 vccd1 _04952_
+ sky130_fd_sc_hd__o221a_1
X_07714_ _04257_ _04295_ _04296_ net1619 net449 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__o32a_1
X_08694_ _02566_ top.header_synthesis.start _03389_ vssd1 vssd1 vccd1 vccd1 _04895_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout448_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05720__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ _02551_ _04175_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__or2_4
X_09315_ net1002 net224 net215 _04515_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__a22o_1
X_06527_ net1643 _03336_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__nor2_1
X_09246_ _05207_ _05209_ _05210_ _05208_ net1713 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[1\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout615_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06458_ _03249_ _03252_ _03302_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05409_ top.cb_syn.zeroes\[7\] vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06389_ top.hist_data_o\[13\] top.hist_data_o\[12\] vssd1 vssd1 vccd1 vccd1 _03254_
+ sky130_fd_sc_hd__and2_1
X_09177_ net1511 _05054_ _05090_ top.hTree.state\[6\] vssd1 vssd1 vccd1 vccd1 _00025_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__05484__B2 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ top.cb_syn.cb_length\[4\] _04618_ _04621_ net172 vssd1 vssd1 vccd1 vccd1
+ _04622_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08059_ _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11070_ clknet_leaf_57_clk _01635_ _00460_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XANTENNA__06984__A1 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
X_10021_ net830 net665 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__and2_1
XANTENNA__09383__C1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05539__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ clknet_leaf_71_clk _01488_ _00313_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10854_ clknet_leaf_116_clk _01448_ _00244_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05711__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10785_ clknet_leaf_114_clk _01391_ _00175_ vssd1 vssd1 vccd1 vccd1 top.path\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05475__B2 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11406_ clknet_leaf_87_clk _01971_ _00796_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[10\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_74_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11337_ clknet_leaf_84_clk _01902_ _00727_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11268_ clknet_leaf_69_clk net1451 _00658_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_11199_ clknet_leaf_29_clk _01764_ _00589_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_118_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10219_ net807 net642 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__and2_1
XANTENNA__07924__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05760_ net544 net536 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05691_ top.cb_syn.char_path\[38\] net529 net310 top.cb_syn.char_path\[102\] vssd1
+ vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05702__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07430_ top.dut.bits_in_buf\[3\] _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07361_ _03801_ _03802_ _03999_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a21o_1
XANTENNA__09687__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06312_ _03170_ _03173_ _03176_ _03181_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__or4_1
X_09100_ _05119_ _05120_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__or2_1
XANTENNA__08591__A _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07292_ top.findLeastValue.sum\[32\] net276 _03953_ _03954_ vssd1 vssd1 vccd1 vccd1
+ _01919_ sky130_fd_sc_hd__a22o_1
X_09031_ top.WB.CPU_DAT_O\[19\] net1202 net313 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06243_ net458 _03095_ _03101_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05466__B2 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 top.hTree.node_reg\[18\] vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
X_06174_ net445 top.TRN_char_index\[1\] vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nand2_1
XANTENNA__10345__B net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold334 net100 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 net84 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 top.path\[113\] vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 top.cb_syn.char_path\[95\] vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 net75 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05769__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 top.path\[54\] vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top.hTree.tree_reg\[4\] vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09933_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__and2_1
XANTENNA__08530__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 top.hTree.nulls\[56\] vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout814 net816 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout803 net808 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_2
Xfanout825 net826 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_2
X_09864_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__and2_1
Xfanout847 net854 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout836 net845 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 net876 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__dlymetal6s2s_1
X_08815_ top.path\[108\] top.path\[109\] top.path\[110\] top.path\[111\] net511 net507
+ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__mux4_1
X_09795_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07391__B2 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05958_ top.compVal\[3\] net160 net143 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ _02220_ sky130_fd_sc_hd__a22o_1
X_08746_ top.path\[116\] net403 net323 top.path\[117\] net505 vssd1 vssd1 vccd1 vccd1
+ _04935_ sky130_fd_sc_hd__o221a_1
XANTENNA__05941__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _04884_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__and2_1
X_05889_ top.hist_data_o\[9\] top.WB.CPU_DAT_O\[9\] net352 vssd1 vssd1 vccd1 vccd1
+ _02261_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout732_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ top.cb_syn.h_element\[58\] top.cb_syn.h_element\[49\] _04176_ vssd1 vssd1
+ vccd1 vccd1 _04225_ sky130_fd_sc_hd__mux2_1
XANTENNA__08891__A1 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07559_ top.cb_syn.char_path_n\[46\] top.cb_syn.char_path_n\[45\] top.cb_syn.char_path_n\[48\]
+ top.cb_syn.char_path_n\[47\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ net839 net674 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ top.header_synthesis.header\[3\] top.cb_syn.char_index\[3\] net490 vssd1
+ vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05457__B2 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08440__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ clknet_leaf_71_clk _01687_ _00512_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[68\]
+ sky130_fd_sc_hd__dfrtp_1
X_11053_ clknet_leaf_25_clk _01618_ _00443_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10271__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ net840 net675 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__and2_1
XANTENNA__06895__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05932__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10906_ clknet_leaf_33_clk _01478_ _00296_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08882__A1 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11886_ net441 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10837_ clknet_leaf_115_clk _01431_ _00227_ vssd1 vssd1 vccd1 vccd1 top.path\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08634__A1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ clknet_leaf_111_clk _01374_ _00158_ vssd1 vssd1 vccd1 vccd1 top.path\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10699_ clknet_leaf_21_clk _01330_ _00089_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_57_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06930_ top.findLeastValue.val1\[27\] net134 net115 top.compVal\[27\] vssd1 vssd1
+ vccd1 vccd1 _01988_ sky130_fd_sc_hd__o22a_1
X_08600_ _04818_ _04819_ _02542_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__mux2_1
X_06861_ top.compVal\[23\] top.findLeastValue.val1\[23\] net156 vssd1 vssd1 vccd1
+ vccd1 _03636_ sky130_fd_sc_hd__mux2_1
X_05812_ top.findLeastValue.least2\[6\] top.findLeastValue.least2\[5\] top.findLeastValue.least2\[4\]
+ top.findLeastValue.least2\[7\] vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_66_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09580_ net798 net633 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__and2_1
X_06792_ _02430_ top.findLeastValue.val2\[22\] _03576_ vssd1 vssd1 vccd1 vccd1 _03590_
+ sky130_fd_sc_hd__or3b_1
X_08531_ net1068 top.cb_syn.char_path_n\[28\] net234 vssd1 vssd1 vccd1 vccd1 _01511_
+ sky130_fd_sc_hd__mux2_1
X_05743_ top.findLeastValue.histo_index\[8\] top.findLeastValue.histo_index\[7\] vssd1
+ vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_38_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05674_ _02733_ _02734_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__or2_1
X_08462_ net1320 top.cb_syn.char_path_n\[97\] net237 vssd1 vssd1 vccd1 vccd1 _01580_
+ sky130_fd_sc_hd__mux2_1
X_07413_ top.findLeastValue.histo_index\[2\] top.findLeastValue.least1\[2\] net148
+ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08873__A1 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ top.cb_syn.char_path_n\[8\] net376 net333 top.cb_syn.char_path_n\[6\] net179
+ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06884__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07344_ net268 _03992_ _03993_ net275 net1630 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_98_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07275_ net270 _03941_ _03942_ net276 net1696 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a32o_1
X_06226_ top.hist_addr\[5\] top.hist_addr\[4\] _03098_ vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__and3_1
X_09014_ net1612 _05081_ _05082_ top.TRN_char_index\[3\] vssd1 vssd1 vccd1 vccd1 _01329_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout313_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 top.cb_syn.char_path\[92\] vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 top.cb_syn.char_path\[16\] vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 top.cb_syn.char_path\[53\] vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net49 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
X_06157_ _03025_ _03031_ _02877_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06088_ _02987_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__inv_2
Xhold186 _01535_ vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 top.cb_syn.char_path\[105\] vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 top.histogram.sram_out\[25\] vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07665__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_2
X_09916_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__and2_1
Xfanout622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_2
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_1
Xfanout633 net638 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_1
Xhold197 top.path\[4\] vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10091__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net661 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_2
Xfanout666 net669 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_2
Xfanout644 net647 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_2
Xfanout688 net689 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_2
X_09847_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__and2_1
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_2
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_2
X_09778_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08729_ top.path\[56\] top.path\[57\] top.path\[58\] top.path\[59\] net508 net506
+ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_107_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ clknet_leaf_106_clk _02290_ _01130_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11671_ clknet_leaf_91_clk _02221_ _01061_ vssd1 vssd1 vccd1 vccd1 top.compVal\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07419__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10622_ clknet_leaf_83_clk _01253_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ net832 net667 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__and2_1
X_10484_ net837 net672 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ clknet_leaf_56_clk _01670_ _00495_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[51\]
+ sky130_fd_sc_hd__dfrtp_2
X_11036_ clknet_leaf_49_clk _01601_ _00426_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08837__C top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11938_ net901 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_82_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06866__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ clknet_leaf_113_clk _02402_ _01241_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_15_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05390_ top.cw2\[5\] vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07060_ _03727_ _03730_ _03728_ _03725_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a211o_1
X_06011_ net481 top.controller.state_reg\[4\] _02878_ vssd1 vssd1 vccd1 vccd1 _02924_
+ sky130_fd_sc_hd__and3_2
XANTENNA__07291__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__and2_1
X_07962_ net477 _04494_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__or2_1
X_07893_ net421 _04439_ _04440_ net263 vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__o211a_1
XANTENNA__09335__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ top.findLeastValue.val1\[44\] net136 net113 net1753 vssd1 vssd1 vccd1 vccd1
+ _02005_ sky130_fd_sc_hd__o22a_1
X_09632_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__and2_1
X_06844_ top.findLeastValue.val2\[32\] net127 net118 _03627_ vssd1 vssd1 vccd1 vccd1
+ _02040_ sky130_fd_sc_hd__o22a_1
X_09563_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__and2_1
XANTENNA__09099__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ net1255 top.cb_syn.char_path_n\[45\] net244 vssd1 vssd1 vccd1 vccd1 _01528_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout263_A _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06775_ _02421_ top.findLeastValue.val2\[31\] top.findLeastValue.val2\[30\] _02422_
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a22oi_1
X_05726_ top.cb_syn.char_path\[0\] net546 net538 top.cb_syn.char_path\[64\] vssd1
+ vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a22o_1
X_09494_ net780 net615 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__and2_1
XANTENNA__06306__C1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net1277 top.cb_syn.char_path_n\[114\] net242 vssd1 vssd1 vccd1 vccd1 _01597_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05657_ top.hTree.node_reg\[44\] net307 _02720_ net467 vssd1 vssd1 vccd1 vccd1 _02721_
+ sky130_fd_sc_hd__a22o_1
X_08376_ top.cb_syn.char_path_n\[16\] net205 _04750_ vssd1 vssd1 vccd1 vccd1 _01635_
+ sky130_fd_sc_hd__o21a_1
X_05588_ top.cb_syn.char_path\[55\] net530 net311 top.cb_syn.char_path\[119\] vssd1
+ vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_83_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05879__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07327_ _03766_ _03980_ _03764_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07258_ _03901_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06209_ top.cw2\[7\] _02600_ _03081_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__a31o_1
X_07189_ _03789_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__B net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05596__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _02548_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_2
Xfanout441 net72 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
Xfanout463 net465 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout452 top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
Xfanout496 top.cb_syn.end_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
Xfanout485 top.findLeastValue.histo_index\[4\] vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11723_ clknet_leaf_74_clk _02273_ _01113_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06848__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ clknet_leaf_115_clk _02204_ _01044_ vssd1 vssd1 vccd1 vccd1 top.path\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_10605_ net743 net578 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ clknet_leaf_30_clk _02150_ _00975_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10536_ net817 net652 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ net829 net664 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__and2_1
X_10398_ net801 net636 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__and2_1
XANTENNA__05587__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ clknet_leaf_64_clk _01584_ _00409_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08620__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06560_ top.histogram.total\[0\] _03322_ _03323_ top.histogram.total\[1\] vssd1 vssd1
+ vccd1 vccd1 _03363_ sky130_fd_sc_hd__a31o_1
X_05511_ net447 top.WorR net533 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__and3_1
X_06491_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__and2_1
X_08230_ net1746 net194 _04677_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__o21a_1
X_05442_ top.cb_syn.zero_count\[5\] vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__inv_2
X_08161_ top.cb_syn.char_path_n\[124\] net369 net326 top.cb_syn.char_path_n\[122\]
+ net173 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a221o_1
X_05373_ top.findLeastValue.val1\[27\] vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__inv_2
X_08092_ top.cb_syn.num_lefts\[3\] _04592_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__nand2_1
X_07112_ top.findLeastValue.val2\[23\] top.findLeastValue.val1\[23\] top.findLeastValue.val1\[22\]
+ top.findLeastValue.val2\[22\] vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07043_ _03394_ _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__and2_1
XANTENNA__08213__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05578__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ top.WB.CPU_DAT_O\[26\] net1192 net365 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout380_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ top.hTree.tree_reg\[8\] top.findLeastValue.sum\[8\] net285 vssd1 vssd1 vccd1
+ vccd1 _04482_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout478_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ top.hTree.tree_reg\[22\] top.findLeastValue.sum\[22\] net265 vssd1 vssd1
+ vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
X_09615_ net733 net568 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__and2_1
X_06827_ top.compVal\[40\] top.findLeastValue.val1\[40\] net153 vssd1 vssd1 vccd1
+ vccd1 _03619_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09546_ net737 net572 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__and2_1
XANTENNA__08774__A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06758_ _03551_ _03555_ _03550_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08819__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05709_ top.cb_syn.char_path\[35\] net529 net310 top.cb_syn.char_path\[99\] vssd1
+ vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a22o_1
X_09477_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout812_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08428_ top.cb_syn.char_index\[1\] _04779_ _04772_ vssd1 vssd1 vccd1 vccd1 _01612_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06689_ top.compVal\[44\] _02480_ _03485_ _03486_ vssd1 vssd1 vccd1 vccd1 _03487_
+ sky130_fd_sc_hd__o211a_1
X_08359_ top.cb_syn.char_path_n\[25\] net374 net330 top.cb_syn.char_path_n\[23\] net177
+ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ clknet_leaf_15_clk _01935_ _00760_ vssd1 vssd1 vccd1 vccd1 top.cw1\[2\] sky130_fd_sc_hd__dfrtp_1
X_10321_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__and2_1
X_11908__939 vssd1 vssd1 vccd1 vccd1 net939 _11908__939/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_115_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10252_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__and2_1
XANTENNA__05569__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ net802 net637 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__and2_1
XANTENNA_input39_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06230__A1 top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 _04249_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
Xfanout260 _04256_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_4
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06469__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07730__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ clknet_leaf_80_clk _02256_ _01096_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ clknet_leaf_98_clk _02187_ _01027_ vssd1 vssd1 vccd1 vccd1 top.path\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_11568_ clknet_leaf_7_clk _02133_ _00958_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold719 top.hTree.nullSumIndex\[5\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08994__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold708 top.findLeastValue.sum\[28\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ net733 net568 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11499_ clknet_leaf_0_clk _02064_ _00889_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10454__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08746__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08859__A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ net257 _04308_ _04309_ net985 net433 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a32o_1
X_05991_ top.WB.CPU_DAT_O\[10\] net1059 net348 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XANTENNA__05980__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ net471 _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__nand2_1
X_07592_ top.cb_syn.h_element\[54\] _04190_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ net975 net220 _05279_ _05280_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06612_ _03400_ _03407_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__or3_1
X_09331_ net1028 net226 net218 _04451_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__a22o_1
X_06543_ top.histogram.total\[10\] top.histogram.total\[9\] _03331_ vssd1 vssd1 vccd1
+ vccd1 _03356_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ top.cb_syn.zero_count\[6\] _05218_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06474_ top.hist_data_o\[4\] _03246_ top.hist_data_o\[5\] vssd1 vssd1 vccd1 vccd1
+ _03313_ sky130_fd_sc_hd__a21o_1
X_05425_ net496 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__inv_2
X_09193_ _04542_ _04543_ _05178_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21o_1
X_08213_ top.cb_syn.char_path_n\[98\] net372 net329 top.cb_syn.char_path_n\[96\] net177
+ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a221o_1
XANTENNA__07003__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _04200_ _04629_ _04632_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08533__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05356_ top.findLeastValue.val2\[13\] vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__inv_2
XANTENNA__08985__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08075_ _04570_ _04576_ _04581_ _04566_ net1722 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a32o_1
X_05287_ net441 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07026_ _03691_ _03696_ _03701_ _02562_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__a31o_1
Xhold13 top.hTree.node_reg\[27\] vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06212__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08977_ top.WB.CPU_DAT_O\[24\] net1780 net367 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout762_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 top.hTree.tree_reg\[48\] vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 top.hTree.node_reg\[26\] vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 top.hTree.node_reg\[59\] vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A1 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold68 top.hTree.node_reg\[56\] vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 top.hTree.node_reg\[51\] vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ net420 _04467_ _04468_ net263 vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__o211a_1
Xhold57 top.hTree.node_reg\[41\] vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05971__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ net432 net1546 net253 top.findLeastValue.sum\[26\] _04413_ vssd1 vssd1 vccd1
+ vccd1 _01815_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ clknet_leaf_27_clk _01455_ _00260_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_3_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05723__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ net801 net636 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11422_ clknet_leaf_103_clk _01987_ _00812_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[26\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__08976__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ clknet_leaf_106_clk _01918_ _00743_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10304_ net844 net679 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__and2_1
X_11284_ clknet_leaf_42_clk _01849_ _00674_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ net800 net635 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__and2_1
XANTENNA__07400__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10166_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__and2_1
X_10097_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__and2_1
XANTENNA__09153__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07522__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05714__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ clknet_leaf_54_clk net1246 _00389_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11889__920 vssd1 vssd1 vccd1 vccd1 net920 _11889__920/LO sky130_fd_sc_hd__conb_1
XFILLER_0_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07562__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06190_ top.cb_syn.char_index\[6\] _03047_ _03063_ vssd1 vssd1 vccd1 vccd1 _03064_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08967__A0 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold516 top.histogram.sram_out\[8\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 top.histogram.total\[12\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold505 top.histogram.total\[23\] vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 top.cb_syn.curr_index\[4\] vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold538 top.sram_interface.zero_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
X_09880_ net858 net693 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__and2_1
X_08900_ net1187 top.WB.CPU_DAT_O\[2\] net305 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08831_ net430 _04985_ _04988_ _04993_ _02546_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__o311ai_1
X_05974_ top.WB.CPU_DAT_O\[27\] net1185 net345 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
X_08762_ top.path\[94\] top.path\[95\] net511 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__mux2_1
XANTENNA__05953__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ net515 _04208_ _04562_ _04894_ net1572 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a32o_1
X_07713_ top.hTree.tree_reg\[54\] net282 net417 vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o21a_1
XANTENNA__09144__B1 top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07644_ top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\] vssd1 vssd1 vccd1 vccd1
+ _04239_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05705__B1 _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _04143_ _04174_ _04107_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__mux2_1
X_09314_ _02851_ net220 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06526_ _03338_ _03349_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__nor2_1
X_09245_ top.cb_syn.zero_count\[0\] top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1 vccd1
+ _05210_ sky130_fd_sc_hd__or2_1
X_06457_ top.hist_data_o\[11\] _03251_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout510_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05408_ net1675 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout608_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06572__A top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06388_ top.hist_data_o\[12\] _03249_ _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__A0 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ _02567_ _02572_ _02618_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__o21ai_1
X_08127_ _02534_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05339_ top.findLeastValue.val2\[42\] vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__inv_2
X_08058_ _02530_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07009_ top.cw1\[1\] net140 _03686_ net487 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XANTENNA__09383__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ net830 net665 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05944__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ clknet_leaf_71_clk _01487_ _00312_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08438__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10853_ clknet_leaf_116_clk _01447_ _00243_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10269__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ clknet_leaf_117_clk _01390_ _00174_ vssd1 vssd1 vccd1 vccd1 top.path\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07544__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05475__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__S0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08949__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ clknet_leaf_87_clk _01970_ _00795_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[9\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_74_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11336_ clknet_leaf_81_clk _01901_ _00726_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11267_ clknet_leaf_68_clk _01832_ _00657_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_11198_ clknet_leaf_32_clk _01763_ _00588_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.left
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07924__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ net807 net642 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07924__B2 net1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__and2_1
XANTENNA__05935__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05690_ top.cb_syn.char_path\[6\] net549 net541 top.cb_syn.char_path\[70\] vssd1
+ vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07360_ top.findLeastValue.sum\[14\] net278 net272 _04004_ vssd1 vssd1 vccd1 vccd1
+ _01901_ sky130_fd_sc_hd__a22o_1
X_11932__895 vssd1 vssd1 vccd1 vccd1 _11932__895/HI net895 sky130_fd_sc_hd__conb_1
XANTENNA__07535__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06311_ top.cb_syn.curr_index\[4\] _02584_ _03180_ net446 _03179_ vssd1 vssd1 vccd1
+ vccd1 _03181_ sky130_fd_sc_hd__a221o_1
XANTENNA__09687__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07291_ _03874_ _03888_ net270 vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o21a_1
X_09030_ top.WB.CPU_DAT_O\[20\] net1382 net313 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
X_06242_ _03109_ _03111_ _03113_ _03114_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__or4_1
XANTENNA__08404__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06173_ _02536_ _02605_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__or3b_1
Xhold302 top.path\[77\] vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold313 top.cb_syn.char_path\[82\] vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 top.hTree.node_reg\[49\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold335 top.path\[110\] vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09932_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__and2_1
Xhold346 top.cb_syn.char_path\[31\] vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 top.cb_syn.char_path\[40\] vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 top.path\[9\] vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold379 _01578_ vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_2
Xfanout804 net808 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net854 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_2
X_09863_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__and2_1
Xfanout837 net845 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout826 net835 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_2
X_09794_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__and2_1
Xfanout859 net865 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_2
X_08814_ top.path\[32\] net405 net325 top.path\[33\] net430 vssd1 vssd1 vccd1 vccd1
+ _05003_ sky130_fd_sc_hd__o221a_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07391__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08745_ net428 _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout460_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05957_ top.compVal\[4\] net160 net143 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ _02221_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout558_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ top.cb_syn.curr_state\[2\] _04878_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__nor2_1
X_05888_ net1634 top.WB.CPU_DAT_O\[10\] net349 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
X_07627_ net1550 _04224_ _04212_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ _04150_ _04157_ _04109_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08782__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06509_ top.histogram.total\[29\] top.histogram.total\[28\] _03341_ vssd1 vssd1 vccd1
+ vccd1 _03342_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07489_ _04082_ _04091_ net342 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ net1081 _05200_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[2\]
+ sky130_fd_sc_hd__mux2_1
X_09159_ top.cb_syn.pulse_first net424 _02890_ net522 vssd1 vssd1 vccd1 vccd1 _05161_
+ sky130_fd_sc_hd__o31a_1
X_11121_ clknet_leaf_63_clk _01686_ _00511_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06957__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ clknet_leaf_24_clk _01617_ _00442_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_10003_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__and2_1
XANTENNA__06709__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ net917 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_103_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10905_ clknet_leaf_37_clk _01477_ _00295_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_11885_ net441 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05696__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836_ clknet_leaf_115_clk _01430_ _00226_ vssd1 vssd1 vccd1 vccd1 top.path\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07517__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07800__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ clknet_leaf_110_clk _01373_ _00157_ vssd1 vssd1 vccd1 vccd1 top.path\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09292__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10698_ clknet_leaf_7_clk net1613 _00088_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ clknet_leaf_43_clk _01884_ _00709_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05620__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ top.findLeastValue.val2\[24\] net132 net122 _03635_ vssd1 vssd1 vccd1 vccd1
+ _02032_ sky130_fd_sc_hd__o22a_1
X_05811_ top.findLeastValue.least2\[3\] top.findLeastValue.least2\[2\] top.findLeastValue.least2\[1\]
+ top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__or4_1
XANTENNA__05990__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ _03564_ _03588_ _03580_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a21bo_1
X_08530_ net1426 top.cb_syn.char_path_n\[29\] net234 vssd1 vssd1 vccd1 vccd1 _01512_
+ sky130_fd_sc_hd__mux2_1
X_05742_ top.findLeastValue.histo_index\[8\] top.findLeastValue.histo_index\[7\] vssd1
+ vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05673_ top.cb_syn.char_path\[41\] net529 net312 top.cb_syn.char_path\[105\] vssd1
+ vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
X_08461_ net1404 top.cb_syn.char_path_n\[98\] net232 vssd1 vssd1 vccd1 vccd1 _01581_
+ sky130_fd_sc_hd__mux2_1
X_07412_ _02518_ net126 net124 _04036_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_18_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05687__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ top.cb_syn.char_path_n\[8\] net201 _04758_ vssd1 vssd1 vccd1 vccd1 _01627_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07343_ _03769_ _03991_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_98_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07274_ _03729_ _03940_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__nand2_1
X_06225_ top.hist_addr\[2\] top.hist_addr\[1\] top.hist_addr\[0\] top.hist_addr\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a31o_1
X_09013_ net1758 _05081_ _05082_ top.TRN_char_index\[4\] vssd1 vssd1 vccd1 vccd1 _01330_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08389__B2 top.cb_syn.char_path_n\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 top.cb_syn.char_path\[112\] vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout306_A _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__S net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 _01536_ vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 top.cb_syn.char_path\[67\] vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 top.header_synthesis.header\[4\] vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ top.sram_interface.init_counter\[9\] _03024_ vssd1 vssd1 vccd1 vccd1 _03031_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06087_ _02985_ _02986_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__or2_1
XANTENNA__07665__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 top.histogram.total\[7\] vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 top.path\[29\] vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 top.compVal\[24\] vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05611__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 top.cb_syn.char_path\[113\] vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__and2_1
Xfanout623 net629 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_2
Xfanout612 net630 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_2
Xfanout601 net612 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09338__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 top.path\[34\] vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
X_09846_ net839 net674 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__and2_1
Xfanout634 net638 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_2
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10091__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 net647 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_1
Xfanout667 net668 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_2
Xfanout689 net712 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_2
X_09777_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__and2_1
X_06989_ _02506_ net125 net123 _03679_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_107_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ net425 net508 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_107_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ top.cb_syn.end_cnt\[3\] _04873_ _04871_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05678__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ clknet_leaf_91_clk _02220_ _01060_ vssd1 vssd1 vccd1 vccd1 top.compVal\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09401__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ clknet_leaf_83_clk _01252_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10547__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ net832 net667 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07824__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10483_ net840 net675 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ clknet_leaf_56_clk _01669_ _00494_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[50\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09329__B1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05602__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ clknet_leaf_49_clk net1273 _00425_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08552__A1 top.cb_syn.char_path_n\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ net900 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_82_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05669__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07530__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__S _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11868_ clknet_leaf_112_clk _02401_ _01240_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_11799_ clknet_leaf_7_clk _02332_ _01171_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_10819_ clknet_leaf_97_clk _01413_ _00209_ vssd1 vssd1 vccd1 vccd1 top.path\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10457__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06010_ net304 _02923_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_93_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ top.hTree.tree_reg\[5\] top.findLeastValue.sum\[5\] net266 vssd1 vssd1 vccd1
+ vccd1 _04495_ sky130_fd_sc_hd__mux2_1
X_09700_ net849 net684 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__and2_1
X_06912_ top.findLeastValue.val1\[45\] net137 net113 net1654 vssd1 vssd1 vccd1 vccd1
+ _02006_ sky130_fd_sc_hd__o22a_1
X_07892_ net478 _04438_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__or2_1
XANTENNA__07346__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06843_ top.compVal\[32\] top.findLeastValue.val1\[32\] net151 vssd1 vssd1 vccd1
+ vccd1 _03627_ sky130_fd_sc_hd__mux2_1
X_09562_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__and2_1
X_06774_ _02421_ top.findLeastValue.val2\[31\] top.findLeastValue.val2\[30\] _02422_
+ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__o22a_1
X_08513_ net1067 top.cb_syn.char_path_n\[46\] net244 vssd1 vssd1 vccd1 vccd1 _01529_
+ sky130_fd_sc_hd__mux2_1
X_05725_ net1274 net170 _02777_ net209 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__a22o_1
X_09493_ net780 net615 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__and2_1
XANTENNA__08536__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05656_ _02718_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__or2_1
X_08444_ net1133 top.cb_syn.char_path_n\[115\] net242 vssd1 vssd1 vccd1 vccd1 _01598_
+ sky130_fd_sc_hd__mux2_1
X_05587_ top.cb_syn.char_path\[23\] net548 net538 top.cb_syn.char_path\[87\] vssd1
+ vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__a22o_1
X_08375_ top.cb_syn.char_path_n\[17\] net385 net340 top.cb_syn.char_path_n\[15\] net188
+ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_102_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07326_ _03779_ _03979_ _03786_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07257_ _03895_ _03898_ _03897_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06208_ _02501_ net361 _03074_ _03075_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__a22o_1
X_07188_ _03855_ _03858_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__a21oi_1
X_06139_ net1032 net166 _03017_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a21o_1
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_2
Xfanout431 net434 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_2
Xfanout475 net480 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_2
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
X_09829_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__and2_1
Xfanout497 top.cb_syn.end_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
Xfanout486 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
XFILLER_0_68_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06997__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11722_ clknet_leaf_72_clk _02272_ _01112_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11653_ clknet_leaf_115_clk _02203_ _01043_ vssd1 vssd1 vccd1 vccd1 top.path\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_10604_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ clknet_leaf_30_clk _02149_ _00974_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535_ net817 net652 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__and2_1
X_10466_ net829 net664 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__and2_1
XANTENNA__05818__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__A1 top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ net801 net636 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07525__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ clknet_leaf_70_clk net1214 _00408_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08620__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08864__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05510_ net444 top.histogram.wr_r_en\[1\] _02594_ top.histogram.wr_r_en\[0\] vssd1
+ vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__or4b_1
X_06490_ top.histogram.eof_n top.histogram.state\[1\] net453 vssd1 vssd1 vccd1 vccd1
+ _03323_ sky130_fd_sc_hd__o21a_1
X_05441_ top.cb_syn.zero_count\[2\] vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__inv_2
X_08160_ net1785 net191 _04642_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07111_ _03785_ _03786_ _03767_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05372_ top.findLeastValue.val1\[32\] vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07042_ _03707_ _03712_ _03717_ _03702_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08993_ top.WB.CPU_DAT_O\[27\] net1164 net366 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07944_ net435 net1599 net251 top.findLeastValue.sum\[9\] _04481_ vssd1 vssd1 vccd1
+ vccd1 _01798_ sky130_fd_sc_hd__a221o_1
X_07875_ top.hTree.tree_reg\[22\] top.findLeastValue.sum\[22\] net281 vssd1 vssd1
+ vccd1 vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout373_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ top.findLeastValue.val2\[41\] net129 net119 _03618_ vssd1 vssd1 vccd1 vccd1
+ _02049_ sky130_fd_sc_hd__o22a_1
X_09614_ net726 net561 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09545_ net737 net572 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__and2_1
X_06757_ top.findLeastValue.val2\[12\] _03552_ top.compVal\[12\] vssd1 vssd1 vccd1
+ vccd1 _03555_ sky130_fd_sc_hd__and3b_1
X_05708_ top.cb_syn.char_path\[3\] net548 net539 top.cb_syn.char_path\[67\] vssd1
+ vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a22o_1
X_09476_ net785 net620 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout638_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06688_ _02408_ top.findLeastValue.val1\[43\] _03484_ vssd1 vssd1 vccd1 vccd1 _03486_
+ sky130_fd_sc_hd__a21oi_1
X_08427_ top.cb_syn.h_element\[56\] top.cb_syn.h_element\[47\] net517 vssd1 vssd1
+ vccd1 vccd1 _04779_ sky130_fd_sc_hd__mux2_1
X_05639_ top.hTree.node_reg\[47\] net355 _02704_ _02705_ vssd1 vssd1 vccd1 vccd1 _02706_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout805_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ net1781 net194 _04741_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ top.cb_syn.char_path_n\[60\] net371 net328 top.cb_syn.char_path_n\[58\] net175
+ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07309_ _03749_ _03762_ _03957_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__nand3_1
X_10320_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10251_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__and2_1
X_10182_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__and2_1
XANTENNA__10560__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 net253 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
Xfanout283 _04249_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_4
Xfanout261 _04256_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08030__A top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11705_ clknet_leaf_80_clk _02255_ _01095_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ clknet_leaf_97_clk _02186_ _01026_ vssd1 vssd1 vccd1 vccd1 top.path\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11567_ clknet_leaf_6_clk _02132_ _00957_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold709 top.cb_syn.num_lefts\[2\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10518_ net733 net568 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11498_ clknet_leaf_0_clk _02063_ _00888_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10449_ net813 net648 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05990_ top.WB.CPU_DAT_O\[11\] net1150 net348 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XANTENNA__06379__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ top.findLeastValue.least1\[8\] net390 net265 top.hTree.tree_reg\[63\] vssd1
+ vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__o22ai_1
X_07591_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06611_ top.compVal\[45\] top.compVal\[44\] _03406_ _03408_ vssd1 vssd1 vccd1 vccd1
+ _03409_ sky130_fd_sc_hd__or4_1
X_09330_ net1021 net226 net217 _04455_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06542_ net1478 _03332_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ top.cb_syn.zero_count\[6\] _05218_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08212_ top.cb_syn.char_path_n\[98\] net200 _04668_ vssd1 vssd1 vccd1 vccd1 _01717_
+ sky130_fd_sc_hd__o21a_1
X_06473_ net1376 net297 _03312_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a21o_1
X_05424_ top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__inv_2
X_09192_ net514 _02888_ net463 vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__mux2_1
XANTENNA__07003__B net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _04200_ _04629_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout121_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05355_ top.findLeastValue.val2\[14\] vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__inv_2
X_08074_ _02530_ _04568_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06996__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ _03697_ _03698_ _03699_ _03700_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 top.sram_interface.init_counter\[15\] vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08976_ top.WB.CPU_DAT_O\[25\] top.cb_syn.h_element\[57\] net367 vssd1 vssd1 vccd1
+ vccd1 _01362_ sky130_fd_sc_hd__mux2_1
Xhold47 top.hTree.node_reg\[21\] vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 top.hTree.node_reg\[22\] vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 top.hTree.node_reg\[35\] vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold58 top.hTree.tree_reg\[52\] vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ net478 _04466_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__or2_1
Xhold69 top.hTree.node_reg\[36\] vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ net422 _04411_ _04412_ net258 vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__o211a_1
X_07789_ net437 net1535 net251 top.findLeastValue.sum\[40\] _04357_ vssd1 vssd1 vccd1
+ vccd1 _01829_ sky130_fd_sc_hd__a221o_1
XANTENNA__07712__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06809_ _02406_ top.findLeastValue.val2\[45\] _03509_ _03606_ top.findLeastValue.val2\[46\]
+ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__06920__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ net797 net632 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ net731 net566 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__A1 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11421_ clknet_leaf_103_clk _01986_ _00811_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[25\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10555__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ clknet_leaf_103_clk _01917_ _00742_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10303_ net844 net679 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__and2_1
XANTENNA__06987__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11283_ clknet_leaf_44_clk _01848_ _00673_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_10234_ net800 net635 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__and2_1
X_10165_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05384__A top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__and2_1
XANTENNA__08361__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__A1 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09290__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ clknet_leaf_58_clk net1113 _00388_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06419__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07562__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ clknet_leaf_22_clk net1102 _01009_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold517 top.path\[92\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 top.hTree.tree_reg\[36\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap247 _04781_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
Xhold539 top.hTree.tree_reg\[30\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 top.histogram.state\[7\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08719__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ net503 _05008_ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__a21bo_1
X_08761_ top.path\[80\] top.path\[81\] top.path\[82\] top.path\[83\] net508 net506
+ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__mux4_1
X_05973_ top.WB.CPU_DAT_O\[28\] net1375 net346 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XANTENNA__05953__B2 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937__900 vssd1 vssd1 vccd1 vccd1 _11937__900/HI net900 sky130_fd_sc_hd__conb_1
X_08692_ _02543_ _04562_ _04208_ _04179_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__o211ai_1
X_07712_ top.findLeastValue.least2\[8\] net390 net265 top.hTree.tree_reg\[54\] net470
+ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__o221a_1
X_07643_ net518 top.cb_syn.h_element\[47\] net525 top.cb_syn.h_element\[56\] _04180_
+ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout169_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06902__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05705__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07574_ _04173_ _04158_ _04108_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09313_ _04257_ _05052_ _00053_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or3b_2
XANTENNA__08655__B1 _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06525_ net1532 _03337_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__nor2_1
X_09244_ top.cb_syn.zero_count\[0\] top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1 vccd1
+ _05209_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_60_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
X_06456_ net299 _03253_ _03300_ _03301_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__o31ai_1
X_05407_ top.WorR vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__inv_2
X_09175_ top.WB.curr_state\[1\] _02567_ top.WB.curr_state\[0\] _02617_ vssd1 vssd1
+ vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
X_08126_ _02535_ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__nand2_1
X_06387_ top.hist_data_o\[11\] top.hist_data_o\[10\] top.hist_data_o\[9\] top.hist_data_o\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__and4_1
X_05338_ top.findLeastValue.val2\[44\] vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08057_ _02531_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05641__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07008_ net1639 net140 _03686_ top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1
+ vccd1 _01935_ sky130_fd_sc_hd__a22o_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_12_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08186__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08959_ top.WB.CPU_DAT_O\[9\] net1453 net320 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__mux2_1
XANTENNA__05944__B2 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877__880 vssd1 vssd1 vccd1 vccd1 _11877__880/HI net880 sky130_fd_sc_hd__conb_1
X_10921_ clknet_leaf_71_clk _01486_ _00311_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10852_ clknet_leaf_116_clk _01446_ _00242_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10269__B net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10783_ clknet_leaf_117_clk _01389_ _00173_ vssd1 vssd1 vccd1 vccd1 top.path\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07544__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09297__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ clknet_leaf_87_clk _01969_ _00794_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[8\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11335_ clknet_leaf_84_clk _01900_ _00725_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11266_ clknet_leaf_82_clk _01831_ _00656_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09285__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__and2_1
X_11197_ clknet_leaf_26_clk _01762_ _00587_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10148_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__and2_1
X_10079_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__and2_1
XANTENNA__05935__B2 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05699__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07535__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06310_ top.cb_syn.max_index\[4\] _03102_ _03104_ top.hTree.nullSumIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__a22o_1
XANTENNA__05988__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07290_ _03874_ _03888_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__nand2_1
X_06241_ _02607_ _03036_ _03112_ _03107_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06172_ top.cb_syn.char_index\[5\] top.cb_syn.char_index\[4\] _03044_ vssd1 vssd1
+ vccd1 vccd1 _03047_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold325 _02301_ vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 top.path\[90\] vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 top.path\[87\] vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold336 top.cb_syn.char_path\[12\] vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__and2_1
Xhold358 top.cb_syn.char_path\[72\] vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 top.cb_syn.char_path\[97\] vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 top.cb_syn.char_path\[38\] vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08168__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout816 net877 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_2
Xfanout805 net808 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_1
Xfanout849 net854 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09862_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__and2_1
Xfanout838 net845 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07376__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout827 net835 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_2
X_09793_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__and2_1
X_08813_ net426 _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout286_A _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05956_ top.compVal\[5\] net160 net143 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ _02222_ sky130_fd_sc_hd__a22o_1
X_08744_ top.path\[118\] top.path\[119\] net512 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__mux2_1
XANTENNA__08539__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ top.cb_syn.curr_state\[2\] _04884_ _04879_ vssd1 vssd1 vccd1 vccd1 _04885_
+ sky130_fd_sc_hd__o21bai_1
X_05887_ net1534 top.WB.CPU_DAT_O\[11\] net349 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout453_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07626_ top.cb_syn.max_index\[5\] _04181_ _04221_ _04223_ vssd1 vssd1 vccd1 vccd1
+ _04224_ sky130_fd_sc_hd__o22a_1
XANTENNA__10089__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07557_ _04153_ _04156_ _04110_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_33_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout718_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06508_ top.histogram.total\[27\] top.histogram.total\[26\] _03340_ vssd1 vssd1 vccd1
+ vccd1 _03341_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07488_ _04086_ _04090_ net393 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ top.header_synthesis.header\[2\] top.cb_syn.char_index\[2\] net490 vssd1
+ vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__mux2_1
X_06439_ top.hist_data_o\[18\] _03271_ _03268_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09158_ top.cb_syn.char_path_n\[2\] net516 net463 _04562_ vssd1 vssd1 vccd1 vccd1
+ _05160_ sky130_fd_sc_hd__and4b_1
X_08109_ _04590_ _04591_ _04604_ _04589_ top.cb_syn.num_lefts\[1\] vssd1 vssd1 vccd1
+ vccd1 _01756_ sky130_fd_sc_hd__a32o_1
X_09089_ net455 top.sram_interface.word_cnt\[4\] _05100_ net1040 vssd1 vssd1 vccd1
+ vccd1 _00040_ sky130_fd_sc_hd__a22o_1
X_11120_ clknet_leaf_63_clk _01685_ _00510_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[66\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05614__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11051_ clknet_leaf_24_clk _01616_ _00441_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10002_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__and2_1
XANTENNA__06590__A1 top.header_synthesis.bit1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ net916 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10904_ clknet_leaf_51_clk _01476_ _00294_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_11884_ net441 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08619__A0 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10835_ clknet_leaf_116_clk _01429_ _00225_ vssd1 vssd1 vccd1 vccd1 top.path\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07517__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ clknet_leaf_111_clk _01372_ _00156_ vssd1 vssd1 vccd1 vccd1 top.path\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09292__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ clknet_leaf_6_clk _01328_ _00087_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09044__A0 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05605__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ clknet_leaf_41_clk _01883_ _00708_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06432__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11249_ clknet_leaf_74_clk net1566 _00639_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07358__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05810_ top.findLeastValue.least1\[8\] _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__nand2_1
X_06790_ _02431_ top.findLeastValue.val2\[20\] _03578_ vssd1 vssd1 vccd1 vccd1 _03588_
+ sky130_fd_sc_hd__or3b_1
X_05741_ top.findLeastValue.alternator_timer\[2\] _02784_ _02783_ top.findLeastValue.alternator_timer\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__a211o_1
X_05672_ top.cb_syn.char_path\[9\] net547 net540 top.cb_syn.char_path\[73\] vssd1
+ vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
X_08460_ net1302 top.cb_syn.char_path_n\[99\] net239 vssd1 vssd1 vccd1 vccd1 _01582_
+ sky130_fd_sc_hd__mux2_1
X_08391_ top.cb_syn.char_path_n\[9\] net381 net337 top.cb_syn.char_path_n\[7\] net184
+ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a221o_1
X_07411_ top.findLeastValue.histo_index\[3\] top.findLeastValue.least1\[3\] net150
+ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
X_07342_ _03769_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06884__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ _03729_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__or2_1
XANTENNA__07833__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06224_ top.hist_addr\[1\] top.hist_addr\[0\] vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__nand2_1
X_09012_ net1575 _05081_ _05082_ top.TRN_char_index\[5\] vssd1 vssd1 vccd1 vccd1 _01331_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09035__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06155_ net1525 net164 _03030_ net207 net157 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a221o_1
Xhold100 top.path\[53\] vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 top.hTree.tree_reg\[57\] vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 top.path\[10\] vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 top.path\[30\] vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 top.path\[108\] vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 top.cb_syn.char_path\[26\] vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06086_ top.cb_syn.i\[5\] top.cb_syn.cb_length\[5\] vssd1 vssd1 vccd1 vccd1 _02986_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold155 top.path\[19\] vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 top.path\[50\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout624 net629 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_2
Xhold188 top.cb_syn.char_path\[126\] vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_2
X_09914_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__and2_1
Xfanout613 net615 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_2
Xhold199 top.path\[43\] vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
X_09845_ net785 net620 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__and2_1
Xfanout646 net647 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_2
Xfanout635 net638 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_1
Xfanout657 net660 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_1
XANTENNA_fanout668_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_2
X_09776_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__and2_1
X_06988_ top.cw1\[6\] net148 _03662_ net482 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a22o_1
X_05939_ top.compVal\[22\] net158 net145 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 _02239_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout835_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08727_ top.sram_interface.TRN_counter\[0\] _04912_ _04916_ vssd1 vssd1 vccd1 vccd1
+ _01450_ sky130_fd_sc_hd__o21a_1
XANTENNA__09889__A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _04866_ net493 _04789_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__or3b_1
X_07609_ top.cb_syn.curr_state\[0\] _04181_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__nor2_1
XANTENNA__07901__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ top.cb_syn.end_cnt\[5\] _04800_ _04808_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or3_1
X_10620_ clknet_leaf_83_clk _01251_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10547__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07824__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__B2 top.findLeastValue.sum\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ net832 net667 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__and2_1
X_10482_ net840 net675 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__and2_1
XANTENNA__09026__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11103_ clknet_leaf_56_clk _01668_ _00493_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[49\]
+ sky130_fd_sc_hd__dfrtp_2
X_11034_ clknet_leaf_55_clk _01599_ _00424_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05807__D top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936_ net899 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__08304__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07811__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05523__C1 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ clknet_leaf_112_clk _02400_ _01239_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06427__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ clknet_leaf_97_clk _01412_ _00208_ vssd1 vssd1 vccd1 vccd1 top.path\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11798_ clknet_leaf_5_clk _02331_ _01170_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_10749_ clknet_leaf_10_clk _00044_ _00139_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07815__A1 top.findLeastValue.sum\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08776__C1 _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ top.hTree.tree_reg\[5\] top.findLeastValue.sum\[5\] net284 vssd1 vssd1 vccd1
+ vccd1 _04494_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_06911_ top.findLeastValue.val1\[46\] net142 _03393_ vssd1 vssd1 vccd1 vccd1 _02007_
+ sky130_fd_sc_hd__a21o_1
X_07891_ top.findLeastValue.sum\[19\] _04438_ net392 vssd1 vssd1 vccd1 vccd1 _04439_
+ sky130_fd_sc_hd__mux2_1
X_09630_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__and2_1
X_06842_ top.findLeastValue.val2\[33\] net127 net118 _03626_ vssd1 vssd1 vccd1 vccd1
+ _02041_ sky130_fd_sc_hd__o22a_1
X_09561_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__and2_1
X_06773_ top.compVal\[26\] _02467_ _03568_ _03569_ vssd1 vssd1 vccd1 vccd1 _03571_
+ sky130_fd_sc_hd__o211a_1
X_08512_ net1157 top.cb_syn.char_path_n\[47\] net242 vssd1 vssd1 vccd1 vccd1 _01530_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09099__A3 _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05724_ top.hTree.node_reg\[33\] net307 _02775_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_
+ sky130_fd_sc_hd__a211o_1
X_09492_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05655_ top.cb_syn.char_path\[12\] net547 net310 top.cb_syn.char_path\[108\] vssd1
+ vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
X_08443_ net1161 top.cb_syn.char_path_n\[116\] net242 vssd1 vssd1 vccd1 vccd1 _01599_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout249_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ net1751 net199 _04749_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__o21a_1
X_05586_ net89 net171 _02661_ net212 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07325_ _03776_ _03978_ _03783_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o21ai_1
X_07256_ net1735 net278 net272 _03928_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06207_ top.cw2\[6\] _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07676__B _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ _03767_ _03784_ _03860_ _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__or4_1
X_06138_ net1043 net166 net157 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a21o_1
X_06069_ top.cb_syn.count\[7\] _02526_ _02953_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__05596__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_2
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_4
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_2
Xfanout454 top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
X_09828_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__and2_1
Xfanout498 top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
Xfanout487 top.findLeastValue.histo_index\[1\] vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_2
Xfanout476 net480 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_2
X_09759_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10558__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ clknet_leaf_72_clk _02271_ _01111_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06848__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11652_ clknet_leaf_115_clk _02202_ _01042_ vssd1 vssd1 vccd1 vccd1 top.path\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_10603_ net743 net578 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ clknet_leaf_4_clk _02148_ _00973_ vssd1 vssd1 vccd1 vccd1 top.histogram.out_of_init
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10534_ net817 net652 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__and2_1
X_10465_ net828 net663 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10396_ net801 net636 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__and2_1
XANTENNA__05587__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07806__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ clknet_leaf_63_clk _01582_ _00407_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08637__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11919_ net950 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05440_ top.cb_syn.zero_count\[3\] vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05371_ top.findLeastValue.val1\[33\] vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__inv_2
X_07110_ _03777_ _03781_ _03779_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08090_ top.cb_syn.num_lefts\[2\] top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__and3_1
XANTENNA__08461__A1 top.cb_syn.char_path_n\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07041_ _03713_ _03714_ _03715_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__and4_1
XANTENNA__08213__B2 top.cb_syn.char_path_n\[96\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__A1 top.cb_syn.char_path_n\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08764__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ top.WB.CPU_DAT_O\[28\] net1249 net366 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__mux2_1
XANTENNA__05578__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07943_ net420 _04479_ _04480_ net260 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout199_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ net438 net1551 net248 net1806 _04425_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__a221o_1
X_06825_ top.compVal\[41\] top.findLeastValue.val1\[41\] net153 vssd1 vssd1 vccd1
+ vccd1 _03618_ sky130_fd_sc_hd__mux2_1
X_09613_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09544_ net737 net572 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__and2_1
X_06756_ _03550_ _03551_ _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nor3_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ net785 net620 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__and2_1
X_05707_ net1290 net170 _02762_ net212 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout533_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06687_ _02406_ top.findLeastValue.val1\[45\] top.findLeastValue.val1\[44\] _02407_
+ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__o22a_1
X_08426_ top.cb_syn.char_index\[2\] _04778_ _04772_ vssd1 vssd1 vccd1 vccd1 _01613_
+ sky130_fd_sc_hd__mux2_1
X_05638_ top.histogram.sram_out\[15\] net358 net409 top.hTree.node_reg\[15\] vssd1
+ vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05569_ top.cb_syn.char_path\[26\] net546 net537 top.cb_syn.char_path\[90\] vssd1
+ vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
X_08357_ top.cb_syn.char_path_n\[26\] net374 net330 top.cb_syn.char_path_n\[24\] net176
+ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout700_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ top.cb_syn.char_path_n\[60\] net192 _04706_ vssd1 vssd1 vccd1 vccd1 _01679_
+ sky130_fd_sc_hd__o21a_1
X_07308_ net268 _03966_ _03967_ net274 net1656 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a32o_1
X_07239_ _03895_ _03912_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a21boi_1
XANTENNA__05919__B _02898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05569__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__and2_1
XANTENNA__10560__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_2
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
Xfanout273 _03922_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
Xfanout295 _04112_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
Xfanout284 _04249_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_2
XANTENNA_hold745_A top.findLeastValue.sum\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954__917 vssd1 vssd1 vccd1 vccd1 _11954__917/HI net917 sky130_fd_sc_hd__conb_1
XFILLER_0_56_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ clknet_leaf_80_clk _02254_ _01094_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ clknet_leaf_98_clk _02185_ _01025_ vssd1 vssd1 vccd1 vccd1 top.path\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_11566_ clknet_leaf_5_clk _02131_ _00956_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
X_10517_ net755 net590 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__and2_1
X_11497_ clknet_leaf_119_clk _02062_ _00887_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08920__S _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10448_ net813 net648 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__and2_1
XANTENNA__06006__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379_ net769 net604 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07954__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06440__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07590_ top.cb_syn.pulse_first _02891_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or2_2
X_06610_ top.compVal\[35\] top.compVal\[34\] top.compVal\[33\] top.compVal\[32\] vssd1
+ vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06541_ _03333_ net1504 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nor2_1
X_09260_ _05207_ _05219_ _05220_ _05208_ net1642 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[5\]
+ sky130_fd_sc_hd__a32o_1
X_06472_ top.hist_data_o\[6\] _03248_ _03311_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__o21a_1
X_05423_ top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__inv_2
X_08211_ top.cb_syn.char_path_n\[99\] net380 net336 top.cb_syn.char_path_n\[97\] net183
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a221o_1
XANTENNA__07003__C net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09191_ net1604 _04257_ _05177_ _03393_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
X_08142_ _04611_ _04630_ _04631_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05354_ top.findLeastValue.val2\[16\] vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__inv_2
X_08073_ _04571_ _04576_ _04580_ _04566_ net1787 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06996__B2 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ top.findLeastValue.val2\[34\] top.findLeastValue.val2\[33\] top.findLeastValue.val2\[32\]
+ top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout114_A _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ top.WB.CPU_DAT_O\[26\] net1769 net367 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__mux2_1
Xhold15 top.sram_interface.init_counter\[12\] vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 top.hTree.node_reg\[62\] vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ top.findLeastValue.sum\[12\] _04466_ net392 vssd1 vssd1 vccd1 vccd1 _04467_
+ sky130_fd_sc_hd__mux2_1
Xhold26 top.controller.fin_FINISHED vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold48 top.hTree.node_reg\[61\] vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 top.hTree.tree_reg\[49\] vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ net475 _04410_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__or2_1
XANTENNA__08785__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07788_ net420 _04355_ _04356_ net262 vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__o211a_1
X_06808_ top.compVal\[40\] _02458_ _03514_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__o21bai_1
XANTENNA__05723__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05490__A top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06739_ top.findLeastValue.val2\[2\] _02444_ top.compVal\[3\] _02478_ vssd1 vssd1
+ vccd1 vccd1 _03537_ sky130_fd_sc_hd__a2bb2o_1
X_09527_ net747 net582 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__and2_1
X_11914__945 vssd1 vssd1 vccd1 vccd1 net945 _11914__945/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_42_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ net731 net566 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__and2_1
X_08409_ _02885_ _04606_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__nor2_1
X_09389_ net399 _04287_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ clknet_leaf_103_clk _01985_ _00810_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[24\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10555__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ clknet_leaf_106_clk _01916_ _00741_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10302_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__and2_1
X_11282_ clknet_leaf_44_clk _01847_ _00672_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10571__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ net803 net638 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__and2_1
XANTENNA__07400__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__and2_1
X_10095_ net833 net668 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05714__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06911__A1 top.findLeastValue.val1\[46\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10997_ clknet_leaf_58_clk _01562_ _00387_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05478__B2 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ clknet_leaf_22_clk _02168_ _01008_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11549_ clknet_leaf_47_clk _02114_ _00939_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold518 net104 vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold507 top.hTree.tree_reg\[0\] vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold529 _00035_ vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08719__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08760_ top.path\[84\] net402 net323 top.path\[85\] net504 vssd1 vssd1 vccd1 vccd1
+ _04949_ sky130_fd_sc_hd__o221a_1
X_05972_ top.WB.CPU_DAT_O\[29\] net1400 net345 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XANTENNA__05953__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08691_ top.cb_syn.end_check _04861_ _04893_ net1482 vssd1 vssd1 vccd1 vccd1 _01463_
+ sky130_fd_sc_hd__a31o_1
X_07711_ net258 _04293_ _04294_ net1175 net432 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a32o_1
X_07642_ top.cb_syn.h_element\[56\] top.cb_syn.h_element\[47\] _04176_ vssd1 vssd1
+ vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05705__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07573_ _04165_ _04172_ _04109_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__mux2_1
X_09312_ _05052_ _00053_ net256 vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__and3b_1
XANTENNA__08655__A1 _02538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06524_ net1456 _03338_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__xor2_1
X_09243_ _05207_ _05208_ top.cb_syn.zero_count\[0\] vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[0\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout231_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06455_ net1472 net298 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nand2_1
XANTENNA__09510__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05469__B2 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06386_ top.hist_data_o\[10\] top.hist_data_o\[9\] _03250_ vssd1 vssd1 vccd1 vccd1
+ _03251_ sky130_fd_sc_hd__and3_1
X_05406_ top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__inv_2
X_09174_ net1378 _02567_ top.WB.curr_state\[0\] _02615_ vssd1 vssd1 vccd1 vccd1 _00002_
+ sky130_fd_sc_hd__a22o_1
X_08125_ _04200_ _04611_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05337_ top.histogram.eof_n vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ top.cb_syn.zeroes\[1\] top.cb_syn.zeroes\[0\] vssd1 vssd1 vccd1 vccd1 _04567_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout698_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
X_07007_ net1671 net140 _03686_ net486 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a22o_1
XANTENNA__10391__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout865_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ top.WB.CPU_DAT_O\[10\] net1394 net320 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__mux2_1
XANTENNA__05944__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ net438 net1567 net252 top.findLeastValue.sum\[16\] _04453_ vssd1 vssd1 vccd1
+ vccd1 _01805_ sky130_fd_sc_hd__a221o_1
X_08889_ net1407 top.WB.CPU_DAT_O\[13\] net306 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__mux2_1
X_10920_ clknet_leaf_47_clk _01485_ _00310_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08894__A1 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10851_ clknet_leaf_2_clk _01445_ _00241_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_10782_ clknet_leaf_118_clk _01388_ _00172_ vssd1 vssd1 vccd1 vccd1 top.path\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05880__A1 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ clknet_leaf_87_clk _01968_ _00793_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08470__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ clknet_leaf_82_clk _01899_ _00724_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11265_ clknet_leaf_81_clk _01830_ _00655_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07909__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__and2_1
X_11196_ clknet_leaf_26_clk _01761_ _00586_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10147_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__and2_1
XANTENNA__05935__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ net786 net621 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05842__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A1 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06896__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_06240_ top.cb_syn.curr_index\[7\] _02584_ _03105_ net446 vssd1 vssd1 vccd1 vccd1
+ _03113_ sky130_fd_sc_hd__a22o_1
XANTENNA__05871__A1 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06171_ top.cb_syn.char_index\[4\] _03044_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold315 top.cb_syn.char_path\[109\] vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 top.cb_syn.char_path\[114\] vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 top.cb_syn.char_path\[45\] vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__and2_1
Xhold359 top.cb_syn.char_path\[48\] vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 top.hTree.node_reg\[37\] vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 top.path\[48\] vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout806 net808 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_2
X_09861_ net867 net702 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__and2_1
Xfanout839 net845 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout817 net826 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07376__B2 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07376__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout828 net835 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_1
X_09792_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ top.path\[34\] top.path\[35\] net510 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__mux2_1
X_05955_ top.compVal\[6\] net160 net143 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ _02223_ sky130_fd_sc_hd__a22o_1
X_08743_ net425 _04930_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout181_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08674_ top.cb_syn.i\[5\] top.cb_syn.i\[4\] _04881_ vssd1 vssd1 vccd1 vccd1 _04884_
+ sky130_fd_sc_hd__and3_1
X_05886_ net1623 top.WB.CPU_DAT_O\[12\] net351 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
XANTENNA__08876__A1 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06887__A0 top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07625_ net521 _04220_ _04222_ net516 vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07556_ _04154_ _04155_ net289 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06507_ top.histogram.total\[25\] _03339_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__and2_1
X_09226_ net1408 _05199_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07487_ top.dut.bit_buf\[2\] net40 net713 vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__mux2_1
X_06438_ net1108 _03290_ net300 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09157_ top.cb_syn.curr_state\[0\] _04206_ _04546_ _04544_ vssd1 vssd1 vccd1 vccd1
+ _00003_ sky130_fd_sc_hd__a31o_1
X_06369_ net1204 net165 _03235_ net208 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\] vssd1 vssd1 vccd1 vccd1
+ _04604_ sky130_fd_sc_hd__or2_1
X_09088_ net527 _05107_ _05111_ _05112_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08039_ net550 _02580_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11050_ clknet_leaf_24_clk _01615_ _00440_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09356__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ net855 net690 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__and2_1
XANTENNA__07634__S _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ net915 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ clknet_leaf_51_clk _01475_ _00293_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_11883_ net441 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06878__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10834_ clknet_leaf_116_clk _01428_ _00224_ vssd1 vssd1 vccd1 vccd1 top.path\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10765_ clknet_leaf_97_clk _01371_ _00155_ vssd1 vssd1 vccd1 vccd1 top.path\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10696_ clknet_leaf_21_clk _01327_ _00086_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11317_ clknet_leaf_44_clk _01882_ _00707_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11248_ clknet_leaf_76_clk net1432 _00638_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07358__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ clknet_leaf_38_clk _01744_ _00569_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07358__B2 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06318__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05740_ top.findLeastValue.alternator_timer\[1\] top.findLeastValue.alternator_timer\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__or2_1
X_05671_ net1411 net168 _02732_ net209 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08390_ top.cb_syn.char_path_n\[9\] net202 _04757_ vssd1 vssd1 vccd1 vccd1 _01628_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05541__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07410_ _02517_ net126 net124 _04035_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_35_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07341_ _03768_ _03770_ _03989_ top.findLeastValue.val1\[18\] top.findLeastValue.val2\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_18_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07818__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09995__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ _03730_ _03933_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06223_ top.sram_interface.init_counter\[7\] _03023_ vssd1 vssd1 vccd1 vccd1 _03096_
+ sky130_fd_sc_hd__xor2_1
X_09011_ net1685 _05081_ _05082_ top.TRN_char_index\[6\] vssd1 vssd1 vccd1 vccd1 _01332_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06154_ net454 _03028_ _03029_ _02608_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a211o_1
Xhold101 top.path\[37\] vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 top.cb_syn.char_path\[110\] vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold123 top.cb_syn.char_path\[94\] vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 top.cb_syn.left vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06085_ top.cb_syn.cb_length\[5\] top.cb_syn.i\[5\] vssd1 vssd1 vccd1 vccd1 _02985_
+ sky130_fd_sc_hd__and2b_1
Xhold167 top.histogram.sram_out\[28\] vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 top.hTree.node_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 top.path\[118\] vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 top.cb_syn.char_path\[50\] vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 net606 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_2
X_09913_ net858 net693 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__and2_1
Xhold189 top.histogram.sram_out\[18\] vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09338__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_2
Xfanout636 net637 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_2
Xfanout658 net660 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_2
Xfanout647 net651 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_2
Xfanout669 net670 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_2
X_09775_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__and2_1
X_06987_ _02505_ net125 _03660_ net1742 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06309__C1 top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05938_ top.compVal\[23\] net159 net145 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 _02240_ sky130_fd_sc_hd__a22o_1
X_08726_ net1678 _04916_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09889__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ top.cb_syn.end_cnt\[4\] _04871_ _04872_ _04868_ vssd1 vssd1 vccd1 vccd1 _01476_
+ sky130_fd_sc_hd__o22a_1
X_05869_ net1529 top.WB.CPU_DAT_O\[29\] net353 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_53_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout828_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ _04802_ _04804_ _04807_ top.cb_syn.end_cnt\[3\] _02540_ vssd1 vssd1 vccd1
+ vccd1 _04808_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07539_ top.cb_syn.char_path_n\[82\] top.cb_syn.char_path_n\[81\] top.cb_syn.char_path_n\[84\]
+ top.cb_syn.char_path_n\[83\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ net832 net667 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__and2_1
X_09209_ net1085 net291 _05188_ top.header_synthesis.write_num_lefts _03375_ vssd1
+ vssd1 vccd1 vccd1 top.header_synthesis.next_write_num_lefts sky130_fd_sc_hd__a32o_1
X_10481_ net840 net675 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_62_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10563__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05599__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold690 top.cb_syn.count\[6\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
X_11102_ clknet_leaf_56_clk _01667_ _00492_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09329__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ clknet_leaf_55_clk _01598_ _00423_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08632__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__A1 top.findLeastValue.sum\[45\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05771__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ net898 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_82_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ clknet_leaf_112_clk _02399_ _01238_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_11797_ clknet_leaf_119_clk net441 _01169_ vssd1 vssd1 vccd1 vccd1 top.WB.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_4
X_10817_ clknet_leaf_98_clk _01411_ _00207_ vssd1 vssd1 vccd1 vccd1 top.path\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08923__S _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ clknet_leaf_13_clk _00038_ _00138_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[0\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__09017__B2 top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ clknet_leaf_11_clk _01310_ _00069_ vssd1 vssd1 vccd1 vccd1 top.path\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08776__B1 _04917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06910_ _03394_ net134 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nand2_1
X_07890_ top.hTree.tree_reg\[19\] top.findLeastValue.sum\[19\] net286 vssd1 vssd1
+ vccd1 vccd1 _04438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06841_ top.compVal\[33\] top.findLeastValue.val1\[33\] net151 vssd1 vssd1 vccd1
+ vccd1 _03626_ sky130_fd_sc_hd__mux2_1
X_09560_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__and2_1
X_06772_ _02427_ top.findLeastValue.val2\[25\] vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__nand2_1
X_08511_ net1310 top.cb_syn.char_path_n\[48\] net243 vssd1 vssd1 vccd1 vccd1 _01531_
+ sky130_fd_sc_hd__mux2_1
X_09491_ net765 net600 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__and2_1
X_05723_ top.histogram.sram_out\[1\] net357 net408 top.hTree.node_reg\[1\] vssd1 vssd1
+ vccd1 vccd1 _02776_ sky130_fd_sc_hd__a22o_1
X_08442_ net1272 top.cb_syn.char_path_n\[117\] net235 vssd1 vssd1 vccd1 vccd1 _01600_
+ sky130_fd_sc_hd__mux2_1
X_05654_ top.cb_syn.char_path\[76\] net540 net529 top.cb_syn.char_path\[44\] vssd1
+ vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
X_08373_ top.cb_syn.char_path_n\[18\] net378 net335 top.cb_syn.char_path_n\[16\] net181
+ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a221o_1
X_05585_ net1019 net354 _02659_ _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_102_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07324_ _03860_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07255_ _03910_ _03924_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout311_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06206_ _02507_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07186_ _03772_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08231__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06137_ net1587 net164 net157 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21o_1
X_06068_ _02967_ _02963_ _02965_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout680_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_2
Xfanout411 _02611_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
Xfanout422 _02560_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
Xfanout433 net434 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_2
XANTENNA__05493__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 top.controller.state_reg\[1\] vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
Xfanout444 net72 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 net457 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
X_09827_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__and2_1
Xfanout499 top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_4
Xfanout488 top.cb_syn.wait_cycle vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
Xfanout477 net480 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_2
X_09758_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__and2_1
XANTENNA__07742__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ top.header_synthesis.enable top.header_synthesis.char_added top.header_synthesis.write_num_lefts
+ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__and2_1
X_11720_ clknet_leaf_72_clk _02270_ _01110_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10558__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ clknet_leaf_115_clk _02201_ _01041_ vssd1 vssd1 vccd1 vccd1 top.path\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_10602_ net743 net578 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ clknet_leaf_5_clk _02147_ _00972_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10533_ net817 net652 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10293__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ net828 net663 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10395_ net801 net636 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07981__A1 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05992__A0 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ clknet_leaf_47_clk _01581_ _00406_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05744__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06011__B top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ net949 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XANTENNA__06438__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11849_ clknet_leaf_114_clk _02382_ _01221_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_05370_ top.findLeastValue.val1\[35\] vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__inv_2
XANTENNA__07249__B1 top.findLeastValue.sum\[44\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08997__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07040_ top.findLeastValue.val1\[18\] top.findLeastValue.val1\[17\] top.findLeastValue.val1\[16\]
+ top.findLeastValue.val1\[15\] vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09992__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08991_ top.WB.CPU_DAT_O\[29\] net1268 net366 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__mux2_1
XANTENNA__06901__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ net476 _04478_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__or2_1
XANTENNA__05983__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ net417 _04423_ _04424_ net258 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__o211a_1
XANTENNA__07724__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06824_ top.findLeastValue.val2\[42\] net129 net119 _03617_ vssd1 vssd1 vccd1 vccd1
+ _02050_ sky130_fd_sc_hd__o22a_1
X_09612_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__and2_1
X_09543_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06755_ top.compVal\[12\] top.findLeastValue.val2\[12\] vssd1 vssd1 vccd1 vccd1 _03553_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout261_A _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__and2_1
X_05706_ top.histogram.sram_out\[4\] net357 net408 top.hTree.node_reg\[4\] _02761_
+ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a221o_1
X_06686_ _02406_ top.findLeastValue.val1\[45\] top.findLeastValue.val1\[46\] vssd1
+ vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a21o_1
XANTENNA__05760__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05637_ _02702_ _02703_ net468 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__o21a_1
X_08425_ top.cb_syn.h_element\[57\] top.cb_syn.h_element\[48\] net517 vssd1 vssd1
+ vccd1 vccd1 _04778_ sky130_fd_sc_hd__mux2_1
XANTENNA__07033__A top.findLeastValue.val1\[46\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ top.cb_syn.char_path_n\[26\] net194 _04740_ vssd1 vssd1 vccd1 vccd1 _01645_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05568_ net1460 net170 _02646_ net209 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07307_ _03746_ _03965_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ top.cb_syn.char_path_n\[61\] net371 net328 top.cb_syn.char_path_n\[59\] net174
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a221o_1
X_05499_ net461 _02583_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__and2_2
XFILLER_0_104_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09166__A_N top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07660__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ _03906_ _03908_ _03911_ _03913_ _03905_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o221a_1
X_07169_ top.findLeastValue.val2\[6\] top.findLeastValue.val1\[6\] vssd1 vssd1 vccd1
+ vccd1 _03845_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ net812 net647 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__and2_1
Xfanout230 net233 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xfanout241 net247 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05974__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 _04256_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
Xfanout274 net276 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
Xfanout296 _03376_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05726__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10569__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06151__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ clknet_leaf_80_clk _02253_ _01093_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08691__A2 _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ clknet_leaf_110_clk _02184_ _01024_ vssd1 vssd1 vccd1 vccd1 top.path\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08473__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11565_ clknet_leaf_7_clk _02130_ _00955_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
X_10516_ net755 net590 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__and2_1
X_11496_ clknet_leaf_119_clk _02061_ _00886_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ net815 net650 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__and2_1
X_11928__891 vssd1 vssd1 vccd1 vccd1 _11928__891/HI net891 sky130_fd_sc_hd__conb_1
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10378_ net759 net594 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__and2_1
XANTENNA__05965__B1 top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__B1 _02770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06540_ top.histogram.total\[12\] _03332_ net1503 vssd1 vssd1 vccd1 vccd1 _03355_
+ sky130_fd_sc_hd__a21oi_1
X_06471_ top.hist_data_o\[6\] _03248_ net298 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a21oi_1
X_05422_ top.cb_syn.left_check vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__inv_2
X_08210_ top.cb_syn.char_path_n\[99\] net200 _04667_ vssd1 vssd1 vccd1 vccd1 _01718_
+ sky130_fd_sc_hd__o21a_1
X_09190_ _02851_ _04255_ _05173_ net470 vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ top.cb_syn.cb_length\[0\] top.cb_syn.cb_length\[1\] vssd1 vssd1 vccd1 vccd1
+ _04631_ sky130_fd_sc_hd__nand2b_1
X_05353_ top.findLeastValue.val2\[18\] vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__inv_2
X_08072_ top.cb_syn.zeroes\[4\] _04569_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__or2_1
XANTENNA__06445__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06996__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07023_ top.findLeastValue.val2\[38\] top.findLeastValue.val2\[37\] top.findLeastValue.val2\[36\]
+ top.findLeastValue.val2\[35\] vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__and4_1
X_08974_ top.WB.CPU_DAT_O\[27\] top.cb_syn.h_element\[59\] net367 vssd1 vssd1 vccd1
+ vccd1 _01364_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 top.sram_interface.init_counter\[19\] vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 top.hTree.node_reg\[57\] vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 top.hTree.node_reg\[13\] vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ top.hTree.tree_reg\[12\] top.findLeastValue.sum\[12\] net285 vssd1 vssd1
+ vccd1 vccd1 _04466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold49 top.hTree.closing vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05708__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ top.hTree.tree_reg\[26\] top.findLeastValue.sum\[26\] net265 vssd1 vssd1
+ vccd1 vccd1 _04411_ sky130_fd_sc_hd__mux2_1
X_07787_ net479 _04354_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout643_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ _03526_ _03527_ _03604_ _02459_ top.compVal\[39\] vssd1 vssd1 vccd1 vccd1
+ _03605_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_65_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05490__B net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06738_ top.compVal\[0\] _02479_ _03533_ _03534_ _03535_ vssd1 vssd1 vccd1 vccd1
+ _03536_ sky130_fd_sc_hd__o311a_1
XANTENNA__06920__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ net747 net582 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__and2_1
X_09457_ net730 net565 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08408_ net1515 _02554_ _04766_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__mux2_1
XANTENNA__06133__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06669_ _02424_ top.findLeastValue.val1\[28\] top.findLeastValue.val1\[24\] _02428_
+ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ net1024 net221 _05271_ _05272_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08339_ top.cb_syn.char_path_n\[35\] net379 net332 top.cb_syn.char_path_n\[33\] net182
+ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ clknet_leaf_103_clk _01915_ _00740_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10301_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11281_ clknet_leaf_44_clk _01846_ _00671_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10571__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ net802 net637 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__and2_1
XANTENNA__05947__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_A gpio_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__and2_1
XANTENNA__08468__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06911__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ clknet_leaf_58_clk _01561_ _00386_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07547__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06124__B1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11617_ clknet_leaf_22_clk _02167_ _01007_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11548_ clknet_leaf_74_clk _02113_ _00938_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08931__S _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 top.path\[104\] vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 top.cb_syn.cb_length\[6\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ clknet_leaf_95_clk _02044_ _00869_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[36\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05938__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896__927 vssd1 vssd1 vccd1 vccd1 net927 _11896__927/LO sky130_fd_sc_hd__conb_1
X_07710_ net475 _04291_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05971_ top.WB.CPU_DAT_O\[30\] net1243 net346 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
X_08690_ top.cb_syn.cb_enable top.cb_syn.curr_state\[5\] net464 _04792_ vssd1 vssd1
+ vccd1 vccd1 _04893_ sky130_fd_sc_hd__and4_1
X_07641_ net1455 _04236_ _04212_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__mux2_1
X_07572_ _04168_ _04171_ _04110_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__mux2_1
XANTENNA__06902__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07538__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06523_ _03339_ net1545 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nor2_1
X_09311_ net754 net589 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ top.header_synthesis.write_zeroes _03388_ net491 vssd1 vssd1 vccd1 vccd1
+ _05208_ sky130_fd_sc_hd__a21oi_4
X_06454_ _03249_ _03252_ top.hist_data_o\[12\] vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09510__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09173_ net524 net424 _04585_ _05086_ _05171_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a221o_1
X_06385_ top.hist_data_o\[8\] _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05405_ top.findLeastValue.least1\[8\] vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05336_ top.cb_syn.count\[0\] vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__inv_2
X_08124_ top.cb_syn.cb_length\[3\] _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout224_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08055_ net514 _04548_ _04558_ _04565_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a211o_2
XANTENNA__05641__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07006_ net1779 net140 _03686_ net484 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a22o_1
XANTENNA__10391__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ top.WB.CPU_DAT_O\[11\] net1345 net320 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__mux2_1
X_07908_ net421 _04451_ _04452_ net263 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o211a_1
X_08888_ net1218 top.WB.CPU_DAT_O\[14\] net305 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__mux2_1
XANTENNA__08343__A1 top.cb_syn.char_path_n\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ net431 net1490 net248 top.findLeastValue.sum\[30\] _04397_ vssd1 vssd1 vccd1
+ vccd1 _01819_ sky130_fd_sc_hd__a221o_1
X_10850_ clknet_leaf_2_clk _01444_ _00240_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[2\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_27_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07529__S0 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__and2_1
X_10781_ clknet_leaf_118_clk _01387_ _00171_ vssd1 vssd1 vccd1 vccd1 top.path\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07854__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08036__B top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ clknet_leaf_89_clk _01967_ _00792_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ clknet_leaf_84_clk _01898_ _00723_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08052__A top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05632__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ clknet_leaf_68_clk _01829_ _00654_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07909__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ net820 net655 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__and2_1
X_11195_ clknet_leaf_28_clk _01760_ _00585_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10146_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__and2_1
X_10077_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__and2_1
XANTENNA__05699__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ clknet_leaf_38_clk _01544_ _00369_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06995__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06170_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold316 top.path\[91\] vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold305 top.path\[46\] vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold327 top.histogram.sram_out\[9\] vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 top.path\[94\] vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 top.path\[114\] vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__and2_1
Xfanout807 net808 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_1
XFILLER_0_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 net826 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_1
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_2
X_09791_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__and2_1
X_08811_ top.path\[36\] top.path\[37\] top.path\[38\] top.path\[39\] net512 net507
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__mux4_1
X_05954_ top.compVal\[7\] net160 net143 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ _02224_ sky130_fd_sc_hd__a22o_1
X_08742_ top.path\[120\] net403 net323 top.path\[121\] net429 vssd1 vssd1 vccd1 vccd1
+ _04931_ sky130_fd_sc_hd__o221a_1
X_08673_ top.cb_syn.i\[4\] _04881_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout174_A _04616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07624_ top.cb_syn.max_index\[5\] _04184_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__xnor2_1
X_05885_ net1562 top.WB.CPU_DAT_O\[13\] net351 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XANTENNA__06336__B1 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07555_ top.cb_syn.char_path_n\[18\] top.cb_syn.char_path_n\[17\] top.cb_syn.char_path_n\[20\]
+ top.cb_syn.char_path_n\[19\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06506_ top.histogram.total\[24\] top.histogram.total\[23\] _03338_ vssd1 vssd1 vccd1
+ vccd1 _03339_ sky130_fd_sc_hd__and3_1
X_07486_ _04045_ _04088_ _04089_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout439_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ top.header_synthesis.header\[1\] top.cb_syn.char_index\[1\] net490 vssd1
+ vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__mux2_1
X_06437_ top.hist_data_o\[19\] _03268_ _03272_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06368_ top.cb_syn.curr_index\[1\] _02584_ _03232_ _03234_ vssd1 vssd1 vccd1 vccd1
+ _03235_ sky130_fd_sc_hd__a211o_1
X_09156_ _05157_ _05159_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__or2_1
X_08107_ _04590_ _04593_ _04603_ _04589_ net1660 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a32o_1
X_06299_ _02600_ _03079_ _03168_ net361 net486 vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__a32o_1
X_09087_ top.sram_interface.CB_write_counter\[1\] top.sram_interface.CB_write_counter\[0\]
+ net460 top.sram_interface.word_cnt\[12\] vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_110_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_05319_ top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ _04549_ _04547_ _04545_ _02891_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__and4bb_1
XANTENNA__05496__A top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05614__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold850 top.findLeastValue.sum\[28\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08564__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ net855 net690 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__and2_1
X_09989_ net832 net667 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__and2_1
X_11951_ net914 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
X_10902_ clknet_leaf_50_clk _01474_ _00292_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11882_ net441 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ clknet_leaf_117_clk _01427_ _00223_ vssd1 vssd1 vccd1 vccd1 top.path\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05550__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ clknet_leaf_111_clk _01370_ _00154_ vssd1 vssd1 vccd1 vccd1 top.path\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09292__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ clknet_leaf_21_clk _01326_ _00085_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_101_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05605__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ clknet_leaf_44_clk _01881_ _00706_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11247_ clknet_leaf_77_clk _01812_ _00637_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11178_ clknet_leaf_38_clk _01743_ _00568_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[124\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_output68_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07825__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05670_ top.hTree.node_reg\[42\] net307 _02730_ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__06965__A _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07340_ _03770_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09995__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ top.histogram.eof_n _05080_ _05081_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__o21ba_2
X_07271_ top.findLeastValue.sum\[38\] net276 _03938_ _03939_ vssd1 vssd1 vccd1 vccd1
+ _01925_ sky130_fd_sc_hd__a22o_1
X_06222_ net482 net361 _02600_ _03094_ _03093_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a221o_1
XANTENNA__08243__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06153_ net458 net533 net407 _02592_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__a31o_1
Xhold102 net61 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 top.header_synthesis.header\[6\] vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 top.cb_syn.char_path\[69\] vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 net69 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ _02982_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nor2_1
Xhold146 top.cb_syn.char_path\[111\] vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 top.cb_syn.char_path\[127\] vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 top.histogram.sram_out\[19\] vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_2
Xhold179 _01533_ vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__and2_1
Xfanout615 net630 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__dlymetal6s2s_1
X_09843_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__and2_1
Xfanout626 net629 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09516__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 net651 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_2
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout389_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_1
X_09774_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__and2_1
X_06986_ _03667_ _03675_ _02504_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout556_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05937_ net1127 net158 net145 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 _02241_
+ sky130_fd_sc_hd__a22o_1
X_08725_ _04913_ top.sram_interface.TRN_counter\[0\] vssd1 vssd1 vccd1 vccd1 _04916_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_107_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _02540_ _04790_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or2_1
X_05868_ net1646 top.WB.CPU_DAT_O\[30\] net353 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ net522 _02890_ net423 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__a21o_1
X_08587_ _04805_ _04806_ net497 vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__mux2_1
X_07538_ top.cb_syn.char_path_n\[86\] top.cb_syn.char_path_n\[85\] top.cb_syn.char_path_n\[88\]
+ top.cb_syn.char_path_n\[87\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout723_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05799_ net455 _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07469_ net1023 net343 _04075_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ top.cb_syn.num_lefts\[7\] top.cb_syn.num_lefts\[6\] _04604_ _05187_ _02566_
+ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__o41a_1
X_10480_ net840 net675 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__and2_1
X_09139_ net543 net452 _02916_ _02921_ _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a41o_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11101_ clknet_leaf_56_clk _01666_ _00491_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[47\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold680 top.sram_interface.write_counter_FLV\[2\] vssd1 vssd1 vccd1 vccd1 net1631
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 top.cb_syn.zero_count\[5\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ clknet_leaf_55_clk _01597_ _00422_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09426__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08632__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05771__B2 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ net897 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_82_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ clknet_leaf_113_clk _02398_ _01237_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_10816_ clknet_leaf_97_clk _01410_ _00206_ vssd1 vssd1 vccd1 vccd1 top.path\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11796_ clknet_leaf_94_clk _02330_ _01168_ vssd1 vssd1 vccd1 vccd1 top.compVal\[45\]
+ sky130_fd_sc_hd__dfrtp_2
X_10747_ clknet_leaf_7_clk _00037_ _00137_ vssd1 vssd1 vccd1 vccd1 top.histogram.wr_r_en\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10678_ clknet_leaf_108_clk _01309_ _00068_ vssd1 vssd1 vccd1 vccd1 top.path\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06251__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ top.findLeastValue.val2\[34\] net128 net118 _03625_ vssd1 vssd1 vccd1 vccd1
+ _02042_ sky130_fd_sc_hd__o22a_1
X_06771_ _02425_ top.findLeastValue.val2\[27\] vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nand2_1
X_08510_ net1416 top.cb_syn.char_path_n\[49\] net243 vssd1 vssd1 vccd1 vccd1 _01532_
+ sky130_fd_sc_hd__mux2_1
X_05722_ _02773_ _02774_ net467 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__o21a_1
X_09490_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__and2_1
X_08441_ net1088 top.cb_syn.char_path_n\[118\] net235 vssd1 vssd1 vccd1 vccd1 _01601_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05653_ net1530 net168 _02717_ net210 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a22o_1
XANTENNA__09071__A _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05514__A1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ top.cb_syn.char_path_n\[18\] net199 _04748_ vssd1 vssd1 vccd1 vccd1 _01637_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05584_ top.histogram.sram_out\[24\] net359 net410 top.hTree.node_reg\[24\] vssd1
+ vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07323_ _03855_ _03858_ _03862_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07254_ net271 _03926_ _03927_ net277 net1727 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout137_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06205_ top.cw2\[3\] _03077_ top.cw2\[4\] vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05758__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ top.findLeastValue.val2\[16\] top.findLeastValue.val1\[16\] vssd1 vssd1 vccd1
+ vccd1 _03861_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout304_A _02918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06136_ net1031 net166 net157 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a21o_1
X_06067_ _02954_ _02957_ _02961_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__or4_1
Xfanout423 _02555_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_4
Xfanout412 _02580_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_2
Xfanout401 _02850_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08150__A _02538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 top.TRN_char_index\[2\] vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_2
Xfanout456 net457 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_2
Xfanout434 _02419_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_2
X_09826_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__and2_1
Xfanout489 top.cb_syn.wait_cycle vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_1
Xfanout467 net469 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_4
Xfanout478 net480 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_2
X_09757_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout840_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06969_ _03667_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__nor2_1
X_08708_ net1508 _04900_ _04901_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_68_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06950__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08639_ top.cb_syn.end_cnt\[4\] _04850_ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a21oi_1
X_11650_ clknet_leaf_115_clk _02200_ _01040_ vssd1 vssd1 vccd1 vccd1 top.path\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11581_ clknet_leaf_27_clk _02146_ _00971_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
X_10601_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ net817 net652 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__and2_1
X_10463_ net828 net663 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10394_ net801 net636 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__and2_1
XANTENNA__10590__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ clknet_leaf_47_clk _01580_ _00405_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06941__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11917_ net948 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11848_ clknet_leaf_112_clk _02381_ _01220_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07249__B2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ clknet_leaf_3_clk _00014_ _01151_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09410__A2 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ top.WB.CPU_DAT_O\[30\] net1206 net366 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__mux2_1
X_07941_ top.hTree.tree_reg\[9\] top.findLeastValue.sum\[9\] net266 vssd1 vssd1 vccd1
+ vccd1 _04479_ sky130_fd_sc_hd__mux2_1
X_07872_ net475 _04422_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05735__A1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06823_ top.compVal\[42\] top.findLeastValue.val1\[42\] net153 vssd1 vssd1 vccd1
+ vccd1 _03617_ sky130_fd_sc_hd__mux2_1
X_09611_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__and2_1
XANTENNA__06932__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09542_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__and2_1
X_06754_ top.compVal\[13\] _02473_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09005__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05705_ top.hTree.node_reg\[36\] net307 _02760_ net469 vssd1 vssd1 vccd1 vccd1 _02761_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ net837 net672 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_90_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
X_06685_ _02414_ top.findLeastValue.val1\[33\] vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nand2_1
X_05636_ top.cb_syn.char_path\[47\] net531 net312 top.cb_syn.char_path\[111\] vssd1
+ vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a22o_1
X_08424_ top.cb_syn.char_index\[3\] _04777_ _04772_ vssd1 vssd1 vccd1 vccd1 _01614_
+ sky130_fd_sc_hd__mux2_1
X_08355_ top.cb_syn.char_path_n\[27\] net373 net327 top.cb_syn.char_path_n\[25\] net176
+ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a221o_1
X_05567_ top.histogram.sram_out\[27\] net359 _02644_ _02645_ vssd1 vssd1 vccd1 vccd1
+ _02646_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_63_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _03746_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__or2_1
X_08286_ top.cb_syn.char_path_n\[61\] net193 _04705_ vssd1 vssd1 vccd1 vccd1 _01680_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06999__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05498_ net535 _02582_ top.sram_interface.word_cnt\[9\] vssd1 vssd1 vccd1 vccd1 _02583_
+ sky130_fd_sc_hd__a21o_1
X_07237_ _03897_ _03900_ _03899_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07168_ top.findLeastValue.val2\[7\] top.findLeastValue.val1\[7\] vssd1 vssd1 vccd1
+ vccd1 _03844_ sky130_fd_sc_hd__or2_1
X_06119_ _02997_ _02998_ _03012_ _02996_ net1673 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07099_ top.findLeastValue.val2\[19\] top.findLeastValue.val1\[19\] top.findLeastValue.val1\[18\]
+ top.findLeastValue.val2\[18\] vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o211a_1
Xfanout231 net233 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout220 net223 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
XANTENNA__08599__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_4
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_4
Xfanout253 _04337_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
X_09809_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__and2_1
Xfanout286 _04249_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_4
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
XANTENNA__06923__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10569__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
X_11702_ clknet_leaf_85_clk _02252_ _01092_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11633_ clknet_leaf_110_clk _02183_ _01023_ vssd1 vssd1 vccd1 vccd1 top.path\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ clknet_leaf_6_clk _02129_ _00954_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ net756 net591 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__and2_1
X_11495_ clknet_leaf_0_clk _02060_ _00885_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10446_ net815 net650 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10377_ net759 net594 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__and2_1
XANTENNA__09614__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06470_ net1527 net297 _03309_ _03310_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05421_ top.cb_syn.char_path_n\[0\] vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\] vssd1 vssd1 vccd1 vccd1
+ _04630_ sky130_fd_sc_hd__nand2b_1
X_05352_ top.findLeastValue.val2\[19\] vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__inv_2
X_08071_ _04573_ _04576_ _04579_ _04566_ top.cb_syn.zeroes\[5\] vssd1 vssd1 vccd1
+ vccd1 _01769_ sky130_fd_sc_hd__a32o_1
X_07022_ top.findLeastValue.val2\[46\] top.findLeastValue.val2\[45\] top.findLeastValue.val2\[44\]
+ top.findLeastValue.val2\[43\] vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__and4_1
X_08973_ top.WB.CPU_DAT_O\[28\] top.cb_syn.h_element\[60\] net368 vssd1 vssd1 vccd1
+ vccd1 _01365_ sky130_fd_sc_hd__mux2_1
XANTENNA__05956__B2 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold17 top.sram_interface.init_counter\[21\] vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 top.hTree.node_reg\[12\] vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ net438 top.hTree.tree_reg\[13\] net251 net1559 _04465_ vssd1 vssd1 vccd1
+ vccd1 _01802_ sky130_fd_sc_hd__a221o_1
XANTENNA__09147__A1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08355__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 top.hTree.node_reg\[58\] vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout371_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ top.hTree.tree_reg\[26\] top.findLeastValue.sum\[26\] net281 vssd1 vssd1
+ vccd1 vccd1 _04410_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout469_A top.controller.state_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07786_ top.hTree.tree_reg\[40\] top.findLeastValue.sum\[40\] net267 vssd1 vssd1
+ vccd1 vccd1 _04355_ sky130_fd_sc_hd__mux2_1
X_06806_ _03599_ _03600_ _03601_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_65_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ net745 net580 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__and2_1
X_06737_ top.compVal\[1\] top.findLeastValue.val2\[1\] vssd1 vssd1 vccd1 vccd1 _03535_
+ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_63_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
X_09456_ net730 net565 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06668_ _02427_ top.findLeastValue.val1\[25\] vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__and2_1
X_08407_ net522 net523 _04559_ _04561_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__o211a_1
X_05619_ _02687_ _02688_ net467 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__o21a_1
XANTENNA__07330__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ top.hTree.nulls\[55\] net398 net228 vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout803_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06599_ top.compVal\[15\] top.compVal\[14\] top.compVal\[13\] top.compVal\[12\] vssd1
+ vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__or4_1
X_08338_ top.cb_syn.char_path_n\[35\] net200 _04731_ vssd1 vssd1 vccd1 vccd1 _01654_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08269_ top.cb_syn.char_path_n\[70\] net375 net333 top.cb_syn.char_path_n\[68\] net178
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05644__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11280_ clknet_leaf_45_clk _01845_ _00670_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_10300_ net855 net690 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10231_ net803 net638 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__and2_1
XANTENNA__07397__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__and2_1
X_10093_ net833 net668 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__and2_1
XANTENNA__05947__B2 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07653__S _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__B1 _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10995_ clknet_leaf_59_clk _01560_ _00385_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[77\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_54_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07547__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ clknet_leaf_24_clk _02166_ _01006_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11547_ clknet_leaf_74_clk _02112_ _00937_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05635__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold509 net92 vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
X_11478_ clknet_leaf_95_clk _02043_ _00868_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[35\]
+ sky130_fd_sc_hd__dfstp_1
X_10429_ net818 net653 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__and2_1
XANTENNA__09129__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05938__B2 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05970_ top.WB.CPU_DAT_O\[31\] net1399 net346 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08352__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ top.cb_syn.max_index\[3\] _04181_ _04232_ _04235_ vssd1 vssd1 vccd1 vccd1
+ _04236_ sky130_fd_sc_hd__o22a_1
XANTENNA__09998__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ _04169_ _04170_ net289 vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
XANTENNA__07538__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ top.header_synthesis.write_zeroes _05194_ _03388_ vssd1 vssd1 vccd1 vccd1
+ top.header_synthesis.next_write_zeroes sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_45_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
X_06522_ top.histogram.total\[23\] _03338_ net1544 vssd1 vssd1 vccd1 vccd1 _03348_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06907__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09241_ top.header_synthesis.write_zeroes _03388_ _05194_ vssd1 vssd1 vccd1 vccd1
+ _05207_ sky130_fd_sc_hd__and3_2
X_06453_ net298 _03255_ _03298_ _03299_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__o31ai_1
XANTENNA__07863__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ _02896_ _05169_ _05170_ net464 vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__o31a_1
X_05404_ top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06384_ top.hist_data_o\[7\] top.hist_data_o\[6\] _03248_ vssd1 vssd1 vccd1 vccd1
+ _03249_ sky130_fd_sc_hd__and3_2
XFILLER_0_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05335_ top.cb_syn.count\[1\] vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__inv_2
X_08123_ top.cb_syn.cb_length\[2\] top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\]
+ _04611_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11944__907 vssd1 vssd1 vccd1 vccd1 _11944__907/HI net907 sky130_fd_sc_hd__conb_1
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ net515 _04563_ _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07005_ net1664 net140 _03686_ net483 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout586_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920__951 vssd1 vssd1 vccd1 vccd1 net951 _11920__951/LO sky130_fd_sc_hd__conb_1
X_08956_ top.WB.CPU_DAT_O\[12\] net1217 net320 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__mux2_1
XANTENNA__05782__A top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07907_ net478 _04450_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__or2_1
X_08887_ net1200 top.WB.CPU_DAT_O\[15\] net305 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout753_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ net417 _04395_ _04396_ net255 vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__o211a_1
XANTENNA__06354__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07529__S1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
X_07769_ net437 net1450 net252 top.findLeastValue.sum\[44\] _04341_ vssd1 vssd1 vccd1
+ vccd1 _01833_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09508_ net733 net568 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ clknet_leaf_118_clk _01386_ _00170_ vssd1 vssd1 vccd1 vccd1 top.path\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06817__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07854__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05865__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ clknet_leaf_91_clk _01966_ _00791_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05617__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__S _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold798_A top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ clknet_leaf_84_clk _01897_ _00722_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ clknet_leaf_81_clk _01828_ _00653_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_11194_ clknet_leaf_27_clk _01759_ _00584_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_10214_ net820 net655 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__and2_1
X_10145_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10076_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__and2_1
XANTENNA__07542__A0 _04134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06896__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10978_ clknet_leaf_38_clk _01543_ _00368_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09047__A0 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05608__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold317 top.hTree.nulls\[61\] vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold306 top.path\[70\] vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 net99 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09058__B _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06820__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold328 top.path\[122\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout808 net816 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout819 net826 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_2
X_08810_ top.path\[40\] net405 _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__o21a_1
X_11904__935 vssd1 vssd1 vccd1 vccd1 net935 _11904__935/LO sky130_fd_sc_hd__conb_1
X_09790_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__and2_1
X_05953_ top.compVal\[8\] net161 net144 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ _02225_ sky130_fd_sc_hd__a22o_1
X_08741_ top.path\[122\] top.path\[123\] net512 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__mux2_1
X_08672_ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05884_ net1606 top.WB.CPU_DAT_O\[14\] net351 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
X_07623_ net517 top.cb_syn.h_element\[50\] net525 top.cb_syn.h_element\[59\] _04180_
+ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout167_A _02621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ top.cb_syn.char_path_n\[22\] top.cb_syn.char_path_n\[21\] top.cb_syn.char_path_n\[24\]
+ top.cb_syn.char_path_n\[23\] net394 net292 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06505_ top.histogram.total\[22\] top.histogram.total\[21\] _03336_ vssd1 vssd1 vccd1
+ vccd1 _03338_ sky130_fd_sc_hd__and3_1
X_07485_ top.dut.out\[3\] net344 _04056_ _04060_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ net296 _05198_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[0\]
+ sky130_fd_sc_hd__and2_1
X_06436_ net1167 _03289_ net300 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XANTENNA__09038__A0 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06367_ _02588_ _03013_ _03233_ net446 _03228_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a221o_1
X_09155_ net447 top.sram_interface.word_cnt\[14\] _05158_ net535 _02607_ vssd1 vssd1
+ vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
X_08106_ top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\] top.cb_syn.num_lefts\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a21o_1
X_06298_ top.cw2\[4\] top.cw2\[3\] _03077_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__or3_1
X_09086_ top.sram_interface.word_cnt\[6\] _02795_ _02839_ net537 _05076_ vssd1 vssd1
+ vccd1 vccd1 _05111_ sky130_fd_sc_hd__a221o_1
XANTENNA__05777__A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05318_ top.compVal\[11\] vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__inv_2
X_08037_ net514 _04548_ net423 vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a21o_1
XANTENNA__05496__B top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold840 top.findLeastValue.sum\[41\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 top.compVal\[45\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__and2_1
X_08939_ top.WB.CPU_DAT_O\[29\] net1414 net319 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__mux2_1
X_11950_ net913 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_10901_ clknet_leaf_51_clk _01473_ _00291_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07931__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ net883 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XANTENNA__06878__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05550__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ clknet_leaf_117_clk _01426_ _00222_ vssd1 vssd1 vccd1 vccd1 top.path\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10763_ clknet_leaf_111_clk _01369_ _00153_ vssd1 vssd1 vccd1 vccd1 top.path\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09029__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10694_ clknet_leaf_107_clk _01325_ _00084_ vssd1 vssd1 vccd1 vccd1 top.path\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11315_ clknet_leaf_43_clk _01880_ _00705_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11246_ clknet_leaf_73_clk _01811_ _00636_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11177_ clknet_leaf_35_clk _01742_ _00567_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10128_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10059_ net719 net554 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__and2_1
XANTENNA__06318__A1 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__B net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07818__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07270_ _03724_ _03934_ net270 vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06221_ _02505_ _03081_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__xnor2_1
X_06152_ top.sram_interface.init_counter\[10\] _03025_ _03026_ vssd1 vssd1 vccd1 vccd1
+ _03028_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08779__C1 top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06083_ top.cb_syn.cb_length\[1\] top.cb_syn.i\[1\] vssd1 vssd1 vccd1 vccd1 _02983_
+ sky130_fd_sc_hd__and2b_1
Xhold114 top.path\[81\] vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 top.path\[3\] vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 top.path\[39\] vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _01594_ vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 top.cb_syn.char_path\[56\] vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold158 top.hTree.node_reg\[2\] vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_2
Xhold169 top.cb_syn.char_path\[68\] vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
X_09842_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__and2_1
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_2
Xfanout616 net630 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09516__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout649 net651 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_2
Xfanout638 net643 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_2
X_09773_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__and2_1
X_06985_ _02574_ _03087_ _03675_ _03667_ net487 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout284_A _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _04915_ top.sram_interface.TRN_counter\[2\] _04913_ vssd1 vssd1 vccd1 vccd1
+ _01452_ sky130_fd_sc_hd__mux2_1
X_05936_ top.compVal\[25\] net158 net146 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 _02242_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _02538_ _04790_ _04866_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a21oi_1
X_05867_ net1526 top.WB.CPU_DAT_O\[31\] net353 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout451_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout549_A top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ net488 net423 vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__or2_1
X_08586_ top.cb_syn.char_path_n\[67\] top.cb_syn.char_path_n\[68\] top.cb_syn.char_path_n\[71\]
+ top.cb_syn.char_path_n\[72\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__mux4_1
X_07537_ _04135_ _04136_ net289 vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05798_ net542 net533 net527 _02821_ _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__o311a_1
XANTENNA__07809__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _04060_ _04070_ _04074_ _04045_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__a22o_1
X_09207_ top.cb_syn.num_lefts\[5\] top.cb_syn.num_lefts\[4\] top.cb_syn.num_lefts\[3\]
+ top.cb_syn.num_lefts\[2\] vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__or4_1
X_06419_ net1653 _03279_ net301 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
X_07399_ _03829_ net271 _04029_ net277 net1724 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a32o_1
X_09138_ _02858_ _02880_ _05143_ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_118_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05300__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05599__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ clknet_leaf_62_clk _01665_ _00490_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07926__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ net460 net526 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nand2_1
Xhold670 top.cb_syn.cb_enable vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 top.histogram.total\[10\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ clknet_leaf_55_clk _01596_ _00421_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[113\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold692 top.histogram.total\[21\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09426__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05771__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ net896 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ clknet_leaf_113_clk _02397_ _01236_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_10815_ clknet_leaf_111_clk _01409_ _00205_ vssd1 vssd1 vccd1 vccd1 top.path\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11795_ clknet_leaf_92_clk _02329_ _01167_ vssd1 vssd1 vccd1 vccd1 top.compVal\[44\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_15_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07897__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ clknet_leaf_6_clk _00036_ _00136_ vssd1 vssd1 vccd1 vccd1 top.histogram.wr_r_en\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ clknet_leaf_108_clk _01308_ _00067_ vssd1 vssd1 vccd1 vccd1 top.path\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07836__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ clknet_leaf_83_clk _01794_ _00619_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06041__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _02425_ top.findLeastValue.val2\[27\] top.findLeastValue.val2\[26\] _02426_
+ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__o22a_1
X_05721_ top.cb_syn.char_path\[33\] net530 net311 top.cb_syn.char_path\[97\] vssd1
+ vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__a22o_1
X_08440_ net1099 top.cb_syn.char_path_n\[119\] net235 vssd1 vssd1 vccd1 vccd1 _01602_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05652_ top.histogram.sram_out\[13\] net358 net409 top.hTree.node_reg\[13\] _02716_
+ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08371_ top.cb_syn.char_path_n\[19\] net378 net334 top.cb_syn.char_path_n\[17\] net181
+ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05583_ _02657_ _02658_ net465 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_102_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07322_ net268 _03955_ _03976_ net274 net1627 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a32o_1
X_07253_ _03907_ _03925_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__nand2_1
XANTENNA__08216__A1 top.cb_syn.char_path_n\[96\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06204_ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__inv_2
X_07184_ _03768_ _03769_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06135_ net1042 net166 net157 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_57_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06066_ top.cb_syn.zeroes\[0\] _02556_ _02956_ _02962_ vssd1 vssd1 vccd1 vccd1 _02966_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09527__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _02810_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_2
X_09825_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__and2_1
Xfanout424 _02555_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_2
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 _02419_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
Xfanout457 top.controller.state_reg\[2\] vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout666_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__and2_1
X_06968_ net485 net486 _03088_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nand3_1
X_09687_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__and2_1
X_08707_ _04904_ _04901_ net1739 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__mux2_1
X_05919_ net442 _02898_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__or2_1
X_08638_ top.cb_syn.end_cnt\[3\] _04857_ _04854_ _02540_ vssd1 vssd1 vccd1 vccd1 _04858_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_68_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ top.compVal\[4\] top.findLeastValue.val1\[4\] net153 vssd1 vssd1 vccd1 vccd1
+ _03655_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net496 net498 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__nor2_1
XANTENNA__06825__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ net799 net634 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ clknet_leaf_5_clk _02145_ _00970_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
X_10531_ net805 net640 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__and2_1
X_10462_ net828 net663 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10393_ net748 net583 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__and2_1
XANTENNA__07966__A0 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ clknet_leaf_46_clk _01579_ _00404_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07718__B1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11916_ net947 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_11847_ clknet_leaf_114_clk _02380_ _01219_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ clknet_leaf_3_clk _00013_ _01150_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ clknet_leaf_17_clk _01360_ _00119_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ top.hTree.tree_reg\[9\] top.findLeastValue.sum\[9\] net285 vssd1 vssd1 vccd1
+ vccd1 _04478_ sky130_fd_sc_hd__mux2_1
X_07871_ top.hTree.tree_reg\[23\] top.findLeastValue.sum\[23\] net264 vssd1 vssd1
+ vccd1 vccd1 _04423_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ top.findLeastValue.val2\[43\] net129 net119 _03616_ vssd1 vssd1 vccd1 vccd1
+ _02051_ sky130_fd_sc_hd__o22a_1
X_09610_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__and2_1
X_06753_ top.compVal\[13\] _02473_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__and2_1
XANTENNA__08134__B1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05704_ _02758_ _02759_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ net837 net672 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__and2_1
XANTENNA__10021__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06684_ top.compVal\[38\] _02485_ _02486_ top.compVal\[37\] _03481_ vssd1 vssd1 vccd1
+ vccd1 _03482_ sky130_fd_sc_hd__a221o_1
X_05635_ top.cb_syn.char_path\[15\] net549 net540 top.cb_syn.char_path\[79\] vssd1
+ vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a22o_1
X_08423_ top.cb_syn.h_element\[58\] top.cb_syn.h_element\[49\] net517 vssd1 vssd1
+ vccd1 vccd1 _04777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07893__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ top.cb_syn.char_path_n\[27\] net194 _04739_ vssd1 vssd1 vccd1 vccd1 _01646_
+ sky130_fd_sc_hd__o21a_1
X_05566_ top.hTree.node_reg\[59\] net354 net410 top.hTree.node_reg\[27\] vssd1 vssd1
+ vccd1 vccd1 _02645_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07305_ _03747_ _03958_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nand2_1
X_08285_ top.cb_syn.char_path_n\[62\] net371 net328 top.cb_syn.char_path_n\[60\] net175
+ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a221o_1
X_05497_ _02581_ top.cb_syn.setup net514 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__or3b_2
XFILLER_0_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07660__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07236_ _03902_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ top.findLeastValue.val2\[7\] top.findLeastValue.val1\[7\] vssd1 vssd1 vccd1
+ vccd1 _03843_ sky130_fd_sc_hd__and2_1
X_06118_ top.cb_syn.count\[1\] top.cb_syn.count\[0\] vssd1 vssd1 vccd1 vccd1 _03012_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07098_ _03768_ _03769_ _03770_ _03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__and4_1
X_06049_ _02947_ _02948_ _02945_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a21o_1
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
Xfanout221 net223 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
Xfanout210 net212 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
XANTENNA__08599__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 net246 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
Xfanout265 _04251_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
XANTENNA__08373__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__and2_1
Xfanout287 _03394_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_2
Xfanout298 net299 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
X_09739_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__and2_1
XANTENNA__05726__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09720__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ clknet_leaf_19_clk net957 _01091_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.CB_read_counter
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11632_ clknet_leaf_10_clk _02182_ _01022_ vssd1 vssd1 vccd1 vccd1 top.TRN_sram_complete
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ clknet_leaf_6_clk _02128_ _00953_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
X_10514_ net756 net591 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__and2_1
X_11494_ clknet_leaf_2_clk _02059_ _00884_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10445_ net806 net641 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ net761 net596 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__and2_1
XANTENNA__09614__B net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08667__B2 _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05420_ top.cb_syn.char_index\[1\] vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__inv_2
X_05351_ top.findLeastValue.val2\[24\] vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__inv_2
X_08070_ _02528_ _04571_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07021_ top.findLeastValue.val2\[42\] top.findLeastValue.val2\[41\] top.findLeastValue.val2\[40\]
+ top.findLeastValue.val2\[39\] vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__and4_1
XANTENNA__06850__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ top.WB.CPU_DAT_O\[29\] top.cb_syn.h_element\[61\] net367 vssd1 vssd1 vccd1
+ vccd1 _01366_ sky130_fd_sc_hd__mux2_1
XANTENNA__10016__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 top.hTree.node_reg\[45\] vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ net420 _04463_ _04464_ net262 vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__o211a_1
Xhold29 top.hTree.finish_check vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout197_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ net434 net1558 net248 top.findLeastValue.sum\[27\] _04409_ vssd1 vssd1 vccd1
+ vccd1 _01816_ sky130_fd_sc_hd__a221o_1
XANTENNA__05708__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ _02415_ top.findLeastValue.val2\[32\] _03517_ _03518_ _03602_ vssd1 vssd1
+ vccd1 vccd1 _03603_ sky130_fd_sc_hd__o2111a_1
X_07785_ top.hTree.tree_reg\[40\] top.findLeastValue.sum\[40\] net285 vssd1 vssd1
+ vccd1 vccd1 _04354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ net797 net632 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__and2_1
X_06736_ top.compVal\[2\] top.findLeastValue.val2\[2\] vssd1 vssd1 vccd1 vccd1 _03534_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__and2_1
XANTENNA__09540__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ _02421_ top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__or2_1
X_05618_ top.cb_syn.char_path\[50\] net530 net311 top.cb_syn.char_path\[114\] vssd1
+ vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a22o_1
XANTENNA__06133__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ top.cb_syn.char_path_n\[1\] net192 _04765_ vssd1 vssd1 vccd1 vccd1 _01620_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07330__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09386_ net399 _04292_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__nand2_1
X_06598_ top.compVal\[11\] top.compVal\[10\] top.compVal\[9\] top.compVal\[8\] vssd1
+ vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__or4_1
XANTENNA__05892__A1 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ top.cb_syn.char_path_n\[36\] net379 net336 top.cb_syn.char_path_n\[34\] net182
+ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a221o_1
X_05549_ top.hTree.node_reg\[62\] net356 _02629_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ net1763 net196 _04696_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__o21a_1
XANTENNA__08830__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07219_ _03733_ _03890_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__o21ai_4
X_08199_ top.cb_syn.char_path_n\[105\] net380 net337 top.cb_syn.char_path_n\[103\]
+ net183 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10230_ net802 net637 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__and2_1
XANTENNA__08594__A0 top.cb_syn.char_path_n\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06123__B net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__and2_1
XANTENNA__05947__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10092_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__and2_1
XANTENNA__08897__A1 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ clknet_leaf_60_clk net1540 _00384_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08649__A1 _02538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05580__B1 _02656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ clknet_leaf_22_clk _02165_ _01005_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05883__A1 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ clknet_leaf_73_clk _02111_ _00936_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06832__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ clknet_leaf_96_clk _02042_ _00867_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08585__A0 top.cb_syn.char_path_n\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09377__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ net818 net653 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__and2_1
X_10359_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__and2_1
XANTENNA__05938__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__A1 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ top.cb_syn.char_path_n\[50\] top.cb_syn.char_path_n\[49\] top.cb_syn.char_path_n\[52\]
+ top.cb_syn.char_path_n\[51\] net396 net292 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__mux4_1
X_06521_ _03340_ _03347_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09240_ net1232 _05206_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[8\]
+ sky130_fd_sc_hd__mux2_1
X_06452_ net1312 net298 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__nand2_1
X_09171_ _02581_ _02887_ _04605_ _02551_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a22o_1
XANTENNA__05874__A1 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05403_ top.findLeastValue.least2\[1\] vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06383_ _03246_ _03247_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__and2_1
XANTENNA__09065__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05334_ top.cb_syn.count\[2\] vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__inv_2
X_08122_ _04560_ _04605_ _04614_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__or3_2
XFILLER_0_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ net515 net522 net523 net514 _04561_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__o41a_1
XFILLER_0_114_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ net1644 net140 _03686_ net482 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout112_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08955_ top.WB.CPU_DAT_O\[13\] net1253 net320 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__mux2_1
X_07906_ top.hTree.tree_reg\[16\] top.findLeastValue.sum\[16\] net267 vssd1 vssd1
+ vccd1 vccd1 _04451_ sky130_fd_sc_hd__mux2_1
XANTENNA__05782__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08886_ net1162 top.WB.CPU_DAT_O\[16\] net302 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__mux2_1
XANTENNA__08879__A1 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07000__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ net470 _04394_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__or2_1
X_07768_ net421 _04339_ _04340_ net262 vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout746_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09507_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__and2_1
X_06719_ _02409_ top.findLeastValue.val2\[38\] vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07699_ net257 _04283_ _04284_ net1073 net432 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_55_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09438_ net733 net568 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ net398 _04317_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__nand2_1
XANTENNA__05865__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05865__B2 top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ clknet_leaf_90_clk _01965_ _00790_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06833__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ clknet_leaf_84_clk _01896_ _00721_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09359__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11262_ clknet_leaf_81_clk _01827_ _00652_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_11193_ clknet_leaf_27_clk _01758_ _00583_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10213_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__and2_1
X_10144_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__and2_1
XANTENNA_input42_A gpio_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07790__A1 top.findLeastValue.sum\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10075_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__and2_1
XANTENNA__05553__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ clknet_leaf_37_clk _01542_ _00367_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11529_ clknet_leaf_81_clk _02094_ _00919_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold307 top.path\[66\] vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 top.cb_syn.char_path\[85\] vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold329 top.cb_syn.char_path\[122\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11885__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net812 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07781__A1 top.findLeastValue.sum\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05952_ top.compVal\[9\] net161 net144 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ _02226_ sky130_fd_sc_hd__a22o_1
X_08740_ top.path\[124\] net405 _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__o21a_1
X_08671_ top.cb_syn.i\[3\] top.cb_syn.i\[2\] top.cb_syn.i\[1\] top.cb_syn.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05883_ net1790 top.WB.CPU_DAT_O\[15\] net351 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07622_ top.cb_syn.h_element\[59\] top.cb_syn.h_element\[50\] _04176_ vssd1 vssd1
+ vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
X_07553_ _04151_ _04152_ net289 vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06219__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06504_ top.histogram.total\[21\] _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__and2_1
X_07484_ _04077_ _04087_ net342 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ top.header_synthesis.header\[0\] top.cb_syn.char_index\[0\] net490 vssd1
+ vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__mux2_1
X_06435_ top.hist_data_o\[20\] _03272_ _03258_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout327_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ net440 net451 net456 net406 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08105_ _04590_ _04594_ _04602_ _04589_ top.cb_syn.num_lefts\[3\] vssd1 vssd1 vccd1
+ vccd1 _01758_ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06366_ top.cb_syn.max_index\[1\] _03102_ _03104_ top.hTree.nullSumIndex\[0\] vssd1
+ vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06297_ _02602_ _03166_ _03165_ net534 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__o211a_1
X_09085_ net459 net534 _02576_ _05110_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__a31o_1
XANTENNA__05777__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05317_ top.compVal\[15\] vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__inv_2
Xhold830 top.cb_syn.char_path_n\[25\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08036_ top.cb_syn.end_cond top.CB_write_complete vssd1 vssd1 vccd1 vccd1 _04548_
+ sky130_fd_sc_hd__nand2b_1
Xhold841 top.cb_syn.char_path_n\[75\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold852 top.histogram.total\[14\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__and2_1
X_08938_ top.WB.CPU_DAT_O\[30\] net1289 net319 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _05035_ _05048_ _05049_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__and3_1
X_10900_ clknet_leaf_51_clk _01472_ _00290_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_11880_ net882 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__05535__B1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10831_ clknet_leaf_116_clk _01425_ _00221_ vssd1 vssd1 vccd1 vccd1 top.path\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10762_ clknet_leaf_12_clk _00043_ _00152_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ clknet_leaf_107_clk _01324_ _00083_ vssd1 vssd1 vccd1 vccd1 top.path\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05968__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11314_ clknet_leaf_41_clk _01879_ _00704_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11245_ clknet_leaf_73_clk net1553 _00635_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08635__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11176_ clknet_leaf_37_clk _01741_ _00566_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08960__A0 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__and2_1
XANTENNA__05774__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ net719 net554 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06318__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06220_ _02602_ _03086_ _03092_ _02603_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06151_ net1048 net164 net157 _03027_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a211o_1
X_06082_ top.cb_syn.i\[1\] top.cb_syn.cb_length\[1\] vssd1 vssd1 vccd1 vccd1 _02982_
+ sky130_fd_sc_hd__and2b_1
Xhold115 top.hTree.tree_reg\[53\] vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 net67 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 top.path\[23\] vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 top.cb_syn.char_path\[118\] vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 top.cb_syn.char_path\[119\] vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ net839 net674 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__and2_1
Xhold159 top.path\[5\] vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout606 net612 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09841_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__and2_1
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_2
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_2
Xfanout639 net643 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08951__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__and2_1
XANTENNA__07754__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06984_ top.findLeastValue.histo_index\[2\] _03667_ _03675_ _03205_ vssd1 vssd1 vccd1
+ vccd1 _01951_ sky130_fd_sc_hd__a22o_1
XANTENNA__05765__B1 _02806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05935_ top.compVal\[26\] net158 net146 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 _02243_ sky130_fd_sc_hd__a22o_1
X_08723_ _02913_ _04914_ _02589_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout277_A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _04867_ _04870_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05866_ net439 net453 top.histogram.state\[2\] vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__and3_1
X_07605_ _02525_ top.cb_syn.curr_state\[0\] _04178_ net488 _04204_ vssd1 vssd1 vccd1
+ vccd1 _04205_ sky130_fd_sc_hd__a221o_1
X_08585_ top.cb_syn.char_path_n\[65\] top.cb_syn.char_path_n\[66\] top.cb_syn.char_path_n\[69\]
+ top.cb_syn.char_path_n\[70\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__mux4_1
X_05797_ net444 net527 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout444_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ top.cb_syn.char_path_n\[90\] top.cb_syn.char_path_n\[89\] top.cb_syn.char_path_n\[92\]
+ top.cb_syn.char_path_n\[91\] net394 net292 vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07467_ _04071_ _04073_ net342 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__mux2_1
X_06418_ top.hist_data_o\[27\] _03262_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__xor2_1
X_07398_ top.findLeastValue.val2\[0\] top.findLeastValue.val1\[0\] vssd1 vssd1 vccd1
+ vccd1 _04029_ sky130_fd_sc_hd__or2_1
X_06349_ net545 _02589_ top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__mux2_1
X_09137_ net443 _02817_ _05144_ _03391_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09068_ net443 net450 _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_118_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07993__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08019_ top.findLeastValue.alternator_timer\[2\] net406 _02790_ vssd1 vssd1 vccd1
+ vccd1 _04535_ sky130_fd_sc_hd__a21oi_1
Xhold671 top.cb_syn.i\[5\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold660 top.histogram.total\[25\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11030_ clknet_leaf_57_clk _01595_ _00420_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[112\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold693 top.cw1\[6\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 top.sram_interface.write_counter_FLV\[0\] vssd1 vssd1 vccd1 vccd1 net1633
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08942__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ net895 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11863_ clknet_leaf_113_clk _02396_ _01235_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_10814_ clknet_leaf_111_clk _01408_ _00204_ vssd1 vssd1 vccd1 vccd1 top.path\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_40_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11794_ clknet_leaf_92_clk _02328_ _01166_ vssd1 vssd1 vccd1 vccd1 top.compVal\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ clknet_leaf_6_clk net1480 _00135_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10676_ clknet_leaf_107_clk _01307_ _00066_ vssd1 vssd1 vccd1 vccd1 top.path\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08608__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05995__A0 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__B2 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ clknet_leaf_84_clk _01793_ _00618_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11159_ clknet_leaf_62_clk _01724_ _00549_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[105\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07736__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05720_ top.cb_syn.char_path\[1\] net548 net539 top.cb_syn.char_path\[65\] vssd1
+ vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a22o_1
X_05651_ net467 _02714_ net307 top.hTree.node_reg\[45\] vssd1 vssd1 vccd1 vccd1 _02716_
+ sky130_fd_sc_hd__a22o_1
X_08370_ top.cb_syn.char_path_n\[19\] net198 _04747_ vssd1 vssd1 vccd1 vccd1 _01638_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_34_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05582_ top.cb_syn.char_path\[56\] net528 net312 top.cb_syn.char_path\[120\] vssd1
+ vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07321_ _03865_ _03868_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_102_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07252_ _03907_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or2_1
XANTENNA__08216__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06203_ _02510_ _03076_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__nor2_1
X_07183_ _03770_ _03771_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__and2_1
X_06134_ net1012 net166 net157 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a21o_1
XANTENNA__07424__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07975__A1 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06065_ _02529_ top.cb_syn.zero_count\[4\] _02955_ _02964_ vssd1 vssd1 vccd1 vccd1
+ _02965_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09527__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05986__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 _02569_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_2
Xfanout403 _02810_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_2
X_09824_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout394_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 net450 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_2
Xfanout425 net428 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_2
Xfanout436 _02419_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
XANTENNA__05738__A0 top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
Xfanout469 top.controller.state_reg\[1\] vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09543__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__and2_1
X_06967_ top.findLeastValue.startup net459 net288 vssd1 vssd1 vccd1 vccd1 _03668_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout561_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__and2_1
X_08706_ net1652 _04902_ _04903_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__o21a_1
X_05918_ net442 _02898_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__nor2_1
XANTENNA__06950__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06898_ top.findLeastValue.val2\[5\] net130 net120 _03654_ vssd1 vssd1 vccd1 vccd1
+ _02013_ sky130_fd_sc_hd__o22a_1
X_08637_ _04855_ _04856_ net497 vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05849_ top.sram_interface.counter_HTREE\[3\] _02868_ vssd1 vssd1 vccd1 vccd1 _02871_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ _02538_ net1541 _04788_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__mux2_1
X_07519_ _04115_ _04118_ _04110_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__mux2_1
X_08499_ net1209 top.cb_syn.char_path_n\[60\] net231 vssd1 vssd1 vccd1 vccd1 _01543_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ net805 net640 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ net828 net663 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__and2_1
XANTENNA__08622__A top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06841__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ net748 net583 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05977__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold773_A top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold490 top.path\[45\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ clknet_leaf_41_clk net1330 _00403_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07718__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07672__S _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05729__B1 _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__B2 top.cb_syn.char_path_n\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06941__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__B1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11915_ net946 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11846_ clknet_leaf_96_clk _02379_ _01218_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11777_ clknet_leaf_3_clk _00012_ _01149_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_10728_ clknet_leaf_40_clk _01359_ _00118_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[54\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06317__A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ clknet_leaf_67_clk _01290_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07406__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07870_ top.hTree.tree_reg\[23\] top.findLeastValue.sum\[23\] net281 vssd1 vssd1
+ vccd1 vccd1 _04422_ sky130_fd_sc_hd__mux2_1
XANTENNA__09363__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ top.compVal\[43\] top.findLeastValue.val1\[43\] net153 vssd1 vssd1 vccd1
+ vccd1 _03616_ sky130_fd_sc_hd__mux2_1
X_09540_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__and2_1
X_06752_ top.compVal\[14\] _02472_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _03550_
+ sky130_fd_sc_hd__a211o_1
X_09471_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__and2_1
X_05703_ top.cb_syn.char_path\[36\] net529 net310 top.cb_syn.char_path\[100\] vssd1
+ vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a22o_1
XANTENNA__09331__B1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ top.cb_syn.char_index\[4\] _04776_ _04772_ vssd1 vssd1 vccd1 vccd1 _01615_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10021__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06683_ top.compVal\[39\] _02484_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__and2_1
X_05634_ net1383 net168 _02701_ net210 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a22o_1
X_08353_ top.cb_syn.char_path_n\[28\] net373 net327 top.cb_syn.char_path_n\[26\] net176
+ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a221o_1
X_05565_ _02642_ _02643_ net465 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__o21a_1
XANTENNA__09302__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ top.cb_syn.char_path_n\[62\] net192 _04704_ vssd1 vssd1 vccd1 vccd1 _01681_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06993__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07304_ net1725 net274 net268 _03964_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
X_05496_ top.CB_read_complete top.CB_write_complete vssd1 vssd1 vccd1 vccd1 _02581_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07235_ _03904_ _03906_ _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__or3_1
XANTENNA__08842__C1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05488__D top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07757__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ _03819_ _03821_ _03838_ _03818_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o31a_1
XANTENNA__09538__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06117_ _02997_ _02999_ _03011_ _02996_ net1463 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07097_ _03771_ _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__nand2_1
X_06048_ _02450_ top.cb_syn.zeroes\[3\] top.cb_syn.zeroes\[2\] _02451_ vssd1 vssd1
+ vccd1 vccd1 _02948_ sky130_fd_sc_hd__o22a_1
Xfanout200 net202 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout244 net246 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_4
Xfanout233 _04781_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
X_09807_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__and2_1
Xfanout299 _03244_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
X_07999_ top.findLeastValue.least2\[6\] top.findLeastValue.least1\[6\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__mux2_1
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout288 _03393_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
X_09738_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__and2_1
XANTENNA__06923__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06136__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__and2_1
XANTENNA__09720__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07884__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ clknet_leaf_8_clk _02250_ _01090_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.CB_write_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11631_ clknet_leaf_28_clk _02181_ _01021_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11562_ clknet_leaf_21_clk _02127_ _00952_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ net755 net590 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ clknet_leaf_3_clk _02058_ _00883_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ net806 net641 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ net761 net596 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09183__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08667__A2 _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11935__898 vssd1 vssd1 vccd1 vccd1 _11935__898/HI net898 sky130_fd_sc_hd__conb_1
X_11829_ clknet_leaf_47_clk _02362_ _01201_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
X_05350_ top.findLeastValue.val2\[26\] vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08824__C1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07020_ _03692_ _03693_ _03694_ _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ top.WB.CPU_DAT_O\[30\] net1598 net368 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__mux2_1
XANTENNA__10016__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 top.sram_interface.init_counter\[18\] vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ net478 _04462_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_110_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07853_ net417 _04407_ _04408_ net259 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o211a_1
X_06804_ _02415_ top.findLeastValue.val2\[32\] top.findLeastValue.val2\[37\] _02410_
+ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__o2bb2a_1
X_07784_ net437 net1645 net251 top.findLeastValue.sum\[41\] _04353_ vssd1 vssd1 vccd1
+ vccd1 _01830_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09821__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06735_ top.findLeastValue.val2\[1\] top.compVal\[1\] vssd1 vssd1 vccd1 vccd1 _03533_
+ sky130_fd_sc_hd__and2b_1
X_09523_ net743 net578 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__and2_1
X_09454_ net732 net567 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__and2_1
X_06666_ _02421_ top.findLeastValue.val1\[31\] top.findLeastValue.val1\[30\] _02422_
+ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05617_ top.cb_syn.char_path\[18\] net548 net539 top.cb_syn.char_path\[82\] vssd1
+ vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a22o_1
X_08405_ top.cb_syn.char_path_n\[2\] net370 net174 net520 vssd1 vssd1 vccd1 vccd1
+ _04765_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ net1244 net228 _05270_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__o21a_1
X_08336_ top.cb_syn.char_path_n\[36\] net200 _04730_ vssd1 vssd1 vccd1 vccd1 _01655_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06597_ top.findLeastValue.startup _02562_ net288 vssd1 vssd1 vccd1 vccd1 _02055_
+ sky130_fd_sc_hd__a21o_1
X_05548_ top.histogram.sram_out\[30\] net360 net411 top.hTree.node_reg\[30\] vssd1
+ vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ top.cb_syn.char_path_n\[71\] net376 net333 top.cb_syn.char_path_n\[69\] net178
+ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a221o_1
X_05479_ net31 net413 net362 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 _02379_
+ sky130_fd_sc_hd__o22a_1
X_08198_ net1765 net201 _04661_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__o21a_1
XANTENNA__05644__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _03733_ _03893_ _03736_ _03735_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_76_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07149_ top.findLeastValue.val2\[2\] top.findLeastValue.val1\[2\] vssd1 vssd1 vccd1
+ vccd1 _03825_ sky130_fd_sc_hd__nand2_1
XANTENNA__08594__A1 top.cb_syn.char_path_n\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07397__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10160_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__and2_1
X_10091_ net834 net669 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__and2_1
XANTENNA__05735__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10993_ clknet_leaf_60_clk _01558_ _00383_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11614_ clknet_leaf_22_clk _02164_ _01004_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08781__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08806__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11545_ clknet_leaf_72_clk _02110_ _00935_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08821__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05635__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11476_ clknet_leaf_97_clk _02041_ _00866_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[33\]
+ sky130_fd_sc_hd__dfstp_1
X_10427_ net818 net653 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09906__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ net720 net555 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10915__918 vssd1 vssd1 vccd1 vccd1 net918 _10915__918/LO sky130_fd_sc_hd__conb_1
X_10289_ net833 net668 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__and2_1
XANTENNA__07793__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07860__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09298__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06520_ net1611 _03339_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__nor2_1
X_06451_ top.hist_data_o\[13\] _03253_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nor2_1
X_05402_ top.findLeastValue.least2\[2\] vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__inv_2
X_09170_ net488 net524 _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_60_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06382_ top.hist_data_o\[5\] top.hist_data_o\[4\] vssd1 vssd1 vccd1 vccd1 _03247_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05333_ top.cb_syn.count\[3\] vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__inv_2
X_08121_ _04560_ _04605_ _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nor3_2
XFILLER_0_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ top.cb_syn.char_path_n\[2\] _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_78_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05626__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ net407 net287 net133 vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__and3_2
XANTENNA__07379__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08954_ top.WB.CPU_DAT_O\[14\] net1398 net321 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__mux2_1
X_07905_ top.hTree.tree_reg\[16\] top.findLeastValue.sum\[16\] net286 vssd1 vssd1
+ vccd1 vccd1 _04450_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout474_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ net1442 top.WB.CPU_DAT_O\[17\] net302 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__mux2_1
XANTENNA__05782__C net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ top.findLeastValue.sum\[30\] _04394_ net390 vssd1 vssd1 vccd1 vccd1 _04395_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07551__A2 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05562__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net478 _04338_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout641_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09551__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05562__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09506_ net732 net567 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__and2_1
XANTENNA__07839__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06718_ _03509_ _03515_ _02406_ top.findLeastValue.val2\[45\] vssd1 vssd1 vccd1 vccd1
+ _03516_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07698_ net473 _04281_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__or2_1
X_06649_ _02435_ top.findLeastValue.val1\[11\] vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__and2_1
X_09437_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ net1405 net222 _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a22o_1
XANTENNA__05865__A2 _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ top.cb_syn.char_path_n\[45\] net381 net338 top.cb_syn.char_path_n\[43\] net184
+ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09299_ net504 _05241_ _05242_ _05240_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05617__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ clknet_leaf_82_clk _01895_ _00720_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11261_ clknet_leaf_81_clk _01826_ _00651_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_11192_ clknet_leaf_27_clk _01757_ _00582_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10212_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__and2_1
X_10143_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10074_ net786 net621 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__and2_1
XANTENNA_input35_A gpio_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ clknet_leaf_37_clk _01541_ _00366_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05608__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11528_ clknet_leaf_85_clk _02093_ _00918_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold308 top.path\[107\] vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 top.hTree.nulls\[46\] vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
X_11459_ clknet_leaf_101_clk _02024_ _00849_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08558__A1 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07855__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05951_ top.compVal\[10\] net160 net143 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 _02227_ sky130_fd_sc_hd__a22o_1
X_08670_ top.cb_syn.i\[1\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05882_ net1689 top.WB.CPU_DAT_O\[16\] net351 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05544__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ net1417 _04219_ _04212_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ top.cb_syn.char_path_n\[26\] top.cb_syn.char_path_n\[25\] top.cb_syn.char_path_n\[28\]
+ top.cb_syn.char_path_n\[27\] net397 net292 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__mux4_1
XANTENNA__05544__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05404__A top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950__913 vssd1 vssd1 vccd1 vccd1 _11950__913/HI net913 sky130_fd_sc_hd__conb_1
X_06503_ top.histogram.total\[20\] top.histogram.total\[19\] _03335_ vssd1 vssd1 vccd1
+ vccd1 _03336_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07483_ _04081_ _04086_ net393 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__mux2_1
X_09222_ _03372_ _05197_ _03376_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_char_added
+ sky130_fd_sc_hd__o21ai_1
X_06434_ net1145 _03288_ _03243_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_86_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06365_ _03019_ _03229_ _03231_ top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1
+ _03232_ sky130_fd_sc_hd__o211a_1
X_09153_ _05155_ _05156_ net536 vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08104_ top.cb_syn.num_lefts\[3\] _04592_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout222_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05316_ top.compVal\[16\] vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06296_ top.cw1\[4\] _03071_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__xor2_1
X_09084_ net460 top.sram_interface.word_cnt\[2\] net356 top.hTree.write_HT_fin _05109_
+ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a221o_1
Xhold820 top.cb_syn.char_path_n\[126\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
X_08035_ top.cb_syn.setup net463 top.cb_syn.curr_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _04547_ sky130_fd_sc_hd__and3_1
Xhold831 top.cb_syn.char_path_n\[11\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold853 top.compVal\[2\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 top.compVal\[6\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_95_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08937_ top.WB.CPU_DAT_O\[31\] net1393 net319 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08596__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ net513 _02808_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__nand2_1
X_07819_ net435 net1313 net249 top.findLeastValue.sum\[34\] _04381_ vssd1 vssd1 vccd1
+ vccd1 _01823_ sky130_fd_sc_hd__a221o_1
X_08799_ top.path\[68\] net404 _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ clknet_leaf_116_clk _01424_ _00220_ vssd1 vssd1 vccd1 vccd1 top.path\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10761_ clknet_leaf_9_clk _00042_ _00151_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ clknet_leaf_108_clk _01323_ _00082_ vssd1 vssd1 vccd1 vccd1 top.path\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05968__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ clknet_leaf_41_clk _01878_ _00703_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11244_ clknet_leaf_77_clk net1396 _00634_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08635__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11175_ clknet_leaf_37_clk _01740_ _00565_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05774__B2 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ net819 net654 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__and2_1
XANTENNA__09903__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ net719 net554 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__and2_1
X_10959_ clknet_leaf_62_clk _01524_ _00349_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11910__941 vssd1 vssd1 vccd1 vccd1 net941 _11910__941/LO sky130_fd_sc_hd__conb_1
XANTENNA__08779__A1 _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06150_ _02417_ _03026_ net207 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06081_ top.cb_syn.cb_length\[0\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _02981_
+ sky130_fd_sc_hd__xnor2_1
Xhold105 top.cb_syn.char_path\[23\] vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 top.cb_syn.char_path\[46\] vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 top.cb_syn.char_path\[62\] vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 top.cb_syn.char_path\[63\] vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 top.path\[7\] vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
X_09840_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
Xfanout607 net608 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_2
Xfanout618 net621 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ net788 net623 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__and2_1
X_06983_ _03089_ _03185_ _03675_ _03667_ net486 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05765__B2 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05934_ top.compVal\[27\] net158 net145 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 _02244_ sky130_fd_sc_hd__a22o_1
X_08722_ top.sram_interface.TRN_counter\[1\] top.sram_interface.TRN_counter\[0\] top.sram_interface.TRN_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout172_A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ top.cb_syn.end_cnt\[4\] _04790_ _04866_ top.cb_syn.end_cnt\[5\] vssd1 vssd1
+ vccd1 vccd1 _04870_ sky130_fd_sc_hd__o31a_1
X_05865_ net448 _02562_ net411 top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 _02284_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08584_ net497 _04803_ _02541_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a21o_1
X_07604_ top.cb_syn.pulse_first net521 _02889_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05796_ net542 _02577_ _02800_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_37_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ top.cb_syn.char_path_n\[94\] top.cb_syn.char_path_n\[93\] top.cb_syn.char_path_n\[96\]
+ top.cb_syn.char_path_n\[95\] net394 net292 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout437_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07466_ _04054_ _04072_ _04049_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__mux2_1
X_09205_ top.header_synthesis.start _03375_ _03372_ vssd1 vssd1 vccd1 vccd1 _05185_
+ sky130_fd_sc_hd__nor3b_1
X_06417_ net1118 _03278_ net301 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ _03831_ net271 _04028_ net277 net1749 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06348_ top.cb_syn.max_index\[2\] _03102_ _03104_ top.hTree.nullSumIndex\[1\] vssd1
+ vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a22o_1
X_09136_ top.findLeastValue.histo_index\[8\] _02575_ _02816_ top.sram_interface.zero_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_17_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06279_ top.sram_interface.init_counter\[5\] _03021_ vssd1 vssd1 vccd1 vccd1 _03150_
+ sky130_fd_sc_hd__nor2_1
X_09067_ _03013_ _05094_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nor2_2
X_08018_ top.findLeastValue.alternator_timer\[1\] top.findLeastValue.alternator_timer\[0\]
+ _03666_ top.findLeastValue.alternator_timer\[2\] vssd1 vssd1 vccd1 vccd1 _04534_
+ sky130_fd_sc_hd__a31o_1
Xhold672 top.hist_data_o\[12\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 _01800_ vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 top.hist_addr\[3\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 top.hTree.tree_reg\[41\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 top.hist_data_o\[10\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__and2_1
XANTENNA__09723__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08155__C1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ net894 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__08170__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11862_ clknet_leaf_112_clk _02395_ _01234_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_10813_ clknet_leaf_25_clk _00011_ _00203_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11793_ clknet_leaf_92_clk _02327_ _01165_ vssd1 vssd1 vccd1 vccd1 top.compVal\[42\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_15_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ clknet_leaf_6_clk _00034_ _00134_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07681__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ clknet_leaf_109_clk _01306_ _00065_ vssd1 vssd1 vccd1 vccd1 top.path\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08608__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ clknet_leaf_84_clk _01792_ _00617_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11158_ clknet_leaf_64_clk _01723_ _00548_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[104\]
+ sky130_fd_sc_hd__dfrtp_2
X_10109_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__and2_1
XANTENNA__06944__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11089_ clknet_leaf_63_clk _01654_ _00479_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_05650_ _02418_ net356 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__and2_1
X_05581_ top.cb_syn.char_path\[24\] top.sram_interface.word_cnt\[0\] net538 top.cb_syn.char_path\[88\]
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07320_ net268 _03974_ _03975_ net274 net1669 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06484__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07251_ _03910_ _03924_ _03908_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__o21ai_1
X_06202_ top.cw2\[1\] top.cw2\[0\] vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__nand2_1
X_07182_ top.findLeastValue.val2\[15\] top.findLeastValue.val1\[15\] _03796_ _03856_
+ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a221oi_4
X_06133_ net1033 net166 net157 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06064_ _02532_ top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__or2_1
Xfanout404 _02810_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_4
X_09823_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__and2_1
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_2
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_2
Xfanout415 _02568_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_2
Xfanout426 net428 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_2
Xfanout459 top.controller.state_reg\[2\] vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06935__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__and2_1
X_06966_ _02793_ net287 vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__and2_1
X_09685_ net863 net698 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__and2_1
X_08705_ net1430 _04903_ _04905_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05917_ net439 net543 net460 vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__and3_1
X_06897_ top.compVal\[5\] top.findLeastValue.val1\[5\] net154 vssd1 vssd1 vccd1 vccd1
+ _03654_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout554_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08152__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08636_ top.cb_syn.char_path_n\[35\] top.cb_syn.char_path_n\[36\] top.cb_syn.char_path_n\[39\]
+ top.cb_syn.char_path_n\[40\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_68_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
X_05848_ _02867_ _02861_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07360__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _04202_ _04771_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_81_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout721_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05779_ net513 top.translation.totalEn _02808_ top.TRN_sram_complete vssd1 vssd1
+ vccd1 vccd1 _02809_ sky130_fd_sc_hd__or4bb_1
X_07518_ _04116_ _04117_ net289 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__mux2_1
X_08498_ net1295 top.cb_syn.char_path_n\[61\] net230 vssd1 vssd1 vccd1 vccd1 _01544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ top.dut.bits_in_buf\[1\] top.dut.bits_in_buf\[2\] net393 vssd1 vssd1 vccd1
+ vccd1 _04057_ sky130_fd_sc_hd__and3_1
X_10460_ net766 net601 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ net453 top.histogram.state\[1\] net1786 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_79_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05738__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ net735 net570 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold480 top.hTree.tree_reg\[24\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ clknet_leaf_39_clk _01577_ _00402_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[94\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold491 top.path\[17\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06926__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05729__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__C1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06154__A1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11914_ net945 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XANTENNA__08784__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
X_11845_ clknet_leaf_96_clk _02378_ _01217_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11776_ clknet_leaf_75_clk _02315_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10727_ clknet_leaf_25_clk _01358_ _00117_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05502__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ clknet_leaf_67_clk _01289_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08813__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ net745 net580 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06820_ top.findLeastValue.val2\[44\] net129 net119 _03615_ vssd1 vssd1 vccd1 vccd1
+ _02052_ sky130_fd_sc_hd__o22a_1
X_06751_ _02472_ top.compVal\[14\] _02434_ top.findLeastValue.val2\[15\] vssd1 vssd1
+ vccd1 vccd1 _03549_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05702_ top.cb_syn.char_path\[4\] net549 net541 top.cb_syn.char_path\[68\] vssd1
+ vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a22o_1
X_09470_ net837 net672 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_75_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
X_06682_ top.compVal\[40\] _02483_ _02484_ top.compVal\[39\] vssd1 vssd1 vccd1 vccd1
+ _03480_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08421_ top.cb_syn.h_element\[59\] top.cb_syn.h_element\[50\] net517 vssd1 vssd1
+ vccd1 vccd1 _04776_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05633_ top.hTree.node_reg\[16\] net409 _02699_ _02700_ vssd1 vssd1 vccd1 vccd1 _02701_
+ sky130_fd_sc_hd__a211o_1
X_08352_ top.cb_syn.char_path_n\[28\] net190 _04738_ vssd1 vssd1 vccd1 vccd1 _01647_
+ sky130_fd_sc_hd__o21a_1
X_05564_ top.cb_syn.char_path\[27\] top.sram_interface.word_cnt\[0\] net309 top.cb_syn.char_path\[123\]
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ top.cb_syn.char_path_n\[63\] net370 net328 top.cb_syn.char_path_n\[61\] net174
+ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a221o_1
X_05495_ top.CB_read_complete top.CB_write_complete vssd1 vssd1 vccd1 vccd1 _02580_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08842__B1 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07303_ _03741_ _03960_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__xnor2_1
X_07234_ _03908_ _03909_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout135_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07165_ _03817_ _03819_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout302_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06116_ _02451_ _02998_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07096_ top.findLeastValue.val2\[16\] top.findLeastValue.val1\[16\] vssd1 vssd1 vccd1
+ vccd1 _03772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06047_ _02451_ top.cb_syn.zeroes\[2\] top.cb_syn.zeroes\[1\] _02452_ _02946_ vssd1
+ vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05959__B2 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
Xfanout223 _05253_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout671_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 net259 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06908__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 _04111_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_4
X_09806_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__and2_1
Xfanout267 _04251_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_4
X_07998_ top.hTree.state\[6\] top.hTree.state\[3\] vssd1 vssd1 vccd1 vccd1 _04523_
+ sky130_fd_sc_hd__nor2_2
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
X_09737_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__and2_1
X_06949_ top.findLeastValue.val1\[8\] net135 net113 net1687 vssd1 vssd1 vccd1 vccd1
+ _01969_ sky130_fd_sc_hd__o22a_1
XANTENNA__07559__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07802__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__and2_1
X_08619_ top.cb_syn.char_path_n\[1\] top.cb_syn.char_path_n\[2\] top.cb_syn.char_path_n\[5\]
+ top.cb_syn.char_path_n\[6\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__mux4_1
XANTENNA__07884__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__and2_1
X_11630_ clknet_leaf_29_clk _02180_ _01020_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11561_ clknet_leaf_21_clk _02126_ _00951_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05647__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512_ net757 net592 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__and2_1
XANTENNA__08633__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ clknet_leaf_4_clk _02057_ _00882_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_HG
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10443_ net807 net642 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__and2_1
XANTENNA__08597__C1 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ net760 net595 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08349__C1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10403__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_57_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08747__S0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ clknet_leaf_67_clk _02361_ _01200_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09077__B1 top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05638__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ clknet_leaf_47_clk _02298_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06850__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08588__C1 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06041__C_N top.WB.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08970_ top.WB.CPU_DAT_O\[31\] net550 net368 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__mux2_1
XANTENNA__09001__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ top.hTree.tree_reg\[13\] top.findLeastValue.sum\[13\] net267 vssd1 vssd1
+ vccd1 vccd1 _04463_ sky130_fd_sc_hd__mux2_1
XANTENNA__08355__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ net471 _04406_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__or2_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__dlymetal6s2s_1
X_06803_ _02413_ top.findLeastValue.val2\[34\] top.findLeastValue.val2\[33\] _02414_
+ _03522_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o221a_1
XANTENNA__08760__C1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
X_07783_ net420 _04351_ _04352_ net262 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o211a_1
X_09522_ net745 net580 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__and2_1
XANTENNA__09821__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06734_ top.compVal\[9\] _02475_ _02476_ top.compVal\[8\] vssd1 vssd1 vccd1 vccd1
+ _03532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout252_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__and2_1
X_06665_ top.compVal\[27\] _02490_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__nor2_1
X_08404_ top.cb_syn.char_path_n\[2\] net197 _04764_ vssd1 vssd1 vccd1 vccd1 _01621_
+ sky130_fd_sc_hd__o21a_1
X_05616_ net1365 net171 _02686_ net211 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a22o_1
X_09384_ net1212 _02851_ net220 _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a211o_1
X_08335_ top.cb_syn.char_path_n\[37\] net379 net336 top.cb_syn.char_path_n\[35\] net182
+ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a221o_1
X_06596_ _02562_ net288 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__nor2_1
XANTENNA__05629__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05547_ _02627_ _02628_ net465 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_22_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08266_ top.cb_syn.char_path_n\[71\] net202 _04695_ vssd1 vssd1 vccd1 vccd1 _01690_
+ sky130_fd_sc_hd__o21a_1
X_05478_ net32 net415 net364 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 _02380_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09549__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ top.cb_syn.char_path_n\[106\] net381 net337 top.cb_syn.char_path_n\[104\]
+ net183 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07217_ _02462_ _02487_ _03881_ _03891_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__o221a_1
X_07148_ top.findLeastValue.val2\[3\] top.findLeastValue.val1\[3\] vssd1 vssd1 vccd1
+ vccd1 _03824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ top.findLeastValue.val2\[27\] top.findLeastValue.val1\[27\] vssd1 vssd1 vccd1
+ vccd1 _03755_ sky130_fd_sc_hd__and2_1
X_10090_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__and2_1
XANTENNA__08346__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08729__S0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10992_ clknet_leaf_61_clk _01557_ _00382_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06847__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11613_ clknet_leaf_22_clk _02163_ _01003_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08806__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11544_ clknet_leaf_72_clk _02109_ _00934_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06832__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11475_ clknet_leaf_97_clk _02040_ _00865_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[32\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09178__B top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10426_ net821 net656 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09906__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357_ net718 net553 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__and2_1
X_10288_ net833 net668 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08742__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09298__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06450_ net298 _03256_ _03296_ _03297_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__o31ai_1
X_05401_ top.findLeastValue.least2\[3\] vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06381_ top.hist_data_o\[3\] top.hist_data_o\[2\] top.hist_data_o\[1\] top.hist_data_o\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05332_ top.cb_syn.count\[4\] vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__inv_2
X_08120_ _04202_ _04586_ _04610_ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_60_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08051_ top.cb_syn.char_path_n\[1\] _04201_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07002_ net1742 net142 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08953_ top.WB.CPU_DAT_O\[15\] net1381 net321 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__mux2_1
XANTENNA__07784__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ net438 net1443 net252 top.findLeastValue.sum\[17\] _04449_ vssd1 vssd1 vccd1
+ vccd1 _01806_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08884_ net1069 top.WB.CPU_DAT_O\[18\] net302 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__mux2_1
XANTENNA__05782__D net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout467_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07000__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ top.hTree.tree_reg\[30\] top.findLeastValue.sum\[30\] net282 vssd1 vssd1
+ vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
XANTENNA__05562__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ top.findLeastValue.sum\[44\] _04338_ net392 vssd1 vssd1 vccd1 vccd1 _04339_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09505_ net732 net567 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__and2_1
XANTENNA__07839__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06717_ _03512_ _03513_ _03514_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a21oi_1
X_07697_ net473 _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__nand2_1
X_09436_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__and2_1
X_06648_ _02435_ top.findLeastValue.val1\[11\] top.findLeastValue.val1\[10\] _02436_
+ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__o22a_1
X_06579_ top.header_synthesis.count\[0\] _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__or2_1
X_09367_ top.hTree.nulls\[48\] net398 net229 vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ top.cb_syn.char_path_n\[45\] net200 _04721_ vssd1 vssd1 vccd1 vccd1 _01664_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09298_ top.histogram.total\[0\] net403 net323 top.histogram.total\[1\] net429 vssd1
+ vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__o221a_1
X_08249_ top.cb_syn.char_path_n\[80\] net385 net340 top.cb_syn.char_path_n\[78\] net188
+ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a221o_1
XANTENNA__08911__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ clknet_leaf_80_clk _01825_ _00650_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_11191_ clknet_leaf_27_clk _01756_ _00581_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10211_ net824 net659 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__and2_1
X_10142_ net735 net570 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__and2_1
X_10073_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07246__B _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07527__A0 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07961__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ clknet_leaf_37_clk _01540_ _00365_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05454__C_N top.WB.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05510__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ clknet_leaf_80_clk _02092_ _00917_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06325__B top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output96_A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 top.hTree.nulls\[49\] vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
X_11458_ clknet_leaf_79_clk _02023_ _00848_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[15\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__07766__A0 top.findLeastValue.sum\[44\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11389_ clknet_leaf_14_clk _01954_ _00779_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10409_ net742 net577 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__and2_1
XANTENNA__07871__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05950_ top.compVal\[11\] net160 net143 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 _02228_ sky130_fd_sc_hd__a22o_1
X_05881_ net1663 top.WB.CPU_DAT_O\[17\] net351 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07620_ top.cb_syn.max_index\[6\] _04181_ _04215_ _04218_ vssd1 vssd1 vccd1 vccd1
+ _04219_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_109_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ top.cb_syn.char_path_n\[30\] top.cb_syn.char_path_n\[29\] top.cb_syn.char_path_n\[32\]
+ top.cb_syn.char_path_n\[31\] net397 net292 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__mux4_1
XANTENNA__05544__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06502_ top.histogram.total\[18\] top.histogram.total\[17\] _03334_ vssd1 vssd1 vccd1
+ vccd1 _03335_ sky130_fd_sc_hd__and3_1
XANTENNA__08494__A1 top.cb_syn.char_path_n\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07482_ top.dut.bit_buf\[3\] net41 net714 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__mux2_1
X_09221_ net490 net1674 vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nor2_1
X_06433_ top.hist_data_o\[21\] _03269_ _03273_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__o21ba_1
X_06364_ _03097_ _03230_ top.histogram.init vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__a21o_1
X_09152_ net442 net462 net451 top.sram_interface.TRN_counter\[2\] _05096_ vssd1 vssd1
+ vccd1 vccd1 _05156_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08103_ top.cb_syn.num_lefts\[4\] _04589_ _04590_ _04601_ vssd1 vssd1 vccd1 vccd1
+ _01759_ sky130_fd_sc_hd__a22o_1
X_05315_ top.compVal\[17\] vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__inv_2
X_06295_ net486 _02787_ _03090_ _03164_ _02601_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a221o_1
X_09083_ net451 _05108_ top.sram_interface.word_cnt\[9\] vssd1 vssd1 vccd1 vccd1 _05109_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout215_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold821 top.cb_syn.char_path_n\[108\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
X_08034_ top.cb_syn.setup net463 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__nand2_1
XANTENNA__08731__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold810 top.sram_interface.counter_HTREE\[3\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 top.cb_syn.i\[4\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 top.cb_syn.char_path_n\[94\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 top.cb_syn.char_path_n\[94\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05480__B2 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout584_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__and2_1
X_08936_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__inv_2
XANTENNA__07781__S _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ _02808_ _02813_ net513 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout751_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ net418 _04379_ _04380_ net260 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o211a_1
X_08798_ top.path\[69\] net324 _04986_ net426 _02547_ vssd1 vssd1 vccd1 vccd1 _04987_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_84_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07749_ top.hTree.tree_reg\[47\] top.findLeastValue.least2\[1\] net281 vssd1 vssd1
+ vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
X_10760_ clknet_leaf_9_clk _00041_ _00150_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_09419_ net965 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__clkbuf_1
X_10691_ clknet_leaf_108_clk _01322_ _00081_ vssd1 vssd1 vccd1 vccd1 top.path\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11312_ clknet_leaf_13_clk _01877_ _00702_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07956__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ clknet_leaf_77_clk net1351 _00633_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05471__B2 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ clknet_leaf_37_clk _01739_ _00564_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[120\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06161__A top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05759__C1 _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05774__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ net820 net655 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__and2_1
X_10056_ net719 net554 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__and2_1
XANTENNA__08173__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ clknet_leaf_65_clk _01523_ _00348_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ clknet_leaf_26_clk top.header_synthesis.next_write_char_path _00279_ vssd1
+ vssd1 vccd1 vccd1 top.header_synthesis.write_char_path sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06080_ top.cb_syn.cb_length\[0\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _02980_
+ sky130_fd_sc_hd__nand2b_1
Xhold117 top.cb_syn.char_path\[28\] vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07866__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold106 top.path\[31\] vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold128 top.cb_syn.char_path\[120\] vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top.cb_syn.char_path\[1\] vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05462__B2 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout608 net611 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout619 net621 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__and2_1
X_06982_ _03669_ _03675_ _03678_ _03667_ net484 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a32o_1
XANTENNA__05765__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05933_ top.compVal\[28\] net159 net144 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 _02245_ sky130_fd_sc_hd__a22o_1
X_08721_ net304 _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__nor2_1
X_08652_ _04867_ _04869_ top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__mux2_1
X_07603_ net489 _02895_ net524 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__or3b_1
XANTENNA__07911__A0 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05864_ net1476 _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_37_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ top.cb_syn.char_path_n\[75\] top.cb_syn.char_path_n\[76\] top.cb_syn.char_path_n\[79\]
+ top.cb_syn.char_path_n\[80\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout165_A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05795_ net1531 net454 _02594_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07534_ _04130_ _04133_ _04110_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ top.dut.bit_buf\[6\] net35 net713 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout332_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06416_ _03263_ _03277_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09204_ _05184_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07690__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07396_ _03828_ _03829_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nand2b_1
X_06347_ _03019_ _03213_ _03214_ top.histogram.init net454 vssd1 vssd1 vccd1 vccd1
+ _03215_ sky130_fd_sc_hd__o221a_1
X_09135_ _02862_ _05142_ net304 _02585_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or4b_1
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06278_ _03099_ _03148_ _02416_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__o21ai_1
X_09066_ net439 top.sram_interface.word_cnt\[9\] _05094_ _05095_ net1581 vssd1 vssd1
+ vccd1 vccd1 _00049_ sky130_fd_sc_hd__a32o_1
XANTENNA__07776__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout799_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ _02562_ _04533_ _04532_ net287 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__o211a_1
Xhold662 _01329_ vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 top.histogram.total\[15\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 top.histogram.total\[2\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 top.hist_data_o\[30\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 top.findLeastValue.sum\[20\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 top.translation.write_fin vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
X_09968_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__and2_1
X_08919_ _05061_ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__nor2_1
X_09899_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__and2_1
X_11930_ net893 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
X_11892__923 vssd1 vssd1 vccd1 vccd1 net923 _11892__923/LO sky130_fd_sc_hd__conb_1
XANTENNA__10231__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ clknet_leaf_112_clk _02394_ _01233_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_10812_ clknet_leaf_26_clk _00010_ _00202_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.pulse_first_n
+ sky130_fd_sc_hd__dfrtp_1
X_11792_ clknet_leaf_92_clk _02326_ _01164_ vssd1 vssd1 vccd1 vccd1 top.compVal\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06855__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10743_ clknet_leaf_6_clk _00033_ _00133_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10674_ clknet_leaf_110_clk _01305_ _00064_ vssd1 vssd1 vccd1 vccd1 top.path\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07969__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11226_ clknet_leaf_83_clk _01791_ _00616_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07197__A1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ clknet_leaf_64_clk _01722_ _00547_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[103\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08933__A2 _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09406__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ net810 net645 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__and2_1
X_11088_ clknet_leaf_63_clk _01653_ _00478_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[34\]
+ sky130_fd_sc_hd__dfrtp_2
X_10039_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05580_ net1447 net168 _02656_ net210 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07250_ _03895_ _03903_ _03913_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a21boi_2
X_06201_ top.findLeastValue.histo_index\[8\] _02501_ net534 _02575_ _02603_ vssd1
+ vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__a41o_1
XANTENNA__06880__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ top.findLeastValue.val2\[14\] top.findLeastValue.val1\[14\] _03794_ vssd1
+ vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__and3_1
X_06132_ net1036 net166 net157 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_57_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06063_ _02526_ top.cb_syn.zero_count\[7\] vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__and2_1
XANTENNA__07188__A1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 _02810_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_2
X_09822_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__and2_1
X_11880__882 vssd1 vssd1 vccd1 vccd1 _11880__882/HI net882 sky130_fd_sc_hd__conb_1
Xfanout438 _02419_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_4
Xfanout416 _02568_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_2
X_09753_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__and2_1
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
X_08704_ top.header_synthesis.count\[7\] top.header_synthesis.count\[6\] top.header_synthesis.count\[5\]
+ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout282_A _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06965_ _02562_ net287 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__nand2_1
X_09684_ net862 net697 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__and2_1
X_05916_ _02888_ _02891_ _02897_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__and3b_1
X_06896_ top.findLeastValue.val2\[6\] net129 net121 _03653_ vssd1 vssd1 vccd1 vccd1
+ _02014_ sky130_fd_sc_hd__o22a_1
X_08635_ top.cb_syn.char_path_n\[33\] top.cb_syn.char_path_n\[34\] top.cb_syn.char_path_n\[37\]
+ top.cb_syn.char_path_n\[38\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_68_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05847_ _02861_ _02868_ _02867_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout547_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ _02538_ net515 _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__o21a_1
X_11917__948 vssd1 vssd1 vccd1 vccd1 net948 _11917__948/LO sky130_fd_sc_hd__conb_1
X_07517_ top.cb_syn.char_path_n\[98\] top.cb_syn.char_path_n\[97\] top.cb_syn.char_path_n\[100\]
+ top.cb_syn.char_path_n\[99\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_81_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05778_ net423 net452 net36 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__and3_1
X_08497_ net1089 top.cb_syn.char_path_n\[62\] net230 vssd1 vssd1 vccd1 vccd1 _01545_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout714_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07448_ _04052_ _04055_ net342 vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__mux2_1
XANTENNA__08860__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ net1743 net278 _04017_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a21o_1
X_09118_ _02417_ top.histogram.eof_n net360 _05122_ _05131_ vssd1 vssd1 vccd1 vccd1
+ _00032_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ net769 net604 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09049_ top.WB.CPU_DAT_O\[1\] net1471 net316 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold470 net91 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _01813_ vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ clknet_leaf_38_clk net1293 _00401_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[93\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold492 top.hTree.tree_reg\[17\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05729__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net944 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ clknet_leaf_113_clk _02377_ _01216_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_11775_ clknet_leaf_41_clk _02314_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10726_ clknet_leaf_17_clk _01357_ _00116_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05502__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10657_ clknet_leaf_66_clk _01288_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06862__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10588_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08367__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ clknet_leaf_107_clk _01774_ _00599_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_06750_ _02434_ top.findLeastValue.val2\[15\] vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09331__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05701_ net1285 net170 _02757_ net209 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a22o_1
X_06681_ _02410_ top.findLeastValue.val1\[37\] top.findLeastValue.val1\[36\] _02411_
+ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__a22o_1
X_08420_ top.cb_syn.char_index\[5\] _04775_ _04772_ vssd1 vssd1 vccd1 vccd1 _01616_
+ sky130_fd_sc_hd__mux2_1
X_05632_ top.histogram.sram_out\[16\] net358 net355 top.hTree.node_reg\[48\] vssd1
+ vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ top.cb_syn.char_path_n\[29\] net369 net327 top.cb_syn.char_path_n\[27\] net173
+ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a221o_1
X_05563_ top.cb_syn.char_path\[91\] net537 net532 top.cb_syn.char_path\[59\] vssd1
+ vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
X_08282_ net1745 net193 _04703_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_63_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05494_ top.FLV_done _02576_ _02577_ net361 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08842__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07302_ net268 _03962_ _03963_ net274 net1705 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a32o_1
X_07233_ top.findLeastValue.val2\[42\] top.findLeastValue.val1\[42\] vssd1 vssd1 vccd1
+ vccd1 _03909_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout128_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ _03821_ _03838_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__or2_1
X_06115_ _02997_ _03001_ _03010_ _02996_ net1438 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a32o_1
X_07095_ top.findLeastValue.val2\[17\] top.findLeastValue.val1\[17\] vssd1 vssd1 vccd1
+ vccd1 _03771_ sky130_fd_sc_hd__nand2_1
X_06046_ _02452_ top.cb_syn.zeroes\[1\] top.cb_syn.zeroes\[0\] _02453_ vssd1 vssd1
+ vccd1 vccd1 _02946_ sky130_fd_sc_hd__o211a_1
Xfanout202 net206 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
Xfanout213 _02616_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
X_09805_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout257 net259 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
X_07997_ _02846_ _04257_ _04518_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__o21a_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_A net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 net270 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
Xfanout279 _03719_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
XANTENNA__05592__B1 _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__and2_1
X_06948_ top.findLeastValue.val1\[9\] net136 net113 net1768 vssd1 vssd1 vccd1 vccd1
+ _01970_ sky130_fd_sc_hd__o22a_1
X_09667_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__and2_1
XANTENNA__06136__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _02541_ _04837_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout831_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ top.compVal\[14\] top.findLeastValue.val1\[14\] net154 vssd1 vssd1 vccd1
+ vccd1 _03645_ sky130_fd_sc_hd__mux2_1
X_09598_ net742 net577 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__and2_1
X_08549_ net1321 top.cb_syn.char_path_n\[10\] net240 vssd1 vssd1 vccd1 vccd1 _01493_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09086__B2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05895__A1 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ clknet_leaf_21_clk _02125_ _00950_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10511_ net757 net592 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__and2_1
XANTENNA__06844__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ clknet_leaf_26_clk _02056_ _00881_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.bit1
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ net807 net642 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ net760 net595 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10403__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05583__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout791 net794 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_2
Xfanout780 net795 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08747__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05886__A1 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ clknet_leaf_66_clk _02360_ _01199_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11758_ clknet_leaf_106_clk _00018_ _01148_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10709_ clknet_leaf_74_clk _01340_ _00099_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ clknet_leaf_76_clk _02239_ _01079_ vssd1 vssd1 vccd1 vccd1 top.compVal\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07260__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ top.hTree.tree_reg\[13\] top.findLeastValue.sum\[13\] net285 vssd1 vssd1
+ vccd1 vccd1 _04462_ sky130_fd_sc_hd__mux2_1
X_07851_ top.hTree.tree_reg\[27\] top.findLeastValue.sum\[27\] net265 vssd1 vssd1
+ vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
XANTENNA__07563__A1 top.cb_syn.char_path_n\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07782_ net479 _04350_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__or2_1
X_06802_ _02411_ top.findLeastValue.val2\[36\] top.findLeastValue.val2\[35\] _02412_
+ _03521_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o221a_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05574__B1 _02651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__and2_1
X_06733_ top.compVal\[9\] _02475_ _03528_ _03530_ vssd1 vssd1 vccd1 vccd1 _03531_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_65_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06664_ _02422_ top.findLeastValue.val1\[30\] top.findLeastValue.val1\[29\] _02423_
+ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__o22ai_2
X_09452_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__and2_1
X_08403_ top.cb_syn.char_path_n\[3\] net376 net332 top.cb_syn.char_path_n\[1\] net179
+ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a221o_1
X_05615_ top.hTree.node_reg\[51\] net354 _02684_ _02685_ vssd1 vssd1 vccd1 vccd1 _02686_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__05877__A1 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ top.findLeastValue.least2\[8\] net390 net265 top.hTree.tree_reg\[54\] net401
+ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__o221a_1
X_06595_ _02865_ _03392_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__or2_2
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout245_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05546_ top.cb_syn.char_path\[62\] net528 net309 top.cb_syn.char_path\[126\] vssd1
+ vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
X_08334_ top.cb_syn.char_path_n\[37\] net200 _04729_ vssd1 vssd1 vccd1 vccd1 _01656_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06826__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08265_ top.cb_syn.char_path_n\[72\] net379 net336 top.cb_syn.char_path_n\[70\] net182
+ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05477_ net33 net413 net363 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 _02381_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__B net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08196_ top.cb_syn.char_path_n\[106\] net203 _04660_ vssd1 vssd1 vccd1 vccd1 _01725_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07216_ _03875_ _03878_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or2_1
XANTENNA__08579__B1 _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ top.findLeastValue.val2\[3\] top.findLeastValue.val1\[3\] vssd1 vssd1 vccd1
+ vccd1 _03823_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout781_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ top.findLeastValue.val2\[27\] top.findLeastValue.val1\[27\] vssd1 vssd1 vccd1
+ vccd1 _03754_ sky130_fd_sc_hd__nor2_1
X_06029_ top.sram_interface.init_counter\[4\] _02928_ top.sram_interface.init_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05565__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__and2_1
X_10991_ clknet_leaf_62_clk _01556_ _00381_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08729__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05868__A1 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ clknet_leaf_22_clk _02162_ _01002_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06863__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11543_ clknet_leaf_72_clk _02108_ _00933_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06293__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11474_ clknet_leaf_98_clk _02039_ _00864_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[31\]
+ sky130_fd_sc_hd__dfstp_2
X_10425_ net766 net601 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08990__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__and2_1
X_10287_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__and2_1
XANTENNA__10414__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08742__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05400_ top.findLeastValue.least2\[4\] vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06380_ top.hist_data_o\[1\] top.hist_data_o\[0\] vssd1 vssd1 vccd1 vccd1 _03245_
+ sky130_fd_sc_hd__nand2_1
X_05331_ top.cb_syn.count\[5\] vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ _04207_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__nor2_1
X_07001_ _02512_ net126 net123 _03685_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08981__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__B2 top.findLeastValue.sum\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ top.WB.CPU_DAT_O\[16\] net1341 net318 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__mux2_1
X_07903_ net421 _04447_ _04448_ net263 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__o211a_1
X_08883_ net1106 top.WB.CPU_DAT_O\[19\] net302 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout195_A _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07834_ net431 net1537 net248 top.findLeastValue.sum\[31\] _04393_ vssd1 vssd1 vccd1
+ vccd1 _01820_ sky130_fd_sc_hd__a221o_1
XANTENNA__05547__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ top.hTree.tree_reg\[44\] top.findLeastValue.sum\[44\] net286 vssd1 vssd1
+ vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07696_ top.findLeastValue.least1\[2\] net264 _04280_ vssd1 vssd1 vccd1 vccd1 _04282_
+ sky130_fd_sc_hd__a21oi_1
X_09504_ net728 net563 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__and2_1
X_06716_ _02407_ top.findLeastValue.val2\[44\] top.findLeastValue.val2\[43\] _02408_
+ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a22o_1
X_06647_ _02437_ top.findLeastValue.val1\[9\] top.findLeastValue.val1\[8\] _02438_
+ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__o221a_1
X_09435_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout627_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06578_ top.cb_syn.num_lefts\[0\] top.cb_syn.num_lefts\[4\] top.cb_syn.num_lefts\[6\]
+ top.cb_syn.num_lefts\[2\] top.header_synthesis.count\[2\] top.header_synthesis.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09366_ net398 _04322_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nand2_1
X_08317_ top.cb_syn.char_path_n\[46\] net379 net338 top.cb_syn.char_path_n\[44\] net182
+ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05529_ net439 top.histogram.wr_r_en\[1\] net360 _02608_ _02613_ vssd1 vssd1 vccd1
+ vccd1 _02614_ sky130_fd_sc_hd__a311o_1
X_09297_ top.histogram.total\[4\] top.histogram.total\[5\] top.histogram.total\[6\]
+ top.histogram.total\[7\] net509 net506 vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__mux4_1
X_08248_ net1719 net205 _04686_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__o21a_1
X_08179_ top.cb_syn.char_path_n\[115\] net378 net334 top.cb_syn.char_path_n\[113\]
+ net181 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a221o_1
X_10210_ net824 net659 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ clknet_leaf_27_clk _01755_ _00580_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08972__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925__888 vssd1 vssd1 vccd1 vccd1 _11925__888/HI net888 sky130_fd_sc_hd__conb_1
X_10141_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05538__B1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10974_ clknet_leaf_50_clk _01539_ _00364_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11526_ clknet_leaf_80_clk _02091_ _00916_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11457_ clknet_leaf_85_clk _02022_ _00847_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output89_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ clknet_leaf_15_clk _01953_ _00778_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10408_ net741 net576 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__and2_1
XANTENNA__08963__A0 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__and2_1
X_05880_ net1686 top.WB.CPU_DAT_O\[18\] net350 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ _04146_ _04149_ _04110_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06501_ top.histogram.total\[16\] top.histogram.total\[15\] top.histogram.total\[14\]
+ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__and4_1
X_09220_ net491 net1704 _03371_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_start
+ sky130_fd_sc_hd__o21a_1
X_07481_ net1338 net344 _04045_ _04083_ _04085_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a221o_1
X_06432_ net1188 _03287_ net300 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06363_ top.hist_addr\[1\] top.hist_addr\[0\] vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__or2_1
X_09151_ _05144_ net456 net443 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ top.cb_syn.num_lefts\[4\] _04594_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__xnor2_1
X_09082_ net443 net450 _05107_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05314_ top.compVal\[20\] vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__inv_2
X_08033_ net514 top.cb_syn.curr_state\[0\] _04181_ vssd1 vssd1 vccd1 vccd1 _04545_
+ sky130_fd_sc_hd__or3_1
X_06294_ net484 _03089_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold800 top.cb_syn.char_path_n\[17\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout208_A _02620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold811 top.compVal\[31\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 top.cb_syn.char_path_n\[69\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold855 top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 top.compVal\[22\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 top.hTree.node_reg\[29\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05768__B1 _02806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout577_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ top.sram_interface.TRN_counter\[2\] top.sram_interface.TRN_counter\[0\] _02914_
+ top.sram_interface.TRN_counter\[1\] vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__or4b_2
X_08866_ net509 _05039_ _05046_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a21bo_1
X_08797_ top.path\[70\] top.path\[71\] net510 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__mux2_1
X_07817_ net476 _04378_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__or2_1
X_07748_ net257 _04323_ _04324_ net997 net433 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout744_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05940__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07679_ net472 _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__nand2_1
X_09418_ net962 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__clkbuf_1
X_10690_ clknet_leaf_107_clk _01321_ _00080_ vssd1 vssd1 vccd1 vccd1 top.path\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_09349_ net1016 net225 net215 _04379_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06991__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06248__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ clknet_leaf_14_clk _01876_ _00701_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11242_ clknet_leaf_69_clk net1571 _00632_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11173_ clknet_leaf_51_clk _01738_ _00563_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[119\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_95_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07748__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ net819 net654 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__and2_1
XANTENNA_input40_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10055_ net719 net554 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__and2_1
XANTENNA__09370__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A1 top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05931__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ clknet_leaf_65_clk _01522_ _00347_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ clknet_leaf_28_clk top.header_synthesis.next_write_zeroes _00278_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.write_zeroes sky130_fd_sc_hd__dfrtp_1
XANTENNA__08228__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07531__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold107 top.histogram.sram_out\[16\] vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
X_11509_ clknet_leaf_119_clk _02074_ _00899_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05998__A0 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 top.cb_syn.char_path\[15\] vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 top.path\[18\] vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09284__S0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 net611 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06981_ net486 _03088_ net484 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06962__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05932_ top.compVal\[29\] net158 net145 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 _02246_ sky130_fd_sc_hd__a22o_1
X_08720_ net542 _02591_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__nor2_1
X_08651_ _04791_ _04868_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__or2_1
X_05863_ net542 net456 _02799_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__and3_1
X_07602_ _02543_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__nor2_1
X_08582_ _02542_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05794_ net1428 _02817_ _02819_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__o21a_1
X_07533_ _04131_ _04132_ net289 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__mux2_1
XANTENNA__07675__B1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07464_ _04051_ _04053_ net393 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06415_ top.hist_data_o\[27\] _03262_ top.hist_data_o\[28\] vssd1 vssd1 vccd1 vccd1
+ _03277_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05431__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09203_ net1679 _05183_ net1592 top.controller.fin_reg\[7\] vssd1 vssd1 vccd1 vccd1
+ _05184_ sky130_fd_sc_hd__or4b_1
X_09134_ _05139_ _05140_ _05141_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__or3_1
X_07395_ _03834_ net271 _04027_ net277 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1
+ vccd1 _01889_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout325_A _04917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06346_ top.hist_addr\[2\] _03097_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06277_ top.hist_addr\[4\] _03098_ top.hist_addr\[5\] vssd1 vssd1 vccd1 vccd1 _03148_
+ sky130_fd_sc_hd__a21oi_1
X_09065_ net444 net455 _03013_ _05093_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a211o_1
XANTENNA__05989__A0 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold630 top.sram_interface.word_cnt\[6\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
X_08016_ net406 _02790_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor2_1
Xhold663 top.sram_interface.init_counter\[2\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 top.controller.fin_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 top.hTree.tree_reg\[7\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 top.cb_syn.end_check vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 top.hist_data_o\[21\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 top.compVal\[42\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ net773 net608 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__and2_1
XANTENNA__09573__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ top.cb_syn.max_index\[5\] _05060_ top.cb_syn.max_index\[6\] vssd1 vssd1 vccd1
+ vccd1 _05064_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06953__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net854 net689 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09352__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ _02808_ _05035_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__nand2_1
X_11860_ clknet_leaf_114_clk _02393_ _01232_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_10811_ clknet_leaf_32_clk _00009_ _00201_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11791_ clknet_leaf_92_clk _02325_ _01163_ vssd1 vssd1 vccd1 vccd1 top.compVal\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10742_ clknet_leaf_6_clk _00032_ _00132_ vssd1 vssd1 vccd1 vccd1 top.histogram.eof_n
+ sky130_fd_sc_hd__dfrtp_4
X_10673_ clknet_leaf_106_clk _01304_ _00063_ vssd1 vssd1 vccd1 vccd1 top.path\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06871__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07513__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07969__B2 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940__903 vssd1 vssd1 vccd1 vccd1 _11940__903/HI net903 sky130_fd_sc_hd__conb_1
XANTENNA__06172__A top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ clknet_leaf_85_clk _01790_ _00615_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08394__A1 top.cb_syn.char_path_n\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07197__A2 _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ clknet_leaf_64_clk _01721_ _00546_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11087_ clknet_leaf_46_clk _01652_ _00477_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[33\]
+ sky130_fd_sc_hd__dfrtp_4
X_10107_ net812 net647 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__and2_1
X_10038_ net837 net672 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__and2_1
XANTENNA__09343__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06200_ top.cw1\[7\] _03073_ _02602_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a21o_1
X_07180_ _03797_ _03802_ _03800_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06131_ net1466 net164 net157 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a21o_1
X_06062_ _02526_ top.cb_syn.zero_count\[7\] vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_57_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07188__A2 _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__and2_1
Xfanout428 _02549_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_2
Xfanout417 net422 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_4
Xfanout406 _02786_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_4
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
X_09752_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__and2_1
XANTENNA__06935__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ top.header_synthesis.count\[0\] _02566_ _03370_ _04897_ vssd1 vssd1 vccd1
+ vccd1 _04904_ sky130_fd_sc_hd__and4_1
XANTENNA__05426__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09334__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06964_ net456 net288 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nor2_1
X_05915_ _02887_ _02896_ _02581_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__o21ai_1
X_09683_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout275_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06895_ top.compVal\[6\] top.findLeastValue.val1\[6\] net153 vssd1 vssd1 vccd1 vccd1
+ _03653_ sky130_fd_sc_hd__mux2_1
X_08634_ _02542_ _04851_ _04853_ _02541_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_68_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05846_ top.sram_interface.counter_HTREE\[2\] _02854_ vssd1 vssd1 vccd1 vccd1 _02868_
+ sky130_fd_sc_hd__nand2_1
X_08565_ _02543_ top.cb_syn.h_element\[63\] _04562_ vssd1 vssd1 vccd1 vccd1 _04786_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05777_ net423 net36 vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__and2_1
XANTENNA__07360__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ top.cb_syn.char_path_n\[102\] top.cb_syn.char_path_n\[101\] top.cb_syn.char_path_n\[104\]
+ top.cb_syn.char_path_n\[103\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_81_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08496_ net1100 top.cb_syn.char_path_n\[63\] net230 vssd1 vssd1 vccd1 vccd1 _01546_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ _04053_ _04054_ _04049_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07378_ _03850_ net273 _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__and3b_1
X_06329_ top.cb_syn.curr_index\[3\] _02584_ _02607_ _02537_ _03197_ vssd1 vssd1 vccd1
+ vccd1 _03198_ sky130_fd_sc_hd__a221o_1
X_09117_ _03368_ _05124_ top.histogram.eof_n top.dut.out_valid vssd1 vssd1 vccd1 vccd1
+ _05131_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_79_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ top.WB.CPU_DAT_O\[2\] net1373 net316 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 net74 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 top.histogram.total\[5\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ clknet_leaf_35_clk _01575_ _00400_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[92\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold482 top.hTree.tree_reg\[12\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _01806_ vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06926__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900__931 vssd1 vssd1 vccd1 vccd1 net931 _11900__931/LO sky130_fd_sc_hd__conb_1
XANTENNA__06139__B1 _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11912_ net943 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_11843_ clknet_leaf_96_clk _02376_ _01215_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_11774_ clknet_leaf_41_clk _02313_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_10725_ clknet_leaf_25_clk _01356_ _00115_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10656_ clknet_leaf_82_clk _01287_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10417__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ net797 net632 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__and2_1
XANTENNA__07811__A0 top.findLeastValue.sum\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ clknet_leaf_25_clk _01773_ _00598_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.setup
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06917__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ clknet_leaf_53_clk _01704_ _00529_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09316__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05700_ top.hTree.node_reg\[37\] net307 _02755_ _02756_ vssd1 vssd1 vccd1 vccd1 _02757_
+ sky130_fd_sc_hd__a211o_1
X_06680_ top.compVal\[33\] _02488_ _02489_ top.compVal\[32\] vssd1 vssd1 vccd1 vccd1
+ _03478_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05631_ _02697_ _02698_ net468 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_47_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ net1754 net194 _04737_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__o21a_1
X_05562_ net93 net171 _02641_ net213 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a22o_1
XANTENNA__08991__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07301_ _03740_ _03961_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ top.cb_syn.char_path_n\[64\] net371 net328 top.cb_syn.char_path_n\[62\] net175
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05493_ net439 net526 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__and2_1
XANTENNA__08842__A2 top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07232_ top.findLeastValue.val2\[42\] top.findLeastValue.val1\[42\] vssd1 vssd1 vccd1
+ vccd1 _03908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07163_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__inv_2
X_06114_ _02450_ _02999_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ top.findLeastValue.val2\[17\] top.findLeastValue.val1\[17\] vssd1 vssd1 vccd1
+ vccd1 _03770_ sky130_fd_sc_hd__or2_1
X_06045_ _02449_ top.cb_syn.zeroes\[4\] top.cb_syn.zeroes\[3\] _02450_ vssd1 vssd1
+ vccd1 vccd1 _02945_ sky130_fd_sc_hd__a22o_1
Xfanout203 net205 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
Xfanout214 net219 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net247 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_4
X_09804_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__and2_1
Xfanout225 net227 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
XFILLER_0_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06908__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07996_ net1004 net254 _04521_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a21oi_1
X_09735_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06947_ top.findLeastValue.val1\[10\] net136 net113 top.compVal\[10\] vssd1 vssd1
+ vccd1 vccd1 _01971_ sky130_fd_sc_hd__o22a_1
XANTENNA__09570__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ net788 net623 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__and2_1
XANTENNA__07869__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ _04835_ _04836_ _02542_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__mux2_1
X_06878_ top.findLeastValue.val2\[15\] net131 net122 _03644_ vssd1 vssd1 vccd1 vccd1
+ _02023_ sky130_fd_sc_hd__o22a_1
X_05829_ top.hTree.state\[7\] top.hTree.state\[8\] vssd1 vssd1 vccd1 vccd1 _02851_
+ sky130_fd_sc_hd__or2_2
X_09597_ net742 net577 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__and2_1
X_08548_ net1241 top.cb_syn.char_path_n\[11\] net244 vssd1 vssd1 vccd1 vccd1 _01494_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08479_ net1112 top.cb_syn.char_path_n\[80\] net243 vssd1 vssd1 vccd1 vccd1 _01563_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05647__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ net757 net592 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__and2_1
X_11490_ clknet_leaf_12_clk _02055_ _00880_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.startup
+ sky130_fd_sc_hd__dfstp_1
X_10441_ net819 net654 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__and2_1
XANTENNA__08597__B2 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ net760 net595 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__and2_1
Xhold290 top.cb_syn.char_path\[11\] vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout770 net771 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_2
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_2
Xfanout781 net795 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_103_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ clknet_leaf_65_clk _02359_ _01198_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08809__C1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11757_ clknet_leaf_105_clk net1543 _01147_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05638__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ clknet_leaf_47_clk _01339_ _00098_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_11688_ clknet_leaf_78_clk _02238_ _01078_ vssd1 vssd1 vccd1 vccd1 top.compVal\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08037__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10639_ clknet_leaf_74_clk _01270_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08588__B2 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07260__A1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07850_ top.hTree.tree_reg\[27\] top.findLeastValue.sum\[27\] net282 vssd1 vssd1
+ vccd1 vccd1 _04406_ sky130_fd_sc_hd__mux2_1
X_07781_ top.hTree.tree_reg\[41\] top.findLeastValue.sum\[41\] _04251_ vssd1 vssd1
+ vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
X_06801_ _03559_ _03586_ _03595_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a211o_1
X_09520_ net735 net570 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__and2_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_06732_ _02436_ top.findLeastValue.val2\[10\] _03529_ vssd1 vssd1 vccd1 vccd1 _03530_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09451_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__and2_1
X_06663_ _02427_ top.findLeastValue.val1\[25\] top.findLeastValue.val1\[24\] _02428_
+ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__o22a_1
X_08402_ top.cb_syn.char_path_n\[3\] net197 _04763_ vssd1 vssd1 vccd1 vccd1 _01622_
+ sky130_fd_sc_hd__o21a_1
X_05614_ top.histogram.sram_out\[19\] net359 net410 top.hTree.node_reg\[19\] vssd1
+ vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
X_09382_ net960 _05268_ net228 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
X_06594_ _02865_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05545_ top.cb_syn.char_path\[30\] net546 net538 top.cb_syn.char_path\[94\] vssd1
+ vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
X_08333_ top.cb_syn.char_path_n\[38\] net379 net336 top.cb_syn.char_path_n\[36\] net182
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05629__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08264_ top.cb_syn.char_path_n\[72\] net201 _04694_ vssd1 vssd1 vccd1 vccd1 _01691_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout238_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout140_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05476_ net3 net415 net364 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 _02382_
+ sky130_fd_sc_hd__a22o_1
X_08195_ top.cb_syn.char_path_n\[107\] net383 net339 top.cb_syn.char_path_n\[105\]
+ net186 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout405_A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07215_ _03883_ _03886_ _03884_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07146_ top.findLeastValue.val2\[4\] top.findLeastValue.val1\[4\] vssd1 vssd1 vccd1
+ vccd1 _03822_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07077_ _03751_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06028_ _02930_ _02935_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09718_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__and2_1
X_07979_ net436 net1474 net250 top.findLeastValue.sum\[2\] _04509_ vssd1 vssd1 vccd1
+ vccd1 _01791_ sky130_fd_sc_hd__a221o_1
X_10990_ clknet_leaf_65_clk _01555_ _00380_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_09649_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ clknet_leaf_22_clk _02161_ _01001_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08806__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_116_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11542_ clknet_leaf_71_clk _02107_ _00932_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ clknet_leaf_99_clk _02038_ _00863_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[30\]
+ sky130_fd_sc_hd__dfstp_2
X_10424_ net763 net598 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10355_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__and2_1
X_10286_ net828 net663 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_29_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05556__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ clknet_leaf_83_clk _02342_ _01181_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05330_ net981 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_107_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_60_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ top.cw1\[0\] net148 _03662_ top.findLeastValue.histo_index\[0\] vssd1 vssd1
+ vccd1 vccd1 _03685_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07885__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08570__A top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06992__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08951_ top.WB.CPU_DAT_O\[17\] net1065 net318 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__mux2_1
X_07902_ net478 _04446_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__or2_1
X_08882_ net1207 top.WB.CPU_DAT_O\[20\] net302 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08733__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ net417 _04391_ _04392_ net255 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout188_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07764_ net438 net1582 net252 top.findLeastValue.sum\[45\] _04336_ vssd1 vssd1 vccd1
+ vccd1 _01834_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_27_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07695_ top.hTree.tree_reg\[57\] top.findLeastValue.least1\[2\] net280 vssd1 vssd1
+ vccd1 vccd1 _04281_ sky130_fd_sc_hd__mux2_1
X_09503_ net730 net565 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__and2_1
X_06715_ _02456_ top.compVal\[42\] _02408_ top.findLeastValue.val2\[43\] vssd1 vssd1
+ vccd1 vccd1 _03513_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08592__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06646_ _03439_ _03441_ _03443_ top.findLeastValue.val1\[8\] _02438_ vssd1 vssd1
+ vccd1 vccd1 _03444_ sky130_fd_sc_hd__a32o_1
X_09434_ net746 net581 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__and2_1
XANTENNA__08745__A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ net296 top.header_synthesis.header\[8\] vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__and2b_1
X_09365_ net1665 net221 _05256_ _05257_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
X_08316_ top.cb_syn.char_path_n\[46\] net202 _04720_ vssd1 vssd1 vccd1 vccd1 _01665_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_30 top.cb_syn.end_cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05528_ net356 net411 _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__or3_1
X_09296_ net425 _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__or2_1
X_08247_ top.cb_syn.char_path_n\[81\] net385 net340 top.cb_syn.char_path_n\[79\] net188
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05459_ net21 net414 net363 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 _02399_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08178_ top.cb_syn.char_path_n\[115\] net198 _04651_ vssd1 vssd1 vccd1 vccd1 _01734_
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_65_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07129_ top.findLeastValue.val2\[10\] top.findLeastValue.val1\[10\] vssd1 vssd1 vccd1
+ vccd1 _03805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10071_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05538__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ clknet_leaf_49_clk _01538_ _00363_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_74_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08583__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ clknet_leaf_80_clk _02090_ _00915_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11456_ clknet_leaf_86_clk _02021_ _00846_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10425__A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ clknet_leaf_15_clk _01952_ _00777_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10407_ net746 net581 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__and2_1
X_10338_ net730 net565 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10269_ net723 net558 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05529__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08574__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06500_ top.histogram.total\[13\] top.histogram.total\[12\] _03332_ vssd1 vssd1 vccd1
+ vccd1 _03333_ sky130_fd_sc_hd__and3_1
X_07480_ top.dut.bits_in_buf_next\[1\] _04071_ _04084_ _04060_ vssd1 vssd1 vccd1 vccd1
+ _04085_ sky130_fd_sc_hd__o211a_1
X_06431_ top.hist_data_o\[22\] _03273_ _03259_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06362_ top.sram_interface.init_counter\[1\] top.sram_interface.init_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__xor2_1
X_09150_ net455 top.sram_interface.word_cnt\[13\] _05100_ net1047 vssd1 vssd1 vccd1
+ vccd1 _00047_ sky130_fd_sc_hd__a22o_1
X_08101_ _04590_ _04596_ _04600_ _04589_ net1661 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a32o_1
X_06293_ net1075 net165 _03163_ net208 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a22o_1
X_09081_ net443 net459 _05096_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05313_ top.compVal\[22\] vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__inv_2
X_08032_ _02525_ _04544_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold801 top.cb_syn.char_path_n\[82\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 top.cb_syn.char_path_n\[70\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 top.cb_syn.char_path_n\[124\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 net96 vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 top.hist_data_o\[27\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold856 top.findLeastValue.sum\[22\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05429__A top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ net832 net667 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__and2_1
X_08934_ top.cb_syn.max_index\[1\] _05059_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__xnor2_1
XANTENNA__05768__B2 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08865_ _05047_ _05037_ net506 _05046_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a2bb2o_1
X_08796_ net426 _04983_ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__o21a_1
X_07816_ top.findLeastValue.sum\[34\] _04378_ net391 vssd1 vssd1 vccd1 vccd1 _04379_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07747_ net472 _04320_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__or2_1
XANTENNA__05940__B2 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07678_ top.findLeastValue.least1\[5\] net264 _04265_ vssd1 vssd1 vccd1 vccd1 _04267_
+ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ net972 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07693__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06629_ _02429_ top.findLeastValue.val1\[23\] top.findLeastValue.val1\[22\] _02430_
+ _03425_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ net1001 net225 net215 _04383_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06248__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ clknet_leaf_43_clk _01875_ _00700_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ net344 _04050_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[10\] sky130_fd_sc_hd__and2_1
X_11241_ clknet_leaf_69_clk net1444 _00631_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ clknet_leaf_49_clk _01737_ _00562_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10123_ net833 net668 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__and2_1
XANTENNA__06869__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__and2_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05931__B2 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ clknet_leaf_64_clk _01521_ _00346_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ clknet_leaf_26_clk top.header_synthesis.next_start _00277_ vssd1 vssd1 vccd1
+ vccd1 top.header_synthesis.start sky130_fd_sc_hd__dfrtp_1
XANTENNA__05521__B _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07531__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ clknet_leaf_119_clk _02073_ _00898_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold108 top.path\[42\] vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 top.cb_syn.curr_index\[2\] vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ clknet_leaf_91_clk _02004_ _00829_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[43\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09284__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06947__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06980_ net1694 _03670_ _03677_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05931_ top.compVal\[30\] net158 net145 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 _02247_ sky130_fd_sc_hd__a22o_1
X_08650_ net520 _04866_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__or2_2
X_05862_ _02553_ _02562_ _02801_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__or3_1
X_07601_ top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\] _04199_ vssd1 vssd1 vccd1
+ vccd1 _04201_ sky130_fd_sc_hd__or3_2
XANTENNA__07372__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ top.cb_syn.char_path_n\[73\] top.cb_syn.char_path_n\[74\] top.cb_syn.char_path_n\[77\]
+ top.cb_syn.char_path_n\[78\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_37_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05793_ net1489 _02818_ _02820_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__o21ba_1
X_07532_ top.cb_syn.char_path_n\[66\] top.cb_syn.char_path_n\[65\] top.cb_syn.char_path_n\[68\]
+ top.cb_syn.char_path_n\[67\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__mux4_1
XANTENNA__07675__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07463_ _04058_ _04067_ _04069_ _04048_ _04068_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a221o_1
XANTENNA__05686__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06414_ net1461 net301 _03276_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _05181_ _05183_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_1
X_09133_ net455 top.sram_interface.word_cnt\[7\] _02798_ _05096_ net542 vssd1 vssd1
+ vccd1 vccd1 _05141_ sky130_fd_sc_hd__a32o_1
X_07394_ _03825_ _03832_ _03830_ _03827_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06345_ _02926_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout220_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06276_ net484 net361 _03144_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a211o_1
X_09064_ net447 net458 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold620 _01807_ vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
X_08015_ top.findLeastValue.alternator_timer\[2\] top.findLeastValue.alternator_timer\[1\]
+ top.findLeastValue.alternator_timer\[0\] _03666_ top.findLeastValue.alternator_timer\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__a41o_1
XFILLER_0_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold631 top.hTree.tree_reg\[45\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 top.histogram.total\[9\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 top.hTree.state\[1\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold675 top.sram_interface.init_counter\[4\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 top.findLeastValue.sum\[26\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 top.hTree.state\[2\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__and2_1
XANTENNA__09573__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__and2_1
X_08917_ _05063_ top.cb_syn.max_index\[7\] _05059_ vssd1 vssd1 vccd1 vccd1 _01407_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08155__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
X_08848_ net452 _02807_ _05035_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__and3_1
XANTENNA__07363__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _02547_ _04922_ _04967_ top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1
+ _04968_ sky130_fd_sc_hd__o211a_1
X_10810_ clknet_leaf_39_clk _00008_ _00200_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11790_ clknet_leaf_95_clk _02324_ _01162_ vssd1 vssd1 vccd1 vccd1 top.compVal\[39\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10741_ clknet_leaf_6_clk _00031_ _00131_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10672_ clknet_leaf_106_clk _01303_ _00062_ vssd1 vssd1 vccd1 vccd1 top.path\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09748__B net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07513__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ clknet_leaf_83_clk _01789_ _00614_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09040__A0 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ clknet_leaf_64_clk _01720_ _00545_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05601__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ clknet_leaf_42_clk _01651_ _00476_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[32\]
+ sky130_fd_sc_hd__dfrtp_2
X_10106_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__and2_1
X_10037_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_87_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_106_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10939_ clknet_leaf_53_clk _01504_ _00329_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07657__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05668__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06880__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06130_ net458 net361 net208 net407 vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__and4_2
X_06061_ _02959_ _02960_ _02958_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_117_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08989__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__and2_1
Xfanout407 _02786_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_2
Xfanout429 _02548_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_4
Xfanout418 net422 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_4
X_09751_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__and2_1
X_06963_ net1476 _02576_ _03395_ net287 net955 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a32o_1
XANTENNA__08790__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05914_ net489 net524 _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__and3b_1
X_08702_ top.header_synthesis.count\[6\] _04902_ _04895_ vssd1 vssd1 vccd1 vccd1 _04903_
+ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_78_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_09682_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__and2_1
X_06894_ top.findLeastValue.val2\[7\] net129 net120 _03652_ vssd1 vssd1 vccd1 vccd1
+ _02015_ sky130_fd_sc_hd__o22a_1
X_08633_ net497 _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__and2_1
XANTENNA__07922__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05845_ _02858_ _02860_ _02863_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout170_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _04785_ net491 _04783_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__mux2_1
X_05776_ top.compVal\[32\] net162 net147 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ _02317_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout268_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07515_ _04113_ _04114_ net290 vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08495_ net1225 top.cb_syn.char_path_n\[64\] net230 vssd1 vssd1 vccd1 vccd1 _01547_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08845__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06320__A1 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07446_ top.dut.bit_buf\[7\] top.dut.bit_buf\[0\] net713 vssd1 vssd1 vccd1 vccd1
+ _04054_ sky130_fd_sc_hd__mux2_1
X_07377_ _03848_ _03849_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06328_ _03193_ _03195_ _03196_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__or3_1
X_09116_ net353 _05123_ _05130_ net1658 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a22o_1
XANTENNA__07820__A1 top.findLeastValue.sum\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ top.WB.CPU_DAT_O\[3\] net1418 net316 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06259_ top.TRN_char_index\[4\] _03055_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold472 top.cb_syn.char_path\[66\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 top.path\[64\] vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold461 top.path\[35\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09022__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold494 top.hTree.nulls\[50\] vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 net63 vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
X_09949_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_69_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
X_11911_ net942 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_11842_ clknet_leaf_112_clk _02375_ _01214_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07639__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ clknet_leaf_42_clk _02312_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07639__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10724_ clknet_leaf_17_clk _01355_ _00114_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10655_ clknet_leaf_81_clk _01286_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10586_ net797 net632 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ clknet_leaf_26_clk _01772_ _00597_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.wait_cycle
+ sky130_fd_sc_hd__dfstp_1
X_11138_ clknet_leaf_54_clk _01703_ _00528_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[84\]
+ sky130_fd_sc_hd__dfrtp_2
X_11069_ clknet_leaf_58_clk _01634_ _00459_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09941__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07878__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05630_ top.cb_syn.char_path\[48\] net531 net310 top.cb_syn.char_path\[112\] vssd1
+ vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05561_ net1799 net354 _02639_ _02640_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08827__B1 top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07300_ _03740_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__or2_1
X_08280_ top.cb_syn.char_path_n\[64\] net193 _04702_ vssd1 vssd1 vccd1 vccd1 _01683_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05492_ _02563_ _02576_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ _03904_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07162_ _03823_ _03836_ _03820_ _03822_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o211a_1
X_06113_ _02997_ _03002_ _03009_ _02996_ net1662 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07093_ top.findLeastValue.val2\[19\] top.findLeastValue.val1\[19\] vssd1 vssd1 vccd1
+ vccd1 _03769_ sky130_fd_sc_hd__xor2_1
XANTENNA__09004__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06044_ _02447_ _02944_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__nand2_1
XANTENNA__08358__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout204 net205 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlymetal6s2s_1
X_09803_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__and2_1
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06369__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout215 net219 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
XANTENNA__08763__C1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout259 _04256_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
Xfanout248 net253 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09307__A1 top.header_synthesis.bit1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ top.hTree.state\[1\] net254 net953 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a21oi_1
X_09734_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__and2_1
XANTENNA__05871__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ top.findLeastValue.val1\[11\] net135 net113 net1731 vssd1 vssd1 vccd1 vccd1
+ _01972_ sky130_fd_sc_hd__o22a_1
X_09665_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__and2_1
XANTENNA__07869__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ top.compVal\[15\] top.findLeastValue.val1\[15\] net152 vssd1 vssd1 vccd1
+ vccd1 _03644_ sky130_fd_sc_hd__mux2_1
X_08616_ top.cb_syn.char_path_n\[9\] top.cb_syn.char_path_n\[10\] top.cb_syn.char_path_n\[13\]
+ top.cb_syn.char_path_n\[14\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__mux4_1
X_05828_ top.hTree.state\[7\] top.hTree.state\[8\] vssd1 vssd1 vccd1 vccd1 _02850_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09596_ net742 net577 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__and2_1
X_08547_ net1287 top.cb_syn.char_path_n\[12\] net245 vssd1 vssd1 vccd1 vccd1 _01495_
+ sky130_fd_sc_hd__mux2_1
X_05759_ net542 _02799_ _02802_ _02562_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a211o_1
X_08478_ net1245 top.cb_syn.char_path_n\[81\] net246 vssd1 vssd1 vccd1 vccd1 _01564_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06844__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07429_ top.dut.bits_in_buf\[1\] top.dut.bits_in_buf\[0\] top.dut.bits_in_buf\[2\]
+ net713 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__o31a_1
X_10440_ net827 net662 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__and2_1
X_10371_ net760 net595 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__and2_1
XANTENNA__08422__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07827__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 top.cb_syn.char_path\[84\] vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 top.cb_syn.char_path\[101\] vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold764_A top.findLeastValue.sum\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net762 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08658__A _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 net794 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_2
Xfanout771 net777 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_2
Xfanout782 net783 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06877__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ clknet_leaf_66_clk _02358_ _01197_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ clknet_leaf_105_clk _00026_ _01146_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10707_ clknet_leaf_47_clk _01338_ _00097_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ clknet_leaf_102_clk _02237_ _01077_ vssd1 vssd1 vccd1 vccd1 top.compVal\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_10638_ clknet_leaf_72_clk _01269_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09936__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ net860 net695 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__and2_1
X_11907__938 vssd1 vssd1 vccd1 vccd1 net938 _11907__938/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07548__A0 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ top.hTree.tree_reg\[41\] top.findLeastValue.sum\[41\] net285 vssd1 vssd1
+ vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
X_06800_ _03565_ _03574_ _03582_ _03593_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a221o_1
XANTENNA__08760__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ _02435_ top.findLeastValue.val2\[11\] _02474_ top.compVal\[10\] vssd1 vssd1
+ vccd1 vccd1 _03529_ sky130_fd_sc_hd__a2bb2o_1
X_09450_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__and2_1
X_08401_ top.cb_syn.char_path_n\[4\] net375 net332 top.cb_syn.char_path_n\[2\] net179
+ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06662_ top.compVal\[27\] _02490_ top.findLeastValue.val1\[26\] _02426_ vssd1 vssd1
+ vccd1 vccd1 _03460_ sky130_fd_sc_hd__a22o_1
X_05613_ _02682_ _02683_ net467 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__o21a_1
X_09381_ top.hTree.nulls\[53\] _04298_ net400 vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__mux2_1
X_06593_ net431 _02553_ _03390_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__or3b_1
X_08332_ top.cb_syn.char_path_n\[38\] net201 _04728_ vssd1 vssd1 vccd1 vccd1 _01657_
+ sky130_fd_sc_hd__o21a_1
X_05544_ net97 net167 _02626_ net213 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08263_ top.cb_syn.char_path_n\[73\] net380 net337 top.cb_syn.char_path_n\[71\] net184
+ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a221o_1
XANTENNA__07411__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06826__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout133_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05475_ net4 net414 net362 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 _02383_
+ sky130_fd_sc_hd__o22a_1
X_07214_ _03872_ _03873_ _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ top.cb_syn.char_path_n\[107\] net203 _04659_ vssd1 vssd1 vccd1 vccd1 _01726_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout300_A _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07076_ top.findLeastValue.val2\[26\] top.findLeastValue.val1\[26\] vssd1 vssd1 vccd1
+ vccd1 _03752_ sky130_fd_sc_hd__or2_1
X_06027_ net1748 _02929_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nor2_1
XANTENNA__08736__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ net419 _04507_ _04508_ net261 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__o211a_1
X_09717_ net863 net698 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__and2_1
X_06929_ top.findLeastValue.val1\[28\] net133 net114 net1734 vssd1 vssd1 vccd1 vccd1
+ _01989_ sky130_fd_sc_hd__o22a_1
X_09648_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06429__C net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ net798 net633 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__and2_1
X_11610_ clknet_leaf_22_clk _02160_ _01000_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11541_ clknet_leaf_69_clk _02106_ _00931_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ clknet_leaf_99_clk _02037_ _00862_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[29\]
+ sky130_fd_sc_hd__dfstp_1
X_10423_ net739 net574 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__and2_1
X_10354_ net719 net554 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__and2_1
XANTENNA__06461__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10285_ net828 net663 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__and2_1
XANTENNA__05556__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net592 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ clknet_leaf_83_clk _02341_ _01180_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11739_ clknet_leaf_107_clk _02289_ _01129_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09666__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07769__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05795__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ top.WB.CPU_DAT_O\[18\] net1165 net318 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__mux2_1
X_07901_ top.findLeastValue.sum\[17\] _04446_ net392 vssd1 vssd1 vccd1 vccd1 _04447_
+ sky130_fd_sc_hd__mux2_1
X_08881_ net1326 top.WB.CPU_DAT_O\[21\] net302 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07832_ net470 _04390_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__or2_1
XANTENNA__09143__C1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ net431 _04255_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nor2_1
X_09502_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__and2_1
X_07694_ top.hTree.tree_reg\[57\] _04248_ net388 vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__and3_1
X_06714_ _03510_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08592__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06645_ _02443_ top.findLeastValue.val1\[3\] _03435_ _03440_ _03442_ vssd1 vssd1
+ vccd1 vccd1 _03443_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout250_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ net746 net581 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_111_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09364_ top.hTree.nulls\[47\] net401 net229 vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout348_A _02915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ top.cb_syn.char_path_n\[47\] net382 net338 top.cb_syn.char_path_n\[45\] net185
+ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06576_ _03372_ _03375_ _03370_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _02735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05527_ top.sram_interface.check _02610_ top.sram_interface.word_cnt\[13\] net446
+ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_20 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ top.histogram.total\[2\] top.histogram.total\[3\] net509 vssd1 vssd1 vccd1
+ vccd1 _05239_ sky130_fd_sc_hd__mux2_1
X_08246_ net1736 net199 _04685_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__o21a_1
X_05458_ net22 net413 net362 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 _02400_
+ sky130_fd_sc_hd__o22a_1
X_08177_ top.cb_syn.char_path_n\[116\] net377 net334 top.cb_syn.char_path_n\[114\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a221o_1
XANTENNA__05483__B2 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05389_ top.cw2\[6\] vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07128_ _02474_ _02496_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__nor2_1
X_07059_ top.findLeastValue.val2\[39\] top.findLeastValue.val1\[39\] _03734_ vssd1
+ vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10070_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09592__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10972_ clknet_leaf_48_clk _01537_ _00362_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08936__A _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08660__A1 top.cb_syn.char_path_n\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11524_ clknet_leaf_120_clk _02089_ _00914_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07986__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05474__B2 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ clknet_leaf_86_clk _02020_ _00845_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ net746 net581 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11386_ clknet_leaf_15_clk _01951_ _00776_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_111_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10337_ net728 net563 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__and2_1
X_10268_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__and2_1
X_10199_ net819 net654 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08574__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06430_ net1045 net299 _03286_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05701__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06361_ _03225_ _03227_ net459 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o21a_1
X_08100_ top.cb_syn.num_lefts\[4\] top.cb_syn.num_lefts\[3\] _04592_ top.cb_syn.num_lefts\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06292_ net454 _03149_ _03151_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a31o_1
XANTENNA__07896__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ net533 _05106_ _05105_ _05103_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_32_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05312_ top.compVal\[23\] vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__inv_2
X_08031_ top.CB_read_complete top.cb_syn.setup _04542_ vssd1 vssd1 vccd1 vccd1 _04544_
+ sky130_fd_sc_hd__and3_1
XANTENNA__05465__B2 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput40 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
Xhold802 top.compVal\[44\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08403__B2 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold846 top.hist_addr\[1\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 top.compVal\[39\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold835 top.histogram.state\[5\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 top.cb_syn.char_path_n\[89\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08933_ top.cb_syn.max_index\[2\] _05059_ _05072_ _05074_ vssd1 vssd1 vccd1 vccd1
+ _01402_ sky130_fd_sc_hd__a22o_1
XANTENNA__08167__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout298_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _02550_ net402 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__and2_1
X_08795_ top.path\[76\] net404 net324 top.path\[77\] net503 vssd1 vssd1 vccd1 vccd1
+ _04984_ sky130_fd_sc_hd__o221a_1
X_07815_ top.hTree.tree_reg\[34\] top.findLeastValue.sum\[34\] net283 vssd1 vssd1
+ vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07746_ net472 _04322_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05940__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ net970 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07677_ top.hTree.tree_reg\[60\] top.findLeastValue.least1\[5\] net280 vssd1 vssd1
+ vccd1 vccd1 _04266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08890__A1 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06628_ _02429_ top.findLeastValue.val1\[23\] top.findLeastValue.val1\[22\] _02430_
+ _03424_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__o221ai_1
X_09347_ net973 net225 net215 _04387_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__a22o_1
X_06559_ net1602 _03325_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ net343 _04051_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[9\] sky130_fd_sc_hd__and2_1
X_11931__894 vssd1 vssd1 vccd1 vccd1 _11931__894/HI net894 sky130_fd_sc_hd__conb_1
X_08229_ top.cb_syn.char_path_n\[90\] net373 net331 top.cb_syn.char_path_n\[88\] net176
+ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05456__B2 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ clknet_leaf_69_clk net1568 _00630_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11171_ clknet_leaf_49_clk _01736_ _00561_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[117\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_95_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10122_ net817 net652 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__and2_1
XANTENNA__08430__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ net759 net594 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__and2_1
XANTENNA_hold844_A top.hTree.node_reg\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06885__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05931__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ clknet_leaf_64_clk _01520_ _00345_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_10886_ clknet_leaf_23_clk top.header_synthesis.next_header\[8\] _00276_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07684__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08881__A1 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06892__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ clknet_leaf_119_clk _02072_ _00897_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11438_ clknet_leaf_95_clk _02003_ _00828_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[42\]
+ sky130_fd_sc_hd__dfstp_1
Xhold109 top.path\[26\] vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
X_11369_ clknet_leaf_41_clk _01934_ _00759_ vssd1 vssd1 vccd1 vccd1 top.cw1\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06947__B2 top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05930_ top.compVal\[31\] net159 net144 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 _02248_ sky130_fd_sc_hd__a22o_1
X_05861_ _02417_ _02447_ _02878_ net481 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__o31a_1
X_07600_ top.cb_syn.cb_length\[2\] top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__or3_1
X_08580_ top.cb_syn.end_cnt\[3\] _04795_ _04797_ _04799_ top.cb_syn.end_cnt\[4\] vssd1
+ vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__o221a_1
X_07531_ top.cb_syn.char_path_n\[70\] top.cb_syn.char_path_n\[69\] top.cb_syn.char_path_n\[72\]
+ top.cb_syn.char_path_n\[71\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__mux4_1
X_05792_ _02820_ net1390 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_37_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06332__C1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07462_ _04050_ _04063_ top.dut.bits_in_buf_next\[0\] vssd1 vssd1 vccd1 vccd1 _04069_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08872__A1 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06413_ _03264_ _03275_ net301 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o21ai_1
X_07393_ _03837_ net271 _04026_ net277 top.findLeastValue.sum\[3\] vssd1 vssd1 vccd1
+ vccd1 _01890_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_17_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09201_ top.controller.fin_reg\[1\] top.controller.fin_reg\[2\] net1681 top.controller.fin_reg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or4_1
X_06344_ top.sram_interface.init_counter\[1\] top.sram_interface.init_counter\[0\]
+ top.sram_interface.init_counter\[2\] vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09132_ _02906_ _02795_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__and2b_1
X_06275_ _03080_ _03145_ _02600_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__and3b_1
X_09063_ net447 net455 vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__nor2_1
Xhold610 top.cb_syn.zero_count\[3\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold621 top.cb_syn.pulse_first vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
X_08014_ top.findLeastValue.alternator_timer\[1\] top.findLeastValue.alternator_timer\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__nand2_1
XANTENNA__09854__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 top.cb_syn.zero_count\[2\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold643 top.hTree.tree_reg\[37\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 top.histogram.total\[6\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05874__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top.findLeastValue.sum\[24\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 _00020_ vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 top.cb_syn.i\[6\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net773 net608 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__and2_1
X_09896_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08916_ _04186_ _05062_ _04255_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__mux2_1
X_08847_ net513 top.translation.totalEn _05024_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__or3_1
XANTENNA__09352__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06166__A2 top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__B2 net1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08778_ _04924_ _04925_ _04926_ net505 net503 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__a221o_1
X_07729_ net472 _04305_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__or2_1
X_10740_ clknet_leaf_4_clk _00030_ _00130_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06874__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ clknet_leaf_106_clk _01302_ _00061_ vssd1 vssd1 vccd1 vccd1 top.path\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07823__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11223_ clknet_leaf_12_clk _01788_ _00613_ vssd1 vssd1 vccd1 vccd1 top.WorR sky130_fd_sc_hd__dfrtp_4
X_11154_ clknet_leaf_63_clk _01719_ _00544_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[100\]
+ sky130_fd_sc_hd__dfrtp_2
X_11085_ clknet_leaf_37_clk _01650_ _00475_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_10105_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__and2_1
XANTENNA__09780__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_106_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10938_ clknet_leaf_55_clk _01503_ _00328_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07657__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ clknet_leaf_27_clk _01454_ _00259_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06060_ top.cb_syn.zeroes\[2\] _02558_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09955__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout419 net422 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_2
Xfanout408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_2
X_09750_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__and2_1
X_06962_ net1711 net133 _03664_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__o21a_1
XANTENNA__08790__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05913_ _02551_ _02894_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__nor2_1
X_08701_ top.header_synthesis.count\[5\] _04896_ _04897_ vssd1 vssd1 vccd1 vccd1 _04902_
+ sky130_fd_sc_hd__and3_1
X_09681_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__and2_1
XANTENNA__09334__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ top.cb_syn.char_path_n\[43\] top.cb_syn.char_path_n\[44\] top.cb_syn.char_path_n\[47\]
+ top.cb_syn.char_path_n\[48\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__mux4_1
X_06893_ top.compVal\[7\] top.findLeastValue.val1\[7\] net153 vssd1 vssd1 vccd1 vccd1
+ _03652_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05844_ net448 net544 _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__and3_1
X_08563_ _04195_ _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09098__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05775_ top.compVal\[33\] net162 net147 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ _02318_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout163_A _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ top.cb_syn.char_path_n\[106\] top.cb_syn.char_path_n\[105\] top.cb_syn.char_path_n\[108\]
+ top.cb_syn.char_path_n\[107\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__mux4_1
X_08494_ net1385 top.cb_syn.char_path_n\[65\] net238 vssd1 vssd1 vccd1 vccd1 _01548_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ top.dut.bit_buf\[8\] top.dut.bit_buf\[1\] net714 vssd1 vssd1 vccd1 vccd1
+ _04053_ sky130_fd_sc_hd__mux2_1
XANTENNA__06856__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05869__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06320__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07376_ net273 _04014_ _04015_ net279 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1
+ vccd1 _01896_ sky130_fd_sc_hd__a32o_1
X_06327_ top.TRN_char_index\[1\] _02591_ _03191_ net446 vssd1 vssd1 vccd1 vccd1 _03196_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _05079_ _05124_ _05130_ net1446 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a22o_1
X_06258_ _03035_ _03129_ _02607_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__and3b_1
X_09046_ top.WB.CPU_DAT_O\[4\] net1369 net316 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout797_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold451 top.cb_syn.char_path\[43\] vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 top.cb_syn.char_path\[125\] vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ top.cb_syn.char_index\[6\] _03047_ _02605_ vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__a21oi_1
Xhold440 top.path\[49\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold473 _01549_ vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 top.path\[84\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 top.histogram.state\[2\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09948_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__and2_1
XANTENNA__05595__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06139__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__and2_1
X_11910_ net941 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_11841_ clknet_leaf_112_clk _02374_ _01213_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05898__A1 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ clknet_leaf_75_clk _02311_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10723_ clknet_leaf_17_clk _01354_ _00113_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08663__B _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10654_ clknet_leaf_81_clk _01285_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10585_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06614__D _03411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__C1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ clknet_leaf_26_clk _01771_ _00596_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11137_ clknet_leaf_54_clk _01702_ _00527_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[83\]
+ sky130_fd_sc_hd__dfrtp_2
X_11068_ clknet_leaf_59_clk _01633_ _00458_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__and2_1
XANTENNA__05889__A1 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05560_ top.histogram.sram_out\[28\] net360 net411 top.hTree.node_reg\[28\] vssd1
+ vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08827__A1 _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08854__A top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05491_ _02500_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__nor2_2
XANTENNA__06838__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07230_ top.findLeastValue.val2\[43\] top.findLeastValue.val1\[43\] vssd1 vssd1 vccd1
+ vccd1 _03906_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07161_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06112_ top.cb_syn.count\[4\] _03000_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or2_1
XANTENNA__06093__B net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07092_ top.findLeastValue.val2\[18\] top.findLeastValue.val1\[18\] vssd1 vssd1 vccd1
+ vccd1 _03768_ sky130_fd_sc_hd__xor2_2
X_06043_ _02876_ _02940_ _02941_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07409__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__and2_1
Xfanout238 net241 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout227 _05253_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
Xfanout216 net219 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05577__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout249 net253 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09307__A2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07994_ net448 net977 _04257_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__o21a_1
X_09733_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout280_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06945_ top.findLeastValue.val1\[12\] net136 net116 net1729 vssd1 vssd1 vccd1 vccd1
+ _01973_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout378_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__and2_1
X_06876_ top.findLeastValue.val2\[16\] net128 net121 _03643_ vssd1 vssd1 vccd1 vccd1
+ _02024_ sky130_fd_sc_hd__o22a_1
X_08615_ top.cb_syn.char_path_n\[11\] top.cb_syn.char_path_n\[12\] top.cb_syn.char_path_n\[15\]
+ top.cb_syn.char_path_n\[16\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05453__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09595_ net742 net577 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__and2_1
X_05827_ _02848_ top.sram_interface.counter_HTREE\[3\] top.sram_interface.counter_HTREE\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net1123 top.cb_syn.char_path_n\[13\] net245 vssd1 vssd1 vccd1 vccd1 _01496_
+ sky130_fd_sc_hd__mux2_1
X_05758_ net543 net457 _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__and3_1
X_08477_ net1264 top.cb_syn.char_path_n\[82\] net246 vssd1 vssd1 vccd1 vccd1 _01565_
+ sky130_fd_sc_hd__mux2_1
X_05689_ net1282 net170 _02747_ net209 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout712_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ top.findLeastValue.least1\[0\] net140 _03660_ top.findLeastValue.histo_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07359_ _03792_ _04000_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07254__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ net758 net593 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ top.WB.CPU_DAT_O\[21\] net1403 net313 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
Xhold270 top.cb_syn.char_path\[54\] vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 top.header_synthesis.header\[7\] vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 top.path\[62\] vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05568__B1 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout750 net753 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_2
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_2
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_2
Xfanout783 net786 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06178__B top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11824_ clknet_leaf_65_clk _02357_ _01196_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06893__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11755_ clknet_leaf_105_clk _00025_ _01145_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10706_ clknet_leaf_47_clk _01337_ _00096_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ clknet_leaf_100_clk _02236_ _01076_ vssd1 vssd1 vccd1 vccd1 top.compVal\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ clknet_leaf_77_clk _01268_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10568_ net861 net696 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__and2_1
XANTENNA__08993__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07796__A1 top.findLeastValue.sum\[38\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08840__C net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ net755 net590 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07548__A1 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05559__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ _02435_ top.findLeastValue.val2\[11\] vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__nand2_1
X_06661_ _02423_ top.findLeastValue.val1\[29\] top.findLeastValue.val1\[28\] _02424_
+ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__a22o_1
X_05612_ top.cb_syn.char_path\[51\] net530 net311 top.cb_syn.char_path\[115\] vssd1
+ vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a22o_1
X_08400_ top.cb_syn.char_path_n\[4\] net196 _04762_ vssd1 vssd1 vccd1 vccd1 _01623_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09380_ net1022 net222 _05266_ _05267_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
X_06592_ net448 net544 _03390_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__and3_1
X_08331_ top.cb_syn.char_path_n\[39\] net380 net337 top.cb_syn.char_path_n\[37\] net183
+ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a221o_1
X_05543_ top.hTree.node_reg\[63\] net356 _02624_ _02625_ vssd1 vssd1 vccd1 vccd1 _02626_
+ sky130_fd_sc_hd__a211o_1
X_08262_ top.cb_syn.char_path_n\[73\] net201 _04693_ vssd1 vssd1 vccd1 vccd1 _01692_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05474_ net5 net413 net362 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 _02384_
+ sky130_fd_sc_hd__o22a_1
X_07213_ _03881_ _03882_ _03884_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or4_1
X_08193_ top.cb_syn.char_path_n\[108\] net383 net339 top.cb_syn.char_path_n\[106\]
+ net186 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ top.findLeastValue.val2\[4\] top.findLeastValue.val1\[4\] vssd1 vssd1 vccd1
+ vccd1 _03820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08984__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07075_ top.findLeastValue.val2\[26\] top.findLeastValue.val1\[26\] vssd1 vssd1 vccd1
+ vccd1 _03751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05448__A top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06026_ net1757 _02930_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__xor2_1
XANTENNA__08736__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__A top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ net477 _04506_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__or2_1
X_09716_ net862 net697 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__and2_1
XANTENNA__05970__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06928_ top.findLeastValue.val1\[29\] net133 net115 top.compVal\[29\] vssd1 vssd1
+ vccd1 vccd1 _01990_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09647_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07711__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ top.compVal\[24\] top.findLeastValue.val1\[24\] net156 vssd1 vssd1 vccd1
+ vccd1 _03635_ sky130_fd_sc_hd__mux2_1
XANTENNA__05722__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ net798 net633 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__and2_1
X_08529_ net1152 top.cb_syn.char_path_n\[30\] net234 vssd1 vssd1 vccd1 vccd1 _01513_
+ sky130_fd_sc_hd__mux2_1
X_11540_ clknet_leaf_70_clk _02105_ _00930_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07570__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ clknet_leaf_99_clk _02036_ _00861_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[28\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08019__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ net739 net574 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__and2_1
XANTENNA__08975__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06450__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10284_ net833 net668 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__and2_1
Xfanout591 net592 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_2
Xfanout580 net583 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ clknet_leaf_83_clk _02340_ _01179_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ clknet_leaf_106_clk _02288_ _01128_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09947__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ clknet_leaf_91_clk _02219_ _01059_ vssd1 vssd1 vccd1 vccd1 top.compVal\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07769__B2 top.findLeastValue.sum\[44\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__A0 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06992__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07900_ top.hTree.tree_reg\[17\] top.findLeastValue.sum\[17\] net286 vssd1 vssd1
+ vccd1 vccd1 _04446_ sky130_fd_sc_hd__mux2_1
X_08880_ net1046 top.WB.CPU_DAT_O\[22\] net303 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07831_ top.hTree.tree_reg\[31\] top.findLeastValue.sum\[31\] net265 vssd1 vssd1
+ vccd1 vccd1 _04391_ sky130_fd_sc_hd__mux2_1
XANTENNA__07941__A1 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07762_ net421 _04334_ _04335_ net263 vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o211a_1
X_09501_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__and2_1
XANTENNA__05952__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07693_ net258 _04278_ _04279_ net1092 net432 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a32o_1
X_06713_ top.compVal\[42\] _02456_ _02457_ top.compVal\[41\] vssd1 vssd1 vccd1 vccd1
+ _03511_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06644_ _03436_ _03437_ _03431_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__or3b_1
X_09432_ net746 net581 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__and2_1
X_06575_ top.header_synthesis.count\[3\] _03374_ _03373_ vssd1 vssd1 vccd1 vccd1 _03375_
+ sky130_fd_sc_hd__a21oi_2
X_09363_ net401 _04327_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout243_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ top.cb_syn.char_path_n\[47\] net202 _04719_ vssd1 vssd1 vccd1 vccd1 _01666_
+ sky130_fd_sc_hd__o21a_1
X_05526_ net448 net536 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__and2_1
XANTENNA__07552__S0 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _04150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 top.cb_syn.end_cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _05232_ _05237_ net502 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__mux2_1
XANTENNA_32 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ top.cb_syn.char_path_n\[82\] net385 net335 top.cb_syn.char_path_n\[80\] net188
+ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05457_ net23 net413 net362 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 _02401_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ top.cb_syn.char_path_n\[116\] net198 _04650_ vssd1 vssd1 vccd1 vccd1 _01735_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05877__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05388_ top.cw2\[7\] vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__inv_2
XANTENNA__07658__A top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__A0 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07127_ _03796_ _03799_ _03801_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__nand4_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ _02459_ _02484_ _03722_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09592__B net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06009_ _02917_ _02921_ top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05943__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ clknet_leaf_48_clk net1072 _00361_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08428__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ clknet_leaf_120_clk _02088_ _00913_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11454_ clknet_leaf_87_clk _02019_ _00844_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_10405_ net746 net581 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__and2_1
XANTENNA__08948__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11385_ clknet_leaf_15_clk _01950_ _00775_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09783__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10336_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__and2_1
X_10267_ net718 net553 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06411__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05816__A top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05529__A3 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ net817 net652 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__and2_1
XANTENNA__05934__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06360_ _02600_ _03076_ _03226_ _02578_ top.findLeastValue.histo_index\[0\] vssd1
+ vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a32o_1
X_06291_ net458 _03147_ _03152_ _02607_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05311_ top.compVal\[24\] vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__inv_2
X_08030_ top.CB_read_complete top.cb_syn.setup vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__nand2_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
Xhold803 top.cb_syn.char_path_n\[29\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xinput41 gpio_in[7] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08939__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold836 top.cb_syn.zeroes\[4\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold814 top.cb_syn.char_path_n\[105\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold825 top.compVal\[23\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 top.histogram.total\[17\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ net755 net590 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__and2_1
X_08932_ _04239_ _04254_ _05059_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09364__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07417__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07914__B2 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout193_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08863_ net509 _05037_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__or2_1
X_08794_ top.path\[78\] top.path\[79\] net511 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__mux2_1
X_07814_ net435 net1492 net249 top.findLeastValue.sum\[35\] _04377_ vssd1 vssd1 vccd1
+ vccd1 _01824_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ _02519_ net387 _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout458_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ net967 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__clkbuf_1
X_07676_ top.hTree.tree_reg\[60\] _04248_ net387 vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06627_ _03414_ _03423_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o21ai_1
X_09346_ top.hTree.node_reg\[31\] net220 net214 _04391_ vssd1 vssd1 vccd1 vccd1 _01279_
+ sky130_fd_sc_hd__a22o_1
X_06558_ _03326_ net1609 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__nor2_1
X_05509_ _02416_ net453 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__nand2_1
X_09277_ net344 _04053_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[8\] sky130_fd_sc_hd__and2_1
X_06489_ _02454_ _03321_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__or2_1
X_08228_ top.cb_syn.char_path_n\[90\] net190 _04676_ vssd1 vssd1 vccd1 vccd1 _01709_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08159_ top.cb_syn.char_path_n\[125\] net369 net326 top.cb_syn.char_path_n\[123\]
+ net173 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a221o_1
X_11170_ clknet_leaf_55_clk _01735_ _00560_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10121_ net829 net664 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__and2_1
XANTENNA__06956__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ clknet_leaf_70_clk _01519_ _00344_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ clknet_leaf_23_clk top.header_synthesis.next_header\[7\] _00275_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05695__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11506_ clknet_leaf_118_clk _02071_ _00896_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06406__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11437_ clknet_leaf_95_clk _02002_ _00827_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[41\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08621__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ clknet_leaf_43_clk _01933_ _00758_ vssd1 vssd1 vccd1 vccd1 top.cw1\[0\] sky130_fd_sc_hd__dfrtp_2
X_10319_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09346__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ clknet_leaf_4_clk _01864_ _00689_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_05860_ net439 top.WB.prev_BUSY_O _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__and3_1
XANTENNA__07761__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07372__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05791_ top.sram_interface.zero_cnt\[2\] top.sram_interface.zero_cnt\[1\] _02818_
+ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__and3_1
X_07530_ _04128_ _04129_ net290 vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06096__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09071__C_N _02915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07461_ top.dut.bits_in_buf\[1\] net393 _04062_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__and3_1
X_06412_ top.hist_data_o\[29\] _03263_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nor2_1
X_07392_ _03824_ _03835_ _03833_ _03826_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_17_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09200_ _05181_ _05182_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__nor2_1
X_06343_ net534 _03206_ _03208_ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09131_ top.sram_interface.word_cnt\[9\] net545 _02587_ net460 vssd1 vssd1 vccd1
+ vccd1 _05139_ sky130_fd_sc_hd__o211a_1
X_09062_ net463 _04191_ _04556_ _05092_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a31o_1
XANTENNA__10346__B net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06274_ _02507_ _03079_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout206_A _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold611 top.hist_data_o\[13\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold600 top.hTree.tree_reg\[23\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
X_08013_ net1699 _04518_ _04519_ net254 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08531__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold644 top.cb_syn.count\[5\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 top.hTree.tree_reg\[14\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 top.hTree.tree_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 top.hist_data_o\[14\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 top.cw1\[2\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 top.dut.out\[0\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__and2_1
XANTENNA__09337__B1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold699 top.compVal\[5\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
X_09895_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__and2_1
X_08915_ top.cb_syn.max_index\[7\] _05061_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout575_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ net1103 _05034_ _05032_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__mux2_1
XANTENNA__09362__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06166__A3 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05890__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _04938_ _04964_ _04965_ _04940_ net504 vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a221o_1
X_05989_ top.WB.CPU_DAT_O\[12\] net1208 net348 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout742_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05903__B _02538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07728_ net472 _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__nand2_1
X_07659_ _04248_ net388 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__nand2_2
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ clknet_leaf_110_clk _01301_ _00060_ vssd1 vssd1 vccd1 vccd1 top.path\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_09329_ net1025 net227 net218 _04459_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08441__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ clknet_leaf_106_clk _01787_ _00612_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_FINISHED
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06929__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ clknet_leaf_63_clk _01718_ _00543_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10272__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ clknet_leaf_37_clk _01649_ _00474_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__and2_1
XANTENNA__09780__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__and2_1
XANTENNA__08551__A1 top.cb_syn.char_path_n\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10937_ clknet_leaf_54_clk _01502_ _00327_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ clknet_leaf_26_clk top.header_synthesis.next_enable _00258_ vssd1 vssd1 vccd1
+ vccd1 top.header_synthesis.enable sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ clknet_leaf_18_clk _01402_ _00189_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07814__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05840__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout409 net411 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
X_06961_ net407 net287 net149 net142 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__a31o_1
X_08700_ _04896_ _04897_ _04895_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a21oi_1
X_05912_ _02892_ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__nor2_1
X_09680_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__and2_1
X_08631_ top.cb_syn.char_path_n\[41\] top.cb_syn.char_path_n\[42\] top.cb_syn.char_path_n\[45\]
+ top.cb_syn.char_path_n\[46\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__mux4_1
X_06892_ top.findLeastValue.val2\[8\] net130 net121 _03651_ vssd1 vssd1 vccd1 vccd1
+ _02016_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_68_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05843_ _02832_ _02836_ _02864_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__and3_1
X_08562_ net519 net515 top.cb_syn.curr_state\[5\] _02895_ vssd1 vssd1 vccd1 vccd1
+ _04784_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_68_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05774_ top.compVal\[34\] net162 net147 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ _02319_ sky130_fd_sc_hd__a22o_1
X_07513_ top.cb_syn.char_path_n\[110\] top.cb_syn.char_path_n\[109\] top.cb_syn.char_path_n\[112\]
+ top.cb_syn.char_path_n\[111\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__mux4_1
X_08493_ net1423 top.cb_syn.char_path_n\[66\] net232 vssd1 vssd1 vccd1 vccd1 _01549_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07444_ _04050_ _04051_ net393 vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout323_A _04917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ _03851_ _04013_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__nand2_1
X_06326_ _03053_ _03194_ _02585_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__a21oi_1
X_09114_ net444 _05124_ _02417_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a21o_1
X_06257_ top.cb_syn.char_index\[3\] top.cb_syn.char_index\[2\] top.cb_syn.char_index\[1\]
+ top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a31o_1
X_09045_ top.WB.CPU_DAT_O\[5\] net1406 net315 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06188_ _03024_ _03061_ _02877_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__o21a_1
Xhold441 net101 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 top.path\[93\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 top.path\[79\] vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 top.path\[117\] vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold474 top.hTree.nulls\[52\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 top.hTree.tree_reg\[15\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 net90 vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
X_09947_ net794 net629 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__and2_1
X_09878_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__and2_1
X_08829_ net503 _05011_ _05014_ top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1
+ _05018_ sky130_fd_sc_hd__o31a_1
X_11840_ clknet_leaf_113_clk _02373_ _01212_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11771_ clknet_leaf_74_clk net991 vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_10722_ clknet_leaf_17_clk _01353_ _00112_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08436__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10653_ clknet_leaf_80_clk _01284_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ net797 net632 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ clknet_leaf_30_clk _01770_ _00595_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11136_ clknet_leaf_54_clk _01701_ _00526_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[82\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05586__A1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05586__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ clknet_leaf_59_clk _01632_ _00457_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07515__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05490_ top.findLeastValue.histo_index\[7\] net482 _02573_ _02574_ vssd1 vssd1 vccd1
+ vccd1 _02575_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_63_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07160_ _03826_ _03833_ _03835_ _03824_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o211a_1
X_06111_ _02997_ _03004_ _03008_ _02996_ net1595 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07091_ _03763_ _03764_ _03765_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__nand3_1
XANTENNA__09685__B net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06042_ top.sram_interface.init_counter\[1\] top.sram_interface.init_counter\[0\]
+ _02610_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout206 _04615_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
X_09801_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__and2_1
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08763__B2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ net847 net682 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__and2_1
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_4
X_07993_ net431 top.WorR _04520_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a21o_1
X_06944_ top.findLeastValue.val1\[13\] net136 net116 top.compVal\[13\] vssd1 vssd1
+ vccd1 vccd1 _01974_ sky130_fd_sc_hd__o22a_1
XANTENNA__09307__A3 top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__and2_1
X_06875_ top.compVal\[16\] top.findLeastValue.val1\[16\] net155 vssd1 vssd1 vccd1
+ vccd1 _03643_ sky130_fd_sc_hd__mux2_1
X_08614_ top.cb_syn.end_cnt\[3\] _04833_ _04830_ top.cb_syn.end_cnt\[4\] vssd1 vssd1
+ vccd1 vccd1 _04834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05453__B top.WB.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09594_ net726 net561 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__and2_1
X_05826_ top.sram_interface.counter_HTREE\[1\] top.sram_interface.counter_HTREE\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__or2_1
X_08545_ net1179 top.cb_syn.char_path_n\[14\] net245 vssd1 vssd1 vccd1 vccd1 _01497_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout538_A top.sram_interface.word_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05757_ _02794_ _02796_ _02800_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__and3b_1
X_08476_ net1184 top.cb_syn.char_path_n\[83\] net243 vssd1 vssd1 vccd1 vccd1 _01566_
+ sky130_fd_sc_hd__mux2_1
X_05688_ top.hTree.node_reg\[39\] net307 _02745_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout705_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07427_ top.findLeastValue.least1\[1\] net140 _03660_ net1143 vssd1 vssd1 vccd1 vccd1
+ _01870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07358_ net272 _04002_ _04003_ net278 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1
+ vccd1 _01902_ sky130_fd_sc_hd__a32o_1
X_06309_ net445 _03053_ _03178_ top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1
+ _03179_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07254__A1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ net270 _03951_ _03952_ net276 net1715 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a32o_1
XANTENNA__05909__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ top.WB.CPU_DAT_O\[22\] net1107 net314 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
Xhold271 top.hTree.nulls\[48\] vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 net88 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 top.hTree.node_reg\[54\] vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 net70 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 net749 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout751 net753 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_2
Xfanout773 net776 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout784 net786 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_2
Xfanout762 net777 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10550__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_2
XFILLER_0_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11823_ clknet_leaf_65_clk _02356_ _01195_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11754_ clknet_leaf_105_clk _00024_ _01144_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10705_ clknet_leaf_73_clk _01336_ _00095_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ clknet_leaf_100_clk _02235_ _01075_ vssd1 vssd1 vccd1 vccd1 top.compVal\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_10636_ clknet_leaf_73_clk _01267_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ net862 net697 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__and2_1
X_10498_ net751 net586 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11119_ clknet_leaf_49_clk _01684_ _00509_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[65\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10460__A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_11953__916 vssd1 vssd1 vccd1 vccd1 _11953__916/HI net916 sky130_fd_sc_hd__conb_1
XFILLER_0_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06660_ _03426_ _03454_ _03457_ _03427_ _03413_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o32a_1
X_05611_ top.cb_syn.char_path\[19\] net548 net539 top.cb_syn.char_path\[83\] vssd1
+ vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06591_ _02843_ _02852_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__nand2_1
X_08330_ top.cb_syn.char_path_n\[39\] net201 _04727_ vssd1 vssd1 vccd1 vccd1 _01658_
+ sky130_fd_sc_hd__o21a_1
X_05542_ top.histogram.sram_out\[31\] net360 net411 top.hTree.node_reg\[31\] vssd1
+ vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
X_08261_ top.cb_syn.char_path_n\[74\] net380 net337 top.cb_syn.char_path_n\[72\] net183
+ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05473_ net6 net413 net363 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 _02385_
+ sky130_fd_sc_hd__o22a_1
X_07212_ _03886_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__nand2_1
X_08192_ net1772 net203 _04658_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__o21a_1
X_07143_ _02477_ _02498_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_76_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout119_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07074_ _03742_ _03749_ _03744_ _03743_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or4b_2
XFILLER_0_112_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06025_ _02931_ _02934_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__nor2_1
XANTENNA__06995__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ top.findLeastValue.sum\[2\] _04506_ net391 vssd1 vssd1 vccd1 vccd1 _04507_
+ sky130_fd_sc_hd__mux2_1
X_09715_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__and2_1
X_06927_ top.findLeastValue.val1\[30\] net133 net115 top.compVal\[30\] vssd1 vssd1
+ vccd1 vccd1 _01991_ sky130_fd_sc_hd__o22a_1
XANTENNA__08595__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout655_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06858_ top.findLeastValue.val2\[25\] net127 net117 _03634_ vssd1 vssd1 vccd1 vccd1
+ _02033_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05809_ _02829_ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__nor2_1
X_09577_ net800 net635 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__and2_1
X_06789_ _03568_ _03569_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__and2b_1
X_08528_ net1297 top.cb_syn.char_path_n\[31\] net231 vssd1 vssd1 vccd1 vccd1 _01514_
+ sky130_fd_sc_hd__mux2_1
X_08459_ net1213 top.cb_syn.char_path_n\[100\] net239 vssd1 vssd1 vccd1 vccd1 _01583_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07570__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ clknet_leaf_102_clk _02035_ _00860_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10421_ net739 net574 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__and2_1
XANTENNA__10545__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10352_ net719 net554 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__and2_1
X_10283_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_2
Xfanout592 net631 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08586__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05961__B2 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07702__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ clknet_leaf_83_clk _02339_ _01178_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11913__944 vssd1 vssd1 vccd1 vccd1 net944 _11913__944/LO sky130_fd_sc_hd__conb_1
X_11737_ clknet_leaf_107_clk _02287_ _01127_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ clknet_leaf_91_clk _02218_ _01058_ vssd1 vssd1 vccd1 vccd1 top.compVal\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10619_ clknet_leaf_83_clk _01250_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11599_ clknet_leaf_0_clk top.dut.bit_buf_next\[6\] _00989_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08570__D net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07830_ top.hTree.tree_reg\[31\] top.findLeastValue.sum\[31\] net282 vssd1 vssd1
+ vccd1 vccd1 _04390_ sky130_fd_sc_hd__mux2_1
X_07761_ net478 _04333_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09143__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__and2_1
X_06712_ top.compVal\[41\] _02457_ _02458_ top.compVal\[40\] vssd1 vssd1 vccd1 vccd1
+ _03510_ sky130_fd_sc_hd__a22o_1
XANTENNA__05952__B2 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07692_ net474 _04276_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06643_ _03431_ _03437_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__or3_1
X_09431_ net755 net590 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06574_ top.header_synthesis.count\[2\] top.header_synthesis.count\[1\] top.header_synthesis.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__or3_1
X_09362_ net1488 _05255_ net228 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
X_08313_ top.cb_syn.char_path_n\[48\] net382 net332 top.cb_syn.char_path_n\[46\] net185
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a221o_1
X_05525_ net481 net453 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout236_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ net504 _05233_ _05235_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_25_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08244_ net1752 net199 _04684_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__o21a_1
XANTENNA__07552__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05456_ net25 net415 net364 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 _02402_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_33 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ top.cb_syn.char_path_n\[117\] net377 net334 top.cb_syn.char_path_n\[115\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a221o_1
X_05387_ top.findLeastValue.histo_index\[0\] vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout403_A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ top.findLeastValue.val2\[13\] top.findLeastValue.val1\[13\] vssd1 vssd1 vccd1
+ vccd1 _03802_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08709__A1 top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07057_ _03725_ _03726_ _03728_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__or4_2
XFILLER_0_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06008_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07393__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__D_N top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ net436 net1573 net250 top.findLeastValue.sum\[6\] _04493_ vssd1 vssd1 vccd1
+ vccd1 _01795_ sky130_fd_sc_hd__a221o_1
XANTENNA__05943__B2 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ clknet_leaf_55_clk net1137 _00360_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_09629_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_50_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
X_11522_ clknet_leaf_120_clk _02087_ _00912_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11453_ clknet_leaf_87_clk _02018_ _00843_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_10404_ net746 net581 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__and2_1
X_11384_ clknet_leaf_15_clk _01949_ _00774_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06959__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10335_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__and2_1
XANTENNA__06899__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05631__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10266_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__and2_1
XANTENNA__07908__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05816__B net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ net817 net652 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__and2_1
XANTENNA__07384__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05934__B2 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07687__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05698__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06290_ net461 _03160_ _03158_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05310_ top.compVal\[25\] vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__inv_2
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput42 gpio_in[8] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold837 top.cb_syn.char_path_n\[92\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 top.cb_syn.char_path_n\[22\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold804 top.cb_syn.char_path_n\[113\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 net94 vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 top.hTree.node_reg\[60\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06414__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09980_ net754 net589 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__and2_1
X_08931_ _05073_ top.cb_syn.max_index\[3\] _05059_ vssd1 vssd1 vccd1 vccd1 _01403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08167__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08862_ _05043_ _05045_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__or2_1
X_07813_ net418 _04375_ _04376_ net260 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_4_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09116__A1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08793_ _02547_ _04976_ _04980_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__o22a_1
XANTENNA__08529__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ net387 _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07675_ net449 net1039 _04257_ _04264_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o22a_1
X_09414_ net971 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06626_ _02430_ top.findLeastValue.val1\[22\] _02492_ top.compVal\[21\] vssd1 vssd1
+ vccd1 vccd1 _03424_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06350__B2 top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_A top.cb_syn.char_path_n\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
X_09345_ top.hTree.node_reg\[30\] net220 net214 _04395_ vssd1 vssd1 vccd1 vccd1 _01278_
+ sky130_fd_sc_hd__a22o_1
X_06557_ top.histogram.total\[2\] _03325_ net1608 vssd1 vssd1 vccd1 vccd1 _03362_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05508_ net481 _02417_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__nor2_1
X_09276_ net343 _04054_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[7\] sky130_fd_sc_hd__and2_1
X_06488_ top.dut.out_valid top.histogram.out_of_init vssd1 vssd1 vccd1 vccd1 _03321_
+ sky130_fd_sc_hd__and2b_1
X_08227_ top.cb_syn.char_path_n\[91\] net369 net326 top.cb_syn.char_path_n\[89\] net173
+ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a221o_1
X_05439_ top.cb_syn.zero_count\[0\] vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08158_ top.cb_syn.char_path_n\[125\] net192 _04641_ vssd1 vssd1 vccd1 vccd1 _01744_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\] vssd1 vssd1 vccd1 vccd1
+ _04591_ sky130_fd_sc_hd__nand2_1
X_07109_ _03784_ _03776_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__nand2b_1
XANTENNA__05613__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05917__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__and2_1
XANTENNA__08158__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_99_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08439__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold732_A top.findLeastValue.sum\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ clknet_leaf_70_clk _01518_ _00343_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ clknet_leaf_23_clk top.header_synthesis.next_header\[6\] _00274_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[6\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_23_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06892__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07579__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ clknet_leaf_119_clk _02070_ _00895_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11436_ clknet_leaf_95_clk _02001_ _00826_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[40\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09043__A0 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ clknet_leaf_94_clk _01932_ _00757_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[45\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07518__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06422__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10318_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09346__A1 top.hTree.node_reg\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11298_ clknet_leaf_5_clk _01863_ _00688_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ net753 net588 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__and2_1
X_05790_ _02816_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__nand2b_1
X_11919__950 vssd1 vssd1 vccd1 vccd1 net950 _11919__950/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_37_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07460_ net342 net393 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__nor2_1
XANTENNA__08609__B1 _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06411_ net1251 _03274_ net301 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
X_07391_ _03839_ net271 _04025_ net277 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1
+ vccd1 _01891_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_17_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06342_ _02600_ _03078_ _03209_ _02578_ net487 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_14_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_09130_ net1517 _05138_ _05134_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__a21o_1
X_09061_ net424 _02969_ _02995_ net523 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08012_ _04530_ net1672 _04522_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__mux2_1
X_06273_ _02601_ _03141_ _03143_ net534 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 top.hTree.tree_reg\[21\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 top.histogram.total\[17\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09034__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold623 top.histogram.wr_r_en\[0\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 top.hTree.tree_reg\[33\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 top.histogram.total\[16\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__and2_1
Xhold667 top.hTree.nullSumIndex\[2\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 top.hTree.tree_reg\[38\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 top.hTree.node_reg\[28\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08914_ top.cb_syn.max_index\[6\] top.cb_syn.max_index\[5\] _05060_ vssd1 vssd1 vccd1
+ vccd1 _05061_ sky130_fd_sc_hd__and3_1
Xhold689 top.sram_interface.counter_HTREE\[2\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
X_09894_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ net513 _05033_ net423 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__o21ai_1
X_08776_ top.path\[16\] net403 _04917_ top.path\[17\] _02547_ vssd1 vssd1 vccd1 vccd1
+ _04965_ sky130_fd_sc_hd__o221a_1
X_07727_ _02516_ net387 _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__o21a_1
X_05988_ top.WB.CPU_DAT_O\[13\] net1441 net348 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ top.hTree.write_HT_fin top.hTree.closing vssd1 vssd1 vccd1 vccd1 _04250_
+ sky130_fd_sc_hd__or2_1
X_07589_ _02993_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06609_ top.compVal\[39\] top.compVal\[38\] top.compVal\[37\] top.compVal\[36\] vssd1
+ vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__or4_1
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06874__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ net989 net226 net217 _04463_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _02559_ _05216_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07823__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09025__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10553__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ clknet_leaf_106_clk net1005 _00611_ vssd1 vssd1 vccd1 vccd1 top.HT_fin_reg
+ sky130_fd_sc_hd__dfrtp_1
X_11152_ clknet_leaf_64_clk _01717_ _00542_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[98\]
+ sky130_fd_sc_hd__dfrtp_4
X_10103_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__and2_1
XANTENNA__08023__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083_ clknet_leaf_36_clk _01648_ _00473_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_10034_ net785 net620 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__and2_1
XANTENNA__07862__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10936_ clknet_leaf_54_clk _01501_ _00326_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10867_ clknet_leaf_14_clk _01453_ _00257_ vssd1 vssd1 vccd1 vccd1 top.hTree.finish_check
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07801__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06417__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10798_ clknet_leaf_18_clk _01401_ _00188_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07814__B2 top.findLeastValue.sum\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07814__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11419_ clknet_leaf_76_clk _01984_ _00809_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[23\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_117_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08775__C1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ _02499_ net125 net123 _03663_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08790__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_05911_ top.cb_syn.h_element\[61\] top.cb_syn.h_element\[60\] top.cb_syn.h_element\[59\]
+ top.cb_syn.h_element\[62\] vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__or4b_1
X_06891_ top.compVal\[8\] top.findLeastValue.val1\[8\] net154 vssd1 vssd1 vccd1 vccd1
+ _03651_ sky130_fd_sc_hd__mux2_1
XANTENNA__05991__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ _04846_ _04849_ _02541_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__mux2_1
X_05842_ _02849_ net440 top.hTree.state\[8\] _02853_ vssd1 vssd1 vccd1 vccd1 _02864_
+ sky130_fd_sc_hd__and4b_1
X_08561_ _04197_ _04609_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_68_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05773_ top.compVal\[35\] net162 net147 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ _02320_ sky130_fd_sc_hd__a22o_1
X_07512_ _02980_ _02984_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__xor2_1
X_08492_ net1094 top.cb_syn.char_path_n\[67\] net237 vssd1 vssd1 vccd1 vccd1 _01550_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07443_ top.dut.bit_buf\[9\] top.dut.bit_buf\[2\] net713 vssd1 vssd1 vccd1 vccd1
+ _04051_ sky130_fd_sc_hd__mux2_1
XANTENNA__06856__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ _03851_ _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__or2_1
X_09113_ _02417_ net1750 _05129_ _02416_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06325_ top.TRN_char_index\[1\] top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 _03194_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07947__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06256_ net481 _03125_ _03127_ _03019_ net454 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__o221a_1
X_09044_ top.WB.CPU_DAT_O\[6\] net1315 net316 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
Xhold420 top.hTree.tree_reg\[63\] vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 top.cb_syn.char_path\[98\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ top.sram_interface.init_counter\[7\] _03023_ top.sram_interface.init_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__a21oi_1
Xhold442 top.path\[95\] vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 top.path\[116\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 top.cb_syn.char_path\[29\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 _01804_ vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 top.hTree.node_reg\[20\] vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09946_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__and2_1
Xhold497 top.histogram.total\[29\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08828_ _02546_ _04982_ _05015_ _05016_ top.translation.index\[6\] vssd1 vssd1 vccd1
+ vccd1 _05017_ sky130_fd_sc_hd__a221o_1
X_08759_ net425 _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__or2_1
X_11770_ clknet_leaf_45_clk _02309_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10721_ clknet_leaf_40_clk _01352_ _00111_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07621__S _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10548__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10652_ clknet_leaf_79_clk _01283_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ net745 net580 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07857__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11204_ clknet_leaf_30_clk _01769_ _00594_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07576__B _04175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ clknet_leaf_58_clk _01700_ _00525_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[81\]
+ sky130_fd_sc_hd__dfrtp_2
X_11066_ clknet_leaf_60_clk _01631_ _00456_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05586__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06299__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10919_ clknet_leaf_48_clk _01484_ _00309_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11899_ net930 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XANTENNA__10458__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06838__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06110_ _02448_ _03002_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__nand2_1
XANTENNA__07767__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ _03764_ _03765_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__nand2_1
X_06041_ net444 top.sram_interface.init_counter\[10\] top.WB.prev_BUSY_O top.sram_interface.init_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_2_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06471__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08212__A1 top.cb_syn.char_path_n\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05287__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__and2_1
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
Xfanout229 _05252_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
X_07992_ top.hTree.state\[4\] top.hTree.state\[3\] _04519_ net254 vssd1 vssd1 vccd1
+ vccd1 _04520_ sky130_fd_sc_hd__o31a_1
XANTENNA__08763__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 _02620_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
X_09731_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06943_ top.findLeastValue.val1\[14\] net139 net116 top.compVal\[14\] vssd1 vssd1
+ vccd1 vccd1 _01975_ sky130_fd_sc_hd__o22a_1
X_09662_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__and2_1
X_06874_ top.findLeastValue.val2\[17\] net128 net121 _03642_ vssd1 vssd1 vccd1 vccd1
+ _02025_ sky130_fd_sc_hd__o22a_1
X_08613_ _04831_ _04832_ net496 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__mux2_1
X_05825_ _02846_ _02842_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__nand2b_1
XANTENNA__05453__C net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ net742 net577 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__and2_1
X_08544_ net1080 top.cb_syn.char_path_n\[15\] net243 vssd1 vssd1 vccd1 vccd1 _01498_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08279__A1 top.cb_syn.char_path_n\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05756_ _02576_ _02798_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__nand2_1
XANTENNA__08537__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ net1231 top.cb_syn.char_path_n\[84\] net242 vssd1 vssd1 vccd1 vccd1 _01567_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout433_A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05687_ top.histogram.sram_out\[7\] net357 net408 top.hTree.node_reg\[7\] vssd1 vssd1
+ vccd1 vccd1 _02746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07426_ top.findLeastValue.least1\[2\] net141 _03660_ top.findLeastValue.histo_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07357_ _03795_ _04001_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__nand2_1
X_06308_ _02589_ _03049_ _03177_ _03054_ net545 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a32o_1
X_07288_ _03885_ _03944_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_1
X_09027_ top.WB.CPU_DAT_O\[23\] net1205 net313 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
X_06239_ top.cb_syn.char_index\[5\] _03035_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__or2_1
XANTENNA__08739__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07408__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 top.hTree.nulls\[54\] vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 top.path\[40\] vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top.cb_syn.char_path\[81\] vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 top.path\[71\] vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 top.path\[123\] vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05568__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net732 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_2
Xfanout741 net749 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_2
Xfanout774 net776 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_2
X_09929_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__and2_1
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_2
Xfanout763 net766 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_2
Xfanout752 net753 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10550__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout796 net34 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_4
X_11822_ clknet_leaf_66_clk _02355_ _01194_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ clknet_leaf_105_clk net1523 _01143_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ clknet_leaf_45_clk _01335_ _00094_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ clknet_leaf_94_clk _02234_ _01074_ vssd1 vssd1 vccd1 vccd1 top.compVal\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ clknet_leaf_69_clk _01266_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10566_ net864 net699 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10497_ net755 net590 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07526__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ clknet_leaf_50_clk _01683_ _00508_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09155__C1 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ clknet_leaf_24_clk _01614_ _00439_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[3\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_05610_ net1477 net169 _02681_ net211 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06590_ top.header_synthesis.bit1 _03388_ _03389_ _03384_ vssd1 vssd1 vccd1 vccd1
+ _02056_ sky130_fd_sc_hd__a31o_1
XANTENNA__05731__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05541_ _02622_ _02623_ net465 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__o21a_1
X_08260_ top.cb_syn.char_path_n\[74\] net203 _04692_ vssd1 vssd1 vccd1 vccd1 _01693_
+ sky130_fd_sc_hd__o21a_1
X_05472_ net7 net415 net364 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 _02386_
+ sky130_fd_sc_hd__a22o_1
X_08191_ top.cb_syn.char_path_n\[109\] net383 net339 top.cb_syn.char_path_n\[107\]
+ net186 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a221o_1
X_07211_ top.findLeastValue.val2\[32\] top.findLeastValue.val1\[32\] vssd1 vssd1 vccd1
+ vccd1 _03887_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07142_ top.findLeastValue.val2\[5\] top.findLeastValue.val1\[5\] vssd1 vssd1 vccd1
+ vccd1 _03818_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07073_ _03747_ _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nand2_1
X_06024_ top.sram_interface.init_counter\[7\] _02930_ top.sram_interface.init_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08820__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11927__890 vssd1 vssd1 vccd1 vccd1 _11927__890/HI net890 sky130_fd_sc_hd__conb_1
XFILLER_0_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08736__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07944__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ top.hTree.tree_reg\[2\] top.findLeastValue.sum\[2\] net284 vssd1 vssd1 vccd1
+ vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_98_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09714_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__and2_1
X_06926_ top.findLeastValue.val1\[31\] net133 net114 net1762 vssd1 vssd1 vccd1 vccd1
+ _01992_ sky130_fd_sc_hd__o22a_1
XANTENNA__08595__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ net762 net597 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__and2_1
X_06857_ top.compVal\[25\] top.findLeastValue.val1\[25\] net150 vssd1 vssd1 vccd1
+ vccd1 _03634_ sky130_fd_sc_hd__mux2_1
X_05808_ _02523_ top.findLeastValue.least1\[6\] top.findLeastValue.least1\[5\] top.findLeastValue.least1\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout648_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ net798 net633 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__and2_1
X_06788_ _02433_ top.findLeastValue.val2\[16\] _03560_ _03563_ _03585_ vssd1 vssd1
+ vccd1 vccd1 _03586_ sky130_fd_sc_hd__a2111oi_1
X_08527_ net1193 top.cb_syn.char_path_n\[32\] net232 vssd1 vssd1 vccd1 vccd1 _01515_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10098__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05739_ top.findLeastValue.histo_index\[8\] _02575_ vssd1 vssd1 vccd1 vccd1 _02783_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ net1242 top.cb_syn.char_path_n\[101\] net239 vssd1 vssd1 vccd1 vccd1 _01584_
+ sky130_fd_sc_hd__mux2_1
X_07409_ net485 top.findLeastValue.least1\[4\] net150 vssd1 vssd1 vccd1 vccd1 _04035_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05486__B2 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08389_ top.cb_syn.char_path_n\[10\] net380 net337 top.cb_syn.char_path_n\[8\] net183
+ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
X_10420_ net739 net574 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_21_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10545__B net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__and2_1
X_10282_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__and2_1
XANTENNA__08730__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_2
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_2
Xfanout571 net631 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_4
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08586__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05713__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ clknet_leaf_83_clk _02338_ _01177_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
X_11736_ clknet_leaf_7_clk _02286_ _01126_ vssd1 vssd1 vccd1 vccd1 top.histogram.init
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_60_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05477__B2 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ clknet_leaf_91_clk _02217_ _01057_ vssd1 vssd1 vccd1 vccd1 top.compVal\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06425__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10618_ clknet_leaf_83_clk _01249_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11598_ clknet_leaf_120_clk top.dut.bit_buf_next\[5\] _00988_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ net834 net669 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__and2_1
XANTENNA__10471__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07760_ top.hTree.tree_reg\[45\] top.findLeastValue.sum\[45\] net267 vssd1 vssd1
+ vccd1 vccd1 _04334_ sky130_fd_sc_hd__mux2_1
X_06711_ _02406_ top.findLeastValue.val2\[45\] _02455_ top.compVal\[44\] vssd1 vssd1
+ vccd1 vccd1 _03509_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__05952__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07691_ net474 _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand2_1
X_09430_ net755 net590 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06642_ _02440_ top.findLeastValue.val1\[6\] _03430_ _03438_ vssd1 vssd1 vccd1 vccd1
+ _03440_ sky130_fd_sc_hd__a211o_1
X_06573_ top.header_synthesis.count\[7\] top.header_synthesis.count\[6\] top.header_synthesis.count\[5\]
+ top.header_synthesis.count\[4\] vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__or4_1
X_09361_ top.hTree.nulls\[46\] _04331_ net398 vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08312_ top.cb_syn.char_path_n\[48\] net196 _04718_ vssd1 vssd1 vccd1 vccd1 _01667_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05524_ net450 _02524_ net533 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__and3_1
X_09292_ top.histogram.total\[24\] net402 net323 top.histogram.total\[25\] net429
+ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__o221a_1
X_08243_ top.cb_syn.char_path_n\[83\] net378 net335 top.cb_syn.char_path_n\[81\] net181
+ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__a221o_1
XANTENNA_23 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05468__B2 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05455_ net26 net414 net363 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 _02403_
+ sky130_fd_sc_hd__o22a_1
X_08174_ net1710 net198 _04649_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__o21a_1
XANTENNA__08406__A1 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05386_ net483 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__inv_2
X_07125_ top.findLeastValue.val2\[13\] top.findLeastValue.val1\[13\] vssd1 vssd1 vccd1
+ vccd1 _03801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07056_ _03730_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06007_ top.translation.totalEn _02814_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11895__926 vssd1 vssd1 vccd1 vccd1 net926 _11895__926/LO sky130_fd_sc_hd__conb_1
X_07958_ net418 _04491_ _04492_ net261 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o211a_1
XANTENNA__05943__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ net435 net1395 net248 top.findLeastValue.sum\[20\] _04437_ vssd1 vssd1 vccd1
+ vccd1 _01809_ sky130_fd_sc_hd__a221o_1
X_06909_ net288 net140 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__nor2_2
X_09628_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__and2_1
XANTENNA__07696__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A1 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09559_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05459__B2 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold608_A top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ clknet_leaf_119_clk _02086_ _00911_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10556__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11452_ clknet_leaf_88_clk _02017_ _00842_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_11383_ clknet_leaf_9_clk _01948_ _00773_ vssd1 vssd1 vccd1 vccd1 top.cw2\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09070__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ net747 net582 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__and2_1
X_10334_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__and2_1
XANTENNA__09070__B2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10265_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__and2_1
XANTENNA__05385__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ net817 net652 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__and2_1
Xfanout390 net392 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
XANTENNA__05934__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08884__A1 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11719_ clknet_leaf_73_clk _02269_ _01109_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05870__A1 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 gpio_in[9] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xhold816 top.cb_syn.char_path_n\[84\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold805 top.cb_syn.char_path_n\[51\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 top.controller.fin_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold838 top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
X_08930_ _04234_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09364__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ net402 _05037_ net504 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_4_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07812_ net476 _04374_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__or2_1
X_08792_ top.translation.index\[2\] _04977_ net503 vssd1 vssd1 vccd1 vccd1 _04981_
+ sky130_fd_sc_hd__a21o_1
X_07743_ top.hTree.tree_reg\[48\] top.findLeastValue.least2\[2\] net280 vssd1 vssd1
+ vccd1 vccd1 _04320_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout179_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _04262_ _04263_ net474 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__mux2_1
XANTENNA__05742__B top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__A1 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ net968 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06886__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06625_ top.compVal\[20\] _02493_ _03417_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout346_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09344_ net1795 net220 net214 _04399_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__a22o_1
X_06556_ _03327_ _03361_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__nor2_1
X_05507_ _02585_ _02591_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__nand2_1
X_06487_ _02420_ net1454 net297 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
X_09275_ _04072_ _05226_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[6\] sky130_fd_sc_hd__and2_1
X_08226_ net1721 net190 _04675_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__o21a_1
X_05438_ net463 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ top.cb_syn.char_path_n\[126\] net370 net328 top.cb_syn.char_path_n\[124\]
+ net174 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a221o_1
XANTENNA__09884__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07108_ _03780_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__nand2_1
X_05369_ top.findLeastValue.val1\[37\] vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__inv_2
X_08088_ net519 net514 _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_95_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07039_ top.findLeastValue.val1\[22\] top.findLeastValue.val1\[21\] top.findLeastValue.val1\[20\]
+ top.findLeastValue.val1\[19\] vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__and4_1
XANTENNA__09355__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10952_ clknet_leaf_47_clk net1355 _00342_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08866__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10883_ clknet_leaf_23_clk top.header_synthesis.next_header\[5\] _00273_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07579__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ clknet_leaf_120_clk _02069_ _00894_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11435_ clknet_leaf_95_clk _02000_ _00825_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[39\]
+ sky130_fd_sc_hd__dfstp_1
X_11366_ clknet_leaf_93_clk _01931_ _00756_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[44\]
+ sky130_fd_sc_hd__dfrtp_2
X_10317_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__and2_1
X_11297_ clknet_leaf_2_clk _01862_ _00687_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10248_ net819 net654 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__and2_1
X_10179_ net810 net645 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__and2_1
XANTENNA__07534__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__A1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06410_ top.hist_data_o\[30\] _03264_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__xor2_1
XANTENNA__05989__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05540__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07390_ _03820_ _03822_ _03823_ _03836_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_17_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06341_ _02510_ _03076_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06272_ _03072_ _03142_ _02601_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__o21ai_1
X_09060_ net1588 _05089_ _05090_ net1542 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08011_ top.findLeastValue.least2\[0\] top.findLeastValue.least1\[0\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 _01810_ vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 top.hTree.tree_reg\[8\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 top.hist_addr\[5\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 _01822_ vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__and2_1
Xhold679 top.findLeastValue.sum\[19\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 top.hTree.tree_reg\[54\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 top.histogram.total\[14\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 top.histogram.total\[3\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
X_08913_ top.cb_syn.max_index\[4\] top.cb_syn.max_index\[3\] top.cb_syn.max_index\[2\]
+ top.cb_syn.max_index\[1\] vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__and4_1
X_09893_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__and2_1
X_08844_ _02813_ _05028_ top.translation.totalEn vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__o21ba_1
X_05987_ top.WB.CPU_DAT_O\[14\] net1256 net347 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
X_08775_ top.path\[24\] net402 net323 top.path\[25\] net502 vssd1 vssd1 vccd1 vccd1
+ _04964_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout463_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ net387 _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ net449 net282 net1000 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a21o_1
X_07588_ _02972_ _04106_ _02971_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__o21a_1
X_06608_ top.compVal\[43\] top.compVal\[42\] top.compVal\[41\] top.compVal\[40\] vssd1
+ vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__or4_1
X_09327_ net979 net226 net218 _04467_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06539_ net1597 _03333_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__xor2_1
XANTENNA__07808__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07284__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08209_ top.cb_syn.char_path_n\[100\] net379 net336 top.cb_syn.char_path_n\[98\]
+ net182 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a221o_1
X_09189_ top.hTree.state\[3\] net254 _05121_ net1637 vssd1 vssd1 vccd1 vccd1 _00020_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ clknet_leaf_43_clk _01785_ _00610_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ clknet_leaf_46_clk _01716_ _00541_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[97\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07587__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07587__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10553__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05598__B1 _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09328__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__and2_1
X_11082_ clknet_leaf_36_clk _01647_ _00472_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08631__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__and2_1
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05770__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ clknet_leaf_58_clk net1199 _00325_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10866_ clknet_leaf_28_clk top.header_synthesis.next_zero_count\[7\] _00256_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07275__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10797_ clknet_leaf_3_clk _00002_ _00187_ vssd1 vssd1 vccd1 vccd1 top.WB.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ clknet_leaf_76_clk _01983_ _00808_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[22\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_117_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08775__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05589__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11349_ clknet_leaf_103_clk _01914_ _00739_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921__885 vssd1 vssd1 vccd1 vccd1 _11921__885/HI net885 sky130_fd_sc_hd__conb_1
X_05910_ top.cb_syn.h_element\[58\] top.cb_syn.h_element\[57\] top.cb_syn.h_element\[56\]
+ top.cb_syn.h_element\[55\] vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__or4_1
X_06890_ top.findLeastValue.val2\[9\] net130 net120 _03650_ vssd1 vssd1 vccd1 vccd1
+ _02017_ sky130_fd_sc_hd__o22a_1
X_05841_ net544 _02861_ net448 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08560_ net515 top.cb_syn.curr_state\[5\] _04178_ _04607_ net464 vssd1 vssd1 vccd1
+ vccd1 _04782_ sky130_fd_sc_hd__o311a_1
X_05772_ top.compVal\[36\] net162 net147 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ _02321_ sky130_fd_sc_hd__a22o_1
XANTENNA__05761__B1 _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ _02975_ _04101_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__xnor2_2
X_08491_ net1120 top.cb_syn.char_path_n\[68\] net237 vssd1 vssd1 vccd1 vccd1 _01551_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07442_ top.dut.bit_buf\[10\] top.dut.bit_buf\[3\] net714 vssd1 vssd1 vccd1 vccd1
+ _04050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07373_ top.findLeastValue.val2\[8\] top.findLeastValue.val1\[8\] _03850_ vssd1 vssd1
+ vccd1 vccd1 _04013_ sky130_fd_sc_hd__a21o_1
X_06324_ _03042_ _03192_ _02605_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09112_ _03369_ _05122_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__nor2_1
XANTENNA__08823__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06255_ _03023_ _03126_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nor2_1
X_09043_ top.WB.CPU_DAT_O\[7\] net1183 net315 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 _01525_ vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08215__C1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06186_ net1548 net164 _03060_ net207 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold454 top.hTree.node_reg\[48\] vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 net80 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07666__C net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 top.path\[74\] vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08766__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 top.path\[124\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 top.cb_syn.count\[3\] vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 top.cb_syn.char_path\[49\] vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _01512_ vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06241__A1 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__and2_1
Xhold498 _03345_ vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
X_09876_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__and2_1
XANTENNA__07682__B _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ _02547_ _04996_ _04999_ top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1
+ _05016_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout845_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ top.path\[86\] top.path\[87\] net508 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__mux2_1
X_08689_ _04886_ _04879_ top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__mux2_1
X_07709_ net475 _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nand2_1
X_10720_ clknet_leaf_17_clk _01351_ _00110_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_109_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10548__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ clknet_leaf_80_clk _01282_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ net745 net580 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10564__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ clknet_leaf_30_clk _01768_ _00593_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08221__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ clknet_leaf_58_clk _01699_ _00524_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[80\]
+ sky130_fd_sc_hd__dfrtp_2
X_11065_ clknet_leaf_60_clk _01630_ _00455_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05991__A0 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A1 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net830 net665 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08288__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ clknet_leaf_46_clk _01483_ _00308_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11898_ net929 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XANTENNA__10458__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849_ clknet_leaf_117_clk _01443_ _00239_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_119_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08996__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__B2 top.findLeastValue.sum\[38\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06040_ top.sram_interface.init_counter\[9\] top.sram_interface.init_counter\[8\]
+ top.sram_interface.init_counter\[7\] top.sram_interface.init_counter\[6\] vssd1
+ vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout208 _02620_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
Xfanout219 _05254_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
X_07991_ top.hTree.state\[5\] top.hTree.state\[2\] vssd1 vssd1 vccd1 vccd1 _04519_
+ sky130_fd_sc_hd__or2_1
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__and2_1
XANTENNA__05982__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06942_ top.findLeastValue.val1\[15\] net138 net116 top.compVal\[15\] vssd1 vssd1
+ vccd1 vccd1 _01976_ sky130_fd_sc_hd__o22a_1
X_09661_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__and2_1
X_06873_ top.compVal\[17\] top.findLeastValue.val1\[17\] net152 vssd1 vssd1 vccd1
+ vccd1 _03642_ sky130_fd_sc_hd__mux2_1
X_08612_ top.cb_syn.char_path_n\[19\] top.cb_syn.char_path_n\[20\] top.cb_syn.char_path_n\[23\]
+ top.cb_syn.char_path_n\[24\] net499 net493 vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__mux4_1
X_05824_ top.hTree.state\[6\] top.hTree.state\[9\] vssd1 vssd1 vccd1 vccd1 _02846_
+ sky130_fd_sc_hd__nor2_1
X_09592_ net723 net558 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__and2_1
X_08543_ net1104 top.cb_syn.char_path_n\[16\] net243 vssd1 vssd1 vccd1 vccd1 _01499_
+ sky130_fd_sc_hd__mux2_1
X_05755_ _02576_ _02798_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout259_A _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_A _02908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08474_ net1269 top.cb_syn.char_path_n\[85\] net235 vssd1 vssd1 vccd1 vccd1 _01568_
+ sky130_fd_sc_hd__mux2_1
X_05686_ _02743_ _02744_ net468 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07425_ top.findLeastValue.least1\[3\] net141 _03660_ net1615 vssd1 vssd1 vccd1 vccd1
+ _01872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout426_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ _03795_ _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__or2_1
XANTENNA__08987__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06307_ net445 top.TRN_char_index\[1\] vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__or2_1
X_07287_ _03885_ _03944_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06238_ top.cb_syn.char_index\[5\] _03046_ _03110_ vssd1 vssd1 vccd1 vccd1 _03111_
+ sky130_fd_sc_hd__o21a_1
X_09026_ top.WB.CPU_DAT_O\[24\] net1294 net313 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout795_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 top.cb_syn.char_path\[100\] vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 top.hTree.tree_reg\[56\] vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
X_06169_ top.cb_syn.char_index\[3\] top.cb_syn.char_index\[2\] _03042_ vssd1 vssd1
+ vccd1 vccd1 _03044_ sky130_fd_sc_hd__and3_1
Xhold251 top.path\[115\] vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold284 top.cb_syn.char_path\[86\] vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _01564_ vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 top.path\[12\] vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__and2_1
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_1
Xfanout720 net736 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_1
Xfanout742 net749 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_2
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_2
Xfanout764 net766 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05973__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout753 net796 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09859_ net867 net702 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__and2_1
Xfanout786 net795 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07714__A1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout797 net803 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07714__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ clknet_leaf_66_clk _02354_ _01193_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10559__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08029__A top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ clknet_leaf_105_clk _00022_ _01142_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10703_ clknet_leaf_46_clk _01334_ _00093_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_11683_ clknet_leaf_100_clk _02233_ _01073_ vssd1 vssd1 vccd1 vccd1 top.compVal\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_10634_ clknet_leaf_73_clk _01265_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ net862 net697 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__and2_1
XANTENNA__06453__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10496_ net755 net590 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07402__A0 top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ clknet_leaf_50_clk _01682_ _00507_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[63\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07953__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ clknet_leaf_24_clk _01613_ _00438_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[2\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07705__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05540_ top.cb_syn.char_path\[63\] net528 net309 top.cb_syn.char_path\[127\] vssd1
+ vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05471_ net8 net413 net362 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 _02387_
+ sky130_fd_sc_hd__o22a_1
X_08190_ top.cb_syn.char_path_n\[109\] net203 _04657_ vssd1 vssd1 vccd1 vccd1 _01728_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05997__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07210_ top.findLeastValue.val2\[32\] top.findLeastValue.val1\[32\] vssd1 vssd1 vccd1
+ vccd1 _03886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07141_ top.findLeastValue.val2\[5\] top.findLeastValue.val1\[5\] vssd1 vssd1 vccd1
+ vccd1 _03817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09993__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ top.findLeastValue.val2\[28\] top.findLeastValue.val1\[28\] vssd1 vssd1 vccd1
+ vccd1 _03748_ sky130_fd_sc_hd__or2_1
X_06023_ _02932_ _02933_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__and2_1
XANTENNA__05798__A3 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07944__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__B2 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ net436 net1229 net250 top.findLeastValue.sum\[3\] _04505_ vssd1 vssd1 vccd1
+ vccd1 _01792_ sky130_fd_sc_hd__a221o_1
X_09713_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__and2_1
X_06925_ top.findLeastValue.val1\[32\] net133 net114 top.compVal\[32\] vssd1 vssd1
+ vccd1 vccd1 _01993_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout376_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ net762 net597 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__and2_1
X_06856_ top.findLeastValue.val2\[26\] net126 net117 _03633_ vssd1 vssd1 vccd1 vccd1
+ _02034_ sky130_fd_sc_hd__o22a_1
X_05807_ top.findLeastValue.least1\[3\] top.findLeastValue.least1\[2\] top.findLeastValue.least1\[1\]
+ top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_2_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ net799 net634 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__and2_1
X_06787_ top.compVal\[19\] _02469_ _02470_ top.compVal\[18\] _03584_ vssd1 vssd1 vccd1
+ vccd1 _03585_ sky130_fd_sc_hd__o221ai_1
X_08526_ net1324 top.cb_syn.char_path_n\[33\] net237 vssd1 vssd1 vccd1 vccd1 _01516_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10098__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05738_ top.TRN_char_index\[0\] net38 net715 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XANTENNA__07555__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06132__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ net1216 top.cb_syn.char_path_n\[102\] net239 vssd1 vssd1 vccd1 vccd1 _01585_
+ sky130_fd_sc_hd__mux2_1
X_05669_ top.histogram.sram_out\[10\] net357 net408 top.hTree.node_reg\[10\] vssd1
+ vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07408_ _02516_ net125 net124 _04034_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout808_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05486__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ top.cb_syn.char_path_n\[10\] net203 _04756_ vssd1 vssd1 vccd1 vccd1 _01629_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06592__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07339_ _03773_ _03977_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__nand2b_1
X_10350_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10281_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__and2_1
X_09009_ _03364_ _05079_ _05080_ net453 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__o31ai_4
XANTENNA__07627__S _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
XANTENNA__05946__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_2
Xfanout572 net575 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_2
Xfanout561 net571 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout594 net612 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_29_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ clknet_leaf_4_clk _02337_ _01176_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_11735_ clknet_leaf_12_clk _02285_ _01125_ vssd1 vssd1 vccd1 vccd1 top.FLV_done sky130_fd_sc_hd__dfrtp_1
X_11666_ clknet_leaf_18_clk _02216_ _01056_ vssd1 vssd1 vccd1 vccd1 top.CB_read_complete
+ sky130_fd_sc_hd__dfrtp_2
X_10617_ clknet_leaf_83_clk _01248_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ clknet_leaf_120_clk top.dut.bit_buf_next\[4\] _00987_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08921__S _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ net834 net669 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__and2_1
XANTENNA__07537__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09376__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ net841 net676 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__and2_1
XANTENNA__10471__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05937__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _03412_ net149 net288 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__a21o_1
X_07690_ top.findLeastValue.least1\[3\] net264 _04275_ vssd1 vssd1 vccd1 vccd1 _04277_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06641_ _03430_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand2b_1
X_06572_ top.header_synthesis.enable top.header_synthesis.write_char_path top.header_synthesis.char_added
+ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__and3_1
X_09360_ net969 net226 net218 _04334_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__a22o_1
X_08311_ top.cb_syn.char_path_n\[49\] net375 net333 top.cb_syn.char_path_n\[47\] net178
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a221o_1
X_05523_ net460 net545 _02604_ net458 _02607_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a221o_1
X_09291_ net425 _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__or2_1
X_08242_ net1720 net198 _04683_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__o21a_1
X_05454_ net72 net415 top.WB.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__or3b_1
XANTENNA_13 gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ top.cb_syn.char_path_n\[118\] net377 net330 top.cb_syn.char_path_n\[116\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__a221o_1
XANTENNA__08406__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05385_ net482 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__inv_2
X_07124_ _02473_ _02495_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07055_ top.findLeastValue.val2\[36\] top.findLeastValue.val1\[36\] vssd1 vssd1 vccd1
+ vccd1 _03731_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05640__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09367__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06006_ net441 net513 _02919_ _02807_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__or4b_1
XFILLER_0_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ net477 _04490_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__or2_1
XANTENNA__07393__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ top.findLeastValue.val2\[0\] net130 net120 _03659_ vssd1 vssd1 vccd1 vccd1
+ _02008_ sky130_fd_sc_hd__o22a_1
XANTENNA__08342__A1 top.cb_syn.char_path_n\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ net421 _04435_ _04436_ net260 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o211a_1
X_09627_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__and2_1
X_06839_ top.compVal\[34\] top.findLeastValue.val1\[34\] net152 vssd1 vssd1 vccd1
+ vccd1 _03625_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09898__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07528__S0 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ net1129 top.cb_syn.char_path_n\[50\] net242 vssd1 vssd1 vccd1 vccd1 _01533_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__and2_1
XANTENNA__05459__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ clknet_leaf_119_clk _02085_ _00910_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10556__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ clknet_leaf_87_clk _02016_ _00841_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[8\]
+ sky130_fd_sc_hd__dfstp_2
X_11382_ clknet_leaf_19_clk _01947_ _00772_ vssd1 vssd1 vccd1 vccd1 top.cw2\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08802__C1 _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ net747 net582 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__and2_1
XANTENNA__08741__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10333_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__and2_1
XANTENNA__06959__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943__906 vssd1 vssd1 vccd1 vccd1 _11943__906/HI net906 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_111_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10572__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__and2_1
X_10195_ net805 net640 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__and2_1
XANTENNA__07384__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout380 net382 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08916__S _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07820__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06436__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ clknet_leaf_73_clk _02268_ _01108_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07844__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ clknet_leaf_115_clk _02199_ _01039_ vssd1 vssd1 vccd1 vccd1 top.path\[48\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 nrst vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
Xhold806 top.sram_interface.init_counter\[7\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 top.cw1\[4\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold817 top.compVal\[9\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 top.hist_data_o\[15\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09349__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ net502 _05043_ _05044_ _05039_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__o22a_1
XANTENNA__08572__B2 top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07811_ top.findLeastValue.sum\[35\] _04374_ net391 vssd1 vssd1 vccd1 vccd1 _04375_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08791_ net426 _04978_ _04979_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__o21a_1
X_07742_ net257 _04318_ _04319_ net1010 net432 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a32o_1
X_07673_ top.findLeastValue.least1\[6\] _04262_ net389 vssd1 vssd1 vccd1 vccd1 _04263_
+ sky130_fd_sc_hd__mux2_1
X_09412_ net958 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05689__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06624_ _03415_ _03418_ _03420_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__a22o_1
X_09343_ net1629 net220 net214 _04403_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout241_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06555_ net1668 _03326_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05506_ net451 _02589_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__nand2_2
X_06486_ net1410 net297 _03245_ _03320_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22o_1
X_09274_ _04057_ _05226_ _04076_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[5\]
+ sky130_fd_sc_hd__o21a_1
X_08225_ top.cb_syn.char_path_n\[92\] net369 net327 top.cb_syn.char_path_n\[90\] net173
+ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a221o_1
X_05437_ net523 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08156_ net1771 net192 _04640_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__o21a_1
X_05368_ top.findLeastValue.val1\[38\] vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__inv_2
X_07107_ _03781_ _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ _04196_ _04549_ _04587_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__or4b_4
X_05299_ net481 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__inv_2
XANTENNA__10392__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07038_ top.findLeastValue.val1\[30\] top.findLeastValue.val1\[29\] top.findLeastValue.val1\[28\]
+ top.findLeastValue.val1\[27\] vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903__934 vssd1 vssd1 vccd1 vccd1 net934 _11903__934/LO sky130_fd_sc_hd__conb_1
X_08989_ top.WB.CPU_DAT_O\[31\] net1301 net366 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ clknet_leaf_47_clk _01516_ _00341_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10882_ clknet_leaf_23_clk top.header_synthesis.next_header\[4\] _00272_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10567__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ clknet_leaf_120_clk _02068_ _00893_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11434_ clknet_leaf_95_clk _01999_ _00824_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[38\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__08471__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11365_ clknet_leaf_93_clk _01930_ _00755_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[43\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_100_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10316_ net731 net566 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__and2_1
X_11296_ clknet_leaf_2_clk _01861_ _00686_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ net819 net654 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__and2_1
XANTENNA__07815__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07550__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06340_ _03070_ _03207_ _02601_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06271_ top.cw1\[4\] _03071_ top.cw1\[5\] vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08010_ _04529_ net1657 _04522_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold603 top.cb_syn.char_path\[89\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold625 top.histogram.sram_out\[10\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 top.hTree.tree_reg\[25\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 net52 vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold647 top.cb_syn.h_element\[62\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A1 _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold658 _03362_ vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 top.dut.out\[1\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ _02866_ _05055_ _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__or4_4
X_09892_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout191_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _05024_ _05029_ _05030_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout289_A _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08774_ net430 _04943_ _04946_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__or3_1
X_05986_ top.WB.CPU_DAT_O\[15\] net1236 net347 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
X_07725_ top.hTree.tree_reg\[51\] top.findLeastValue.least2\[5\] net280 vssd1 vssd1
+ vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ top.findLeastValue.least2\[8\] top.findLeastValue.least1\[8\] _02837_ _04247_
+ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__and4_2
XANTENNA_fanout623_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ net521 _04177_ _04186_ net516 vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06607_ _03401_ _03402_ _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ net1017 net226 net217 _04471_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__a22o_1
X_06538_ _03353_ _03354_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__nor2_1
X_09257_ _02559_ _05216_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__nor2_1
XANTENNA__07284__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ net1770 net200 _04666_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__o21a_1
X_06469_ net298 _03249_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07284__B2 top.findLeastValue.sum\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ _02866_ _05176_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__or2_1
XANTENNA__08233__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\] top.cb_syn.cb_length\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o21ai_1
X_11150_ clknet_leaf_40_clk _01715_ _00540_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[96\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__and2_1
X_11081_ clknet_leaf_36_clk _01646_ _00471_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08631__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__and2_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05770__B2 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ clknet_leaf_58_clk _01499_ _00324_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ clknet_leaf_28_clk top.header_synthesis.next_zero_count\[6\] _00255_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11949__912 vssd1 vssd1 vccd1 vccd1 _11949__912/HI net912 sky130_fd_sc_hd__conb_1
XANTENNA__07275__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10796_ clknet_leaf_3_clk _00001_ _00186_ vssd1 vssd1 vccd1 vccd1 top.WB.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11417_ clknet_leaf_78_clk _01982_ _00807_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[21\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_117_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11348_ clknet_leaf_75_clk _01913_ _00738_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__A1 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ clknet_leaf_44_clk _01844_ _00669_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_05840_ net526 net536 top.sram_interface.word_cnt\[13\] net446 vssd1 vssd1 vccd1
+ vccd1 _02862_ sky130_fd_sc_hd__o31a_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _02991_ _04102_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__xnor2_4
X_05771_ top.compVal\[37\] net162 net147 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ _02322_ sky130_fd_sc_hd__a22o_1
X_08490_ net1086 top.cb_syn.char_path_n\[69\] net237 vssd1 vssd1 vccd1 vccd1 _01552_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ net393 vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf_next\[0\] sky130_fd_sc_hd__inv_2
X_07372_ top.findLeastValue.sum\[10\] net278 net272 _04012_ vssd1 vssd1 vccd1 vccd1
+ _01897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06323_ top.cb_syn.char_index\[1\] top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1
+ _03192_ sky130_fd_sc_hd__nand2_1
X_09111_ top.histogram.state\[0\] _05126_ _05127_ _05128_ vssd1 vssd1 vccd1 vccd1
+ _00028_ sky130_fd_sc_hd__a211o_1
X_06254_ top.sram_interface.init_counter\[6\] _03022_ vssd1 vssd1 vccd1 vccd1 _03126_
+ sky130_fd_sc_hd__nor2_1
X_09042_ top.WB.CPU_DAT_O\[8\] net1459 net315 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold411 top.cb_syn.char_path\[74\] vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ _03033_ _03059_ _03041_ _03048_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__or4b_1
Xhold400 _01808_ vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 top.cb_syn.char_path\[27\] vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 top.hTree.tree_reg\[20\] vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold422 top.path\[98\] vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 top.cb_syn.curr_index\[6\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 top.path\[101\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 top.sram_interface.zero_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__and2_1
Xhold488 top.cb_syn.char_path\[91\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 top.hTree.tree_reg\[44\] vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_09875_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__and2_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08826_ net505 _05000_ _05002_ _05003_ net503 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout838_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ net428 _04944_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout740_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05969_ net452 net536 _02913_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__nand3_1
X_08688_ _04880_ _04886_ _04892_ _04879_ net1688 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a32o_1
X_07708_ top.findLeastValue.least1\[0\] net264 _04290_ vssd1 vssd1 vccd1 vccd1 _04292_
+ sky130_fd_sc_hd__a21oi_1
X_07639_ net521 _04231_ _04234_ net516 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10650_ clknet_leaf_80_clk _01281_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09309_ top.translation.resEn top.translation.totalEn _02807_ _05028_ vssd1 vssd1
+ vccd1 vccd1 top.controller.fin_TRN sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_101_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10581_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10564__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909__940 vssd1 vssd1 vccd1 vccd1 net940 _11909__940/LO sky130_fd_sc_hd__conb_1
X_11202_ clknet_leaf_30_clk _01767_ _00592_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08757__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__B top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ clknet_leaf_58_clk _01698_ _00523_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_11064_ clknet_leaf_60_clk _01629_ _00454_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_10015_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06940__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ clknet_leaf_39_clk _01482_ _00307_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_found
+ sky130_fd_sc_hd__dfrtp_1
X_11897_ net928 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08924__S _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10848_ clknet_leaf_117_clk _01442_ _00238_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_119_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ clknet_leaf_118_clk _01385_ _00169_ vssd1 vssd1 vccd1 vccd1 top.path\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout209 net212 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_07990_ top.hTree.state\[4\] top.hTree.state\[3\] net255 vssd1 vssd1 vccd1 vccd1
+ _04518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06941_ top.findLeastValue.val1\[16\] net138 net115 top.compVal\[16\] vssd1 vssd1
+ vccd1 vccd1 _01977_ sky130_fd_sc_hd__o22a_1
X_09660_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__and2_1
X_08611_ top.cb_syn.char_path_n\[17\] top.cb_syn.char_path_n\[18\] top.cb_syn.char_path_n\[21\]
+ top.cb_syn.char_path_n\[22\] net499 net493 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__mux4_1
X_06872_ top.findLeastValue.val2\[18\] net131 net122 _03641_ vssd1 vssd1 vccd1 vccd1
+ _02026_ sky130_fd_sc_hd__o22a_1
XANTENNA__05734__A1 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05823_ _02844_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__inv_2
X_09591_ net723 net558 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__and2_1
XANTENNA__06931__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ net1198 top.cb_syn.char_path_n\[17\] net243 vssd1 vssd1 vccd1 vccd1 _01500_
+ sky130_fd_sc_hd__mux2_1
X_05754_ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__inv_2
X_08473_ net1235 top.cb_syn.char_path_n\[86\] net235 vssd1 vssd1 vccd1 vccd1 _01569_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07487__A1 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08119__B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05685_ top.cb_syn.char_path\[39\] net529 net310 top.cb_syn.char_path\[103\] vssd1
+ vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
X_07424_ top.findLeastValue.least1\[4\] net141 _03660_ net485 vssd1 vssd1 vccd1 vccd1
+ _01873_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07355_ _03791_ _04000_ _03790_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a21bo_1
X_06306_ top.cb_syn.char_index\[2\] _03042_ _03175_ net465 vssd1 vssd1 vccd1 vccd1
+ _03176_ sky130_fd_sc_hd__o211a_1
X_07286_ net270 _03946_ _03950_ net276 top.findLeastValue.sum\[34\] vssd1 vssd1 vccd1
+ vccd1 _01921_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout419_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06998__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06237_ _02605_ _03047_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__nor2_1
XANTENNA__06462__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09025_ top.WB.CPU_DAT_O\[25\] net1194 net313 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
XANTENNA__05670__B1 _02730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold252 top.cb_syn.char_path\[103\] vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ top.cb_syn.char_index\[2\] _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__nand2_1
Xhold241 top.hTree.nulls\[58\] vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 top.path\[109\] vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
X_06099_ _02451_ _02998_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout788_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 top.cb_syn.char_path\[64\] vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 top.header_synthesis.header\[5\] vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _01583_ vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 top.path\[47\] vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__and2_1
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_2
Xfanout732 net736 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_2
Xfanout721 net723 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08598__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_1
Xfanout743 net748 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_2
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_2
X_09858_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__and2_1
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_2
Xfanout798 net803 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_1
X_09789_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06922__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ top.path\[41\] net325 _04997_ net426 net430 vssd1 vssd1 vccd1 vccd1 _04998_
+ sky130_fd_sc_hd__o221a_1
X_11820_ clknet_leaf_65_clk _02353_ _01192_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10559__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ clknet_leaf_104_clk _00021_ _01141_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_44_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ clknet_leaf_47_clk _01333_ _00092_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[46\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_80_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08744__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11682_ clknet_leaf_94_clk _02232_ _01072_ vssd1 vssd1 vccd1 vccd1 top.compVal\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ clknet_leaf_69_clk _01264_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ net862 net697 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05661__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ net732 net567 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ clknet_leaf_38_clk _01681_ _00506_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[62\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05964__A1 top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09155__B2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ clknet_leaf_24_clk _01612_ _00437_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08902__A1 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06913__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__B1 _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_71_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
X_11949_ net912 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
X_05470_ net9 net413 net363 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 _02388_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08761__S0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ top.findLeastValue.val2\[10\] top.findLeastValue.val1\[10\] _03808_ _03815_
+ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09993__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07071_ top.findLeastValue.val2\[28\] top.findLeastValue.val1\[28\] vssd1 vssd1 vccd1
+ vccd1 _03747_ sky130_fd_sc_hd__nand2_1
XANTENNA__05652__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06022_ top.sram_interface.init_counter\[9\] _02931_ vssd1 vssd1 vccd1 vccd1 _02933_
+ sky130_fd_sc_hd__or2_1
X_09712_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__and2_1
XANTENNA__05955__B2 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ net419 _04503_ _04504_ net261 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__o211a_1
X_06924_ top.findLeastValue.val1\[33\] net133 net114 net1775 vssd1 vssd1 vccd1 vccd1
+ _01994_ sky130_fd_sc_hd__o22a_1
X_09643_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout271_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06855_ top.compVal\[26\] top.findLeastValue.val1\[26\] net150 vssd1 vssd1 vccd1
+ vccd1 _03633_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout369_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06904__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ net747 net582 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__and2_1
XANTENNA__05707__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05806_ net1633 _02825_ _02828_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__o21a_1
X_08525_ net1354 top.cb_syn.char_path_n\[34\] net232 vssd1 vssd1 vccd1 vccd1 _01517_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06349__S top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06786_ _03579_ _03582_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
X_05737_ top.TRN_char_index\[1\] net39 net715 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XANTENNA__07555__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05668_ _02728_ _02729_ net468 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__o21a_1
X_08456_ net1203 top.cb_syn.char_path_n\[103\] net239 vssd1 vssd1 vccd1 vccd1 _01586_
+ sky130_fd_sc_hd__mux2_1
X_08387_ top.cb_syn.char_path_n\[11\] net383 net339 top.cb_syn.char_path_n\[9\] net186
+ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a221o_1
X_07407_ net483 top.findLeastValue.least1\[5\] net149 vssd1 vssd1 vccd1 vccd1 _04034_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07688__B _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05599_ top.cb_syn.char_path\[21\] net548 net539 top.cb_syn.char_path\[85\] vssd1
+ vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout703_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ net269 _03979_ _03988_ net275 net1624 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_21_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07632__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07632__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ _03724_ _03934_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
XANTENNA__05643__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ net444 _02405_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nor2_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
Xfanout551 net553 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05946__B2 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout584 net631 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_2
Xfanout573 net575 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_2
Xfanout562 net564 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08345__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net597 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07699__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09424__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08360__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11803_ clknet_leaf_5_clk _02336_ _01175_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08474__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11734_ clknet_leaf_12_clk _02284_ _01124_ vssd1 vssd1 vccd1 vccd1 top.hTree.write_HT_fin
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09132__A_N _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ clknet_leaf_19_clk _02215_ _01055_ vssd1 vssd1 vccd1 vccd1 top.CB_write_complete
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_10616_ net718 net553 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ clknet_leaf_5_clk top.dut.bit_buf_next\[3\] _00986_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[3\] sky130_fd_sc_hd__dfrtp_1
X_10547_ net832 net667 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10478_ net841 net676 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05937__B2 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07553__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06640_ _02439_ top.findLeastValue.val1\[7\] top.findLeastValue.val1\[6\] _02440_
+ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__o22ai_1
X_06571_ top.header_synthesis.write_char_path top.header_synthesis.start vssd1 vssd1
+ vccd1 vccd1 _03371_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08310_ top.cb_syn.char_path_n\[49\] net196 _04717_ vssd1 vssd1 vccd1 vccd1 _01668_
+ sky130_fd_sc_hd__o21a_1
X_05522_ _02588_ net309 net461 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__o21a_2
X_09290_ top.histogram.total\[26\] top.histogram.total\[27\] net509 vssd1 vssd1 vccd1
+ vccd1 _05234_ sky130_fd_sc_hd__mux2_1
X_08241_ top.cb_syn.char_path_n\[84\] net377 net334 top.cb_syn.char_path_n\[82\] net180
+ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05453_ net440 top.WB.prev_BUSY_O net414 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__and3_1
XANTENNA_14 gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08172_ top.cb_syn.char_path_n\[118\] net193 _04648_ vssd1 vssd1 vccd1 vccd1 _01737_
+ sky130_fd_sc_hd__o21a_1
X_05384_ top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ _03797_ _03798_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__nor2_1
XANTENNA__05625__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA_fanout117_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ top.findLeastValue.val2\[36\] top.findLeastValue.val1\[36\] vssd1 vssd1 vccd1
+ vccd1 _03730_ sky130_fd_sc_hd__nand2_1
X_06005_ top.translation.write_fin top.TRN_sram_complete top.translation.totalEn vssd1
+ vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a21oi_1
X_07956_ top.hTree.tree_reg\[6\] top.findLeastValue.sum\[6\] net266 vssd1 vssd1 vccd1
+ vccd1 _04491_ sky130_fd_sc_hd__mux2_1
X_06907_ top.compVal\[0\] top.findLeastValue.val1\[0\] net154 vssd1 vssd1 vccd1 vccd1
+ _03659_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08342__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07887_ net476 _04434_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout653_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__and2_1
X_06838_ top.findLeastValue.val2\[35\] net128 net118 _03624_ vssd1 vssd1 vccd1 vccd1
+ _02043_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_26_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09898__B net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09557_ net763 net598 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06769_ _02427_ top.findLeastValue.val2\[25\] top.findLeastValue.val2\[24\] _02428_
+ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__o22a_1
XANTENNA__07528__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
X_08508_ net1121 top.cb_syn.char_path_n\[51\] net242 vssd1 vssd1 vccd1 vccd1 _01534_
+ sky130_fd_sc_hd__mux2_1
X_09488_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ net1079 top.cb_syn.char_path_n\[120\] net235 vssd1 vssd1 vccd1 vccd1 _01603_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07302__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07853__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ clknet_leaf_88_clk _02015_ _00840_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11381_ clknet_leaf_19_clk _01946_ _00771_ vssd1 vssd1 vccd1 vccd1 top.cw2\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08802__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10401_ net746 net581 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__and2_1
X_10332_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10572__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10263_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__and2_1
X_10194_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__and2_1
XANTENNA__08469__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout370 _04612_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout392 _04250_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11717_ clknet_leaf_70_clk _02267_ _01107_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_30_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07844__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ clknet_leaf_111_clk _02198_ _01038_ vssd1 vssd1 vccd1 vccd1 top.path\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09046__A0 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ clknet_leaf_6_clk _02144_ _00969_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05607__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold818 top.cb_syn.h_element\[58\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold807 top.hist_addr\[4\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 top.cb_syn.h_element\[56\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ top.hTree.tree_reg\[35\] top.findLeastValue.sum\[35\] net283 vssd1 vssd1
+ vccd1 vccd1 _04374_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08790_ top.path\[0\] net404 net324 top.path\[1\] net429 vssd1 vssd1 vccd1 vccd1
+ _04979_ sky130_fd_sc_hd__o221a_1
X_07741_ net473 _04315_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07672_ top.findLeastValue.least1\[6\] top.hTree.tree_reg\[61\] _04248_ vssd1 vssd1
+ vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
X_09411_ net961 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06886__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06623_ _02432_ top.findLeastValue.val1\[17\] _03419_ vssd1 vssd1 vccd1 vccd1 _03421_
+ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_17_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_09342_ net964 net220 net214 _04407_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__a22o_1
X_06554_ _03325_ _03328_ _03360_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a21oi_1
X_05505_ net451 _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_51_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout234_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ net343 _04067_ _04046_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__o21a_1
X_06485_ top.hist_data_o\[1\] top.hist_data_o\[0\] net300 vssd1 vssd1 vccd1 vccd1
+ _03320_ sky130_fd_sc_hd__o21a_1
X_08224_ net1788 net190 _04674_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__o21a_1
X_05436_ net544 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09037__A0 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08155_ top.cb_syn.char_path_n\[127\] net370 net328 top.cb_syn.char_path_n\[125\]
+ net174 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__a221o_1
X_05367_ top.findLeastValue.val1\[39\] vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__inv_2
X_07106_ top.findLeastValue.val2\[20\] top.findLeastValue.val1\[20\] vssd1 vssd1 vccd1
+ vccd1 _03782_ sky130_fd_sc_hd__or2_1
X_08086_ net519 net524 net514 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05298_ top.compVal\[32\] vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07037_ top.findLeastValue.val1\[26\] top.findLeastValue.val1\[25\] top.findLeastValue.val1\[24\]
+ top.findLeastValue.val1\[23\] vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout770_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net449 net528 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__nand2_1
X_07939_ net436 net1589 net251 top.findLeastValue.sum\[10\] _04477_ vssd1 vssd1 vccd1
+ vccd1 _01799_ sky130_fd_sc_hd__a221o_1
XANTENNA__08315__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ clknet_leaf_46_clk _01515_ _00340_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07921__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ clknet_leaf_23_clk top.header_synthesis.next_header\[3\] _00271_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[3\] sky130_fd_sc_hd__dfrtp_1
X_09609_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10567__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ clknet_leaf_120_clk _02067_ _00892_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08752__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09028__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ clknet_leaf_95_clk _01998_ _00823_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[37\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_59_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11364_ clknet_leaf_81_clk _01929_ _00754_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__and2_1
X_11295_ clknet_leaf_24_clk _01860_ _00685_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08988__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07406__A2_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10246_ net819 net654 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__and2_1
XANTENNA__08306__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05540__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06447__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06270_ _03091_ _03140_ net484 _02787_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06971__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09019__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10493__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__C1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 top.cb_syn.curr_path\[127\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold615 _01814_ vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 top.hist_data_o\[3\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09960_ net770 net605 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold648 top.hTree.tree_reg\[9\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 top.hTree.tree_reg\[39\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 top.hTree.state\[8\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_08911_ net449 _02838_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09891_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__and2_1
X_08842_ net423 top.header_synthesis.enable net36 net452 vssd1 vssd1 vccd1 vccd1 _05031_
+ sky130_fd_sc_hd__o211a_1
X_05985_ top.WB.CPU_DAT_O\[16\] net1299 net345 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
X_08773_ top.translation.index\[5\] _04957_ _04958_ _04961_ vssd1 vssd1 vccd1 vccd1
+ _04962_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07724_ net257 _04303_ _04304_ net1009 net432 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a32o_1
X_07655_ _02837_ _02853_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nand3_4
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout351_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ top.compVal\[19\] top.compVal\[18\] top.compVal\[17\] top.compVal\[16\] vssd1
+ vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07586_ top.cb_syn.max_index\[7\] _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ net995 net224 net216 _04475_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__a22o_1
X_06537_ net1803 _03333_ net1591 vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07808__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _05207_ _05216_ _05217_ _05208_ top.cb_syn.zero_count\[4\] vssd1 vssd1 vccd1
+ vccd1 top.header_synthesis.next_zero_count\[4\] sky130_fd_sc_hd__a32o_1
XANTENNA_fanout616_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ top.hist_data_o\[6\] _03246_ _03247_ top.hist_data_o\[7\] vssd1 vssd1 vccd1
+ vccd1 _03309_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_97_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08207_ top.cb_syn.char_path_n\[101\] net379 net336 top.cb_syn.char_path_n\[99\]
+ net182 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a221o_1
X_05419_ top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06399_ top.hist_data_o\[29\] _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__and2_1
X_09187_ top.hTree.state\[3\] _05057_ net256 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__mux2_1
XANTENNA__08769__C1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__A1 top.cb_syn.char_path_n\[88\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ top.cb_syn.cb_length\[2\] net190 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08069_ net1726 _04578_ _04575_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__o21a_1
X_11080_ clknet_leaf_52_clk _01645_ _00470_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07916__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ net814 net649 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__and2_1
X_10031_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__and2_1
XANTENNA__09135__C net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05770__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10933_ clknet_leaf_58_clk _01498_ _00323_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10864_ clknet_leaf_28_clk top.header_synthesis.next_zero_count\[5\] _00254_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__05522__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10795_ clknet_leaf_4_clk _00000_ _00185_ vssd1 vssd1 vccd1 vccd1 top.WB.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07887__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ clknet_leaf_78_clk _01981_ _00806_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[20\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_117_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11347_ clknet_leaf_76_clk _01912_ _00737_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08775__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ clknet_leaf_104_clk _01843_ _00668_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_10229_ net810 net645 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__and2_1
Xhold1 top.controller.fin_HG vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
X_05770_ top.compVal\[38\] net162 net147 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ _02323_ sky130_fd_sc_hd__a22o_1
XANTENNA__07561__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05761__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07440_ net714 top.dut.bits_in_buf\[0\] vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09996__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07371_ _03806_ _04008_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__xor2_1
X_06322_ top.cb_syn.max_index\[3\] _03102_ _03104_ top.hTree.nullSumIndex\[2\] vssd1
+ vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a22o_1
XANTENNA__07797__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ net439 top.histogram.state\[7\] _05124_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__and3_1
XANTENNA__08463__A1 top.cb_syn.char_path_n\[96\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06905__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09041_ top.WB.CPU_DAT_O\[9\] net1496 net315 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06253_ top.hist_addr\[6\] _03099_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__xor2_1
XANTENNA__08215__A1 top.cb_syn.char_path_n\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06184_ _03051_ _03058_ top.TRN_char_index\[6\] _02592_ vssd1 vssd1 vccd1 vccd1 _03059_
+ sky130_fd_sc_hd__o211a_1
Xhold401 top.path\[68\] vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold434 top.cb_syn.char_path\[65\] vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 top.hTree.node_reg\[19\] vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _01809_ vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 top.path\[89\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 top.histogram.sram_out\[31\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 top.path\[13\] vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 top.path\[99\] vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__and2_1
Xhold489 _01574_ vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09874_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08825_ top.path\[96\] net404 _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__o21a_1
XANTENNA__09191__A2 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ top.path\[20\] net403 net323 top.path\[21\] _02547_ vssd1 vssd1 vccd1 vccd1
+ _04945_ sky130_fd_sc_hd__o221a_1
XANTENNA__05780__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05968_ net452 net536 vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__nand2_1
X_08687_ top.cb_syn.i\[1\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07707_ top.hTree.tree_reg\[55\] top.findLeastValue.least1\[0\] net280 vssd1 vssd1
+ vccd1 vccd1 _04291_ sky130_fd_sc_hd__mux2_1
X_05899_ net461 top.sram_interface.word_cnt\[9\] net956 vssd1 vssd1 vccd1 vccd1 _02251_
+ sky130_fd_sc_hd__a21o_1
X_07638_ _04183_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nand2_1
X_07569_ top.cb_syn.char_path_n\[54\] top.cb_syn.char_path_n\[53\] top.cb_syn.char_path_n\[56\]
+ top.cb_syn.char_path_n\[55\] net394 net295 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09308_ _05250_ _05251_ vssd1 vssd1 vccd1 vccd1 top.translation.writeBin sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_101_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10580_ net799 net634 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09239_ net490 top.header_synthesis.header\[8\] vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11201_ clknet_leaf_29_clk _01766_ _00591_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_11132_ clknet_leaf_59_clk _01697_ _00522_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09427__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ clknet_leaf_61_clk _01628_ _00453_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_10014_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__and2_1
XANTENNA__08477__S net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ clknet_leaf_33_clk _01481_ _00306_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.left_check
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11896_ net927 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_94_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ clknet_leaf_2_clk _01441_ _00237_ vssd1 vssd1 vccd1 vccd1 top.translation.resEn
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10778_ clknet_leaf_113_clk _01384_ _00168_ vssd1 vssd1 vccd1 vccd1 top.path\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07556__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07420__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06940_ top.findLeastValue.val1\[17\] net137 net115 top.compVal\[17\] vssd1 vssd1
+ vccd1 vccd1 _01978_ sky130_fd_sc_hd__o22a_1
X_06871_ top.compVal\[18\] top.findLeastValue.val1\[18\] net155 vssd1 vssd1 vccd1
+ vccd1 _03641_ sky130_fd_sc_hd__mux2_1
X_08610_ _02542_ _04827_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a21o_1
X_05822_ _02840_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09590_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__and2_1
X_08541_ net1170 top.cb_syn.char_path_n\[18\] net246 vssd1 vssd1 vccd1 vccd1 _01501_
+ sky130_fd_sc_hd__mux2_1
X_05753_ top.sram_interface.write_counter_FLV\[1\] top.sram_interface.write_counter_FLV\[0\]
+ top.sram_interface.write_counter_FLV\[2\] vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__or3b_1
X_08472_ net1262 top.cb_syn.char_path_n\[87\] net236 vssd1 vssd1 vccd1 vccd1 _01570_
+ sky130_fd_sc_hd__mux2_1
X_05684_ top.cb_syn.char_path\[7\] net547 net540 top.cb_syn.char_path\[71\] vssd1
+ vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a22o_1
XANTENNA__09800__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07423_ top.findLeastValue.least1\[5\] net141 _03660_ net483 vssd1 vssd1 vccd1 vccd1
+ _01874_ sky130_fd_sc_hd__a22o_1
XANTENNA__05498__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A _02806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07354_ _03802_ _03999_ _03800_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__a21o_1
X_06305_ net545 _03043_ _03174_ _03034_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a22o_1
X_07285_ _03884_ _03945_ _03877_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout314_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06236_ _02591_ _03051_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__nor3_1
X_09024_ top.WB.CPU_DAT_O\[26\] net1279 net314 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
Xhold220 top.cb_syn.char_path\[21\] vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08739__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 top.cb_syn.char_path\[32\] vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 top.cb_syn.char_path\[3\] vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ top.cb_syn.char_index\[1\] top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1
+ _03042_ sky130_fd_sc_hd__or2_1
Xhold253 net65 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
X_06098_ top.cb_syn.count\[1\] top.cb_syn.count\[0\] vssd1 vssd1 vccd1 vccd1 _02998_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout683_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout700 net711 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_2
Xhold286 top.sram_interface.word_cnt\[7\] vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 net59 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 top.path\[86\] vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__and2_1
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_2
Xhold297 net98 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout722 net723 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__clkbuf_2
Xfanout733 net734 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08598__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 net777 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_2
Xfanout744 net748 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_1
Xfanout755 net757 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_2
X_09857_ net871 net706 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout850_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 net794 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_2
Xfanout777 net795 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_2
Xfanout799 net803 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_2
X_09788_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__and2_1
X_08808_ top.path\[42\] top.path\[43\] net511 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__mux2_1
XANTENNA__05725__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ top.path\[125\] net324 _04927_ net427 net505 vssd1 vssd1 vccd1 vccd1 _04928_
+ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_77_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ clknet_leaf_105_clk net1638 _01140_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10701_ clknet_leaf_7_clk _01332_ _00091_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06686__B1 top.findLeastValue.val1\[46\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07883__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ clknet_leaf_86_clk _02231_ _01071_ vssd1 vssd1 vccd1 vccd1 top.compVal\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10632_ clknet_leaf_64_clk _01263_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10563_ net861 net696 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ net752 net587 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ clknet_leaf_38_clk _01680_ _00505_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_11046_ clknet_leaf_24_clk _01611_ _00436_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08363__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ net911 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08761__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ net63 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ _03743_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__and2_1
X_06021_ net1518 _02932_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07929__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09394__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__and2_1
X_07972_ net477 _04502_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__or2_1
X_06923_ top.findLeastValue.val1\[34\] net133 net114 top.compVal\[34\] vssd1 vssd1
+ vccd1 vccd1 _01995_ sky130_fd_sc_hd__o22a_1
X_09642_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__and2_1
XANTENNA__06365__C1 top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05707__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ top.findLeastValue.val2\[27\] net127 net117 _03632_ vssd1 vssd1 vccd1 vccd1
+ _02035_ sky130_fd_sc_hd__o22a_1
X_09573_ net747 net582 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__and2_1
X_06785_ _03564_ _03578_ _03580_ _03581_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__and4_1
X_05805_ net1281 _02828_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__xnor2_1
X_08524_ net1111 top.cb_syn.char_path_n\[35\] net238 vssd1 vssd1 vccd1 vccd1 _01518_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout264_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05736_ net445 net40 net715 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XANTENNA__08657__B2 _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934__897 vssd1 vssd1 vccd1 vccd1 _11934__897/HI net897 sky130_fd_sc_hd__conb_1
XANTENNA__06132__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05667_ top.cb_syn.char_path\[10\] net547 net310 top.cb_syn.char_path\[106\] vssd1
+ vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22o_1
X_08455_ net1238 top.cb_syn.char_path_n\[104\] net240 vssd1 vssd1 vccd1 vccd1 _01587_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout431_A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08386_ net1782 net204 _04755_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout529_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05598_ net1169 net168 _02671_ net210 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a22o_1
X_07406_ _02515_ net126 net123 _04033_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ _03776_ _03783_ _03978_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05891__A1 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ net270 _03936_ _03937_ net276 net1683 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06219_ net482 net534 _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__and3_1
XANTENNA__06840__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ top.findLeastValue.val2\[34\] top.findLeastValue.val1\[34\] vssd1 vssd1 vccd1
+ vccd1 _03875_ sky130_fd_sc_hd__nand2_1
X_09007_ top.histogram.eof_n _03321_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and2_1
XANTENNA__09385__A2 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__B1 _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout541 top.sram_interface.word_cnt\[3\] vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_2
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05946__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__and2_1
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
Xfanout552 net553 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_2
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_1
Xfanout596 net597 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08896__A1 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09424__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net588 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_85_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ clknet_leaf_6_clk _02335_ _01174_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_1_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11733_ clknet_leaf_40_clk _02283_ _01123_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07320__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11664_ clknet_leaf_113_clk _02214_ _01054_ vssd1 vssd1 vccd1 vccd1 top.path\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05882__A1 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ net719 net554 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_94_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09073__A1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11595_ clknet_leaf_0_clk top.dut.bit_buf_next\[2\] _00985_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10546_ net833 net668 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__and2_1
X_10477_ net841 net676 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08584__B1 _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05937__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11029_ clknet_leaf_56_clk net1098 _00419_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06347__C1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06958__B _03609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05862__B _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08887__A1 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05570__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06570_ top.header_synthesis.write_char_path top.header_synthesis.start vssd1 vssd1
+ vccd1 vccd1 _03370_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_86_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05521_ _02563_ _02582_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__nor2_1
X_08240_ net1767 net198 _04682_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05452_ top.WB.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__nand2_1
X_08171_ top.cb_syn.char_path_n\[119\] net371 net329 top.cb_syn.char_path_n\[117\]
+ net175 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a221o_1
XANTENNA__05873__A1 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05383_ top.findLeastValue.histo_index\[8\] vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__inv_2
X_07122_ top.findLeastValue.val2\[12\] top.findLeastValue.val1\[12\] vssd1 vssd1 vccd1
+ vccd1 _03798_ sky130_fd_sc_hd__nor2_1
XANTENNA__06822__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07053_ _03726_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__nor2_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_06004_ _02916_ _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ top.hTree.tree_reg\[6\] top.findLeastValue.sum\[6\] net284 vssd1 vssd1 vccd1
+ vccd1 _04490_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout479_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ top.findLeastValue.val2\[1\] net129 net120 _03658_ vssd1 vssd1 vccd1 vccd1
+ _02009_ sky130_fd_sc_hd__o22a_1
XANTENNA__08878__A1 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ net770 net605 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__and2_1
X_07886_ top.findLeastValue.sum\[20\] _04434_ net391 vssd1 vssd1 vccd1 vccd1 _04435_
+ sky130_fd_sc_hd__mux2_1
X_06837_ top.compVal\[35\] top.findLeastValue.val1\[35\] net152 vssd1 vssd1 vccd1
+ vccd1 _03624_ sky130_fd_sc_hd__mux2_1
X_06768_ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__inv_2
X_09556_ net734 net569 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__and2_1
X_08507_ net1136 top.cb_syn.char_path_n\[52\] net242 vssd1 vssd1 vccd1 vccd1 _01535_
+ sky130_fd_sc_hd__mux2_1
X_09487_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout813_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ _03478_ _03489_ _03490_ _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__or4b_1
XANTENNA__07302__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05719_ net1314 net170 _02772_ net209 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__a22o_1
X_08438_ net1317 top.cb_syn.char_path_n\[121\] net234 vssd1 vssd1 vccd1 vccd1 _01604_
+ sky130_fd_sc_hd__mux2_1
X_08369_ top.cb_syn.char_path_n\[20\] net377 net334 top.cb_syn.char_path_n\[18\] net180
+ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__a221o_1
XANTENNA__09055__A1 top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ clknet_leaf_18_clk _01945_ _00770_ vssd1 vssd1 vccd1 vccd1 top.cw2\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06823__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ net746 net581 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ net728 net563 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09358__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10193_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout371 net374 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
Xfanout382 net386 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_70_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout360 _02593_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
Xfanout393 _04049_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08485__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05552__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11716_ clknet_leaf_69_clk _02266_ _01106_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
X_11647_ clknet_leaf_111_clk _02197_ _01037_ vssd1 vssd1 vccd1 vccd1 top.path\[46\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 gpio_in[10] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
X_11578_ clknet_leaf_5_clk _02143_ _00968_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
Xhold808 top.cb_syn.char_path_n\[112\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 top.cb_syn.char_path_n\[100\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ net805 net640 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__and2_1
XANTENNA__09349__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07564__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ net474 _04317_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__nand2_1
XANTENNA__07780__A1 top.findLeastValue.sum\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07532__A1 top.cb_syn.char_path_n\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ net449 net1160 _04257_ _04261_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__o22a_1
X_09410_ net1580 net229 _05286_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06622_ _02432_ top.findLeastValue.val1\[17\] top.findLeastValue.val1\[16\] _02433_
+ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09341_ net986 net220 net214 _04411_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__a22o_1
X_06553_ net1422 _03327_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nor2_1
X_05504_ net526 _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_51_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06484_ net1498 _03319_ net300 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
X_09272_ net343 _05225_ _04081_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[4\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ top.cb_syn.char_path_n\[93\] net369 net326 top.cb_syn.char_path_n\[91\] net172
+ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a221o_1
X_05435_ top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08154_ top.cb_syn.char_path_n\[127\] net190 _04639_ vssd1 vssd1 vccd1 vccd1 _01746_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_99_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout227_A _05253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05366_ top.findLeastValue.val1\[40\] vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__inv_2
X_08085_ net488 _04178_ _04585_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a211o_1
X_07105_ top.findLeastValue.val2\[20\] top.findLeastValue.val1\[20\] vssd1 vssd1 vccd1
+ vccd1 _03781_ sky130_fd_sc_hd__nand2_1
X_05297_ top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__inv_2
X_07036_ _03708_ _03709_ _03710_ _03711_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_08987_ top.WB.CPU_DAT_O\[14\] top.cb_syn.h_element\[46\] net368 vssd1 vssd1 vccd1
+ vccd1 _01351_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout763_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A1 top.findLeastValue.sum\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06598__B top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ net418 _04475_ _04476_ net261 vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07869_ net431 net1431 net253 top.findLeastValue.sum\[24\] _04421_ vssd1 vssd1 vccd1
+ vccd1 _01813_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10880_ clknet_leaf_23_clk top.header_synthesis.next_header\[2\] _00270_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[2\] sky130_fd_sc_hd__dfrtp_1
X_09608_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__and2_1
X_09539_ net722 net557 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11501_ clknet_leaf_120_clk _02066_ _00891_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11432_ clknet_leaf_95_clk _01997_ _00822_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[36\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ clknet_leaf_91_clk _01928_ _00753_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[41\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10314_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__and2_1
X_11294_ clknet_leaf_22_clk _01859_ _00684_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08988__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net818 net653 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__and2_1
X_10176_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__and2_1
Xfanout190 net192 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05773__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10493__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold605 top.cb_syn.curr_index\[1\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 top.hTree.tree_reg\[16\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09059__B _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold627 top.histogram.total\[0\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 top.hTree.tree_reg\[11\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 top.hTree.tree_reg\[10\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
X_09890_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__and2_1
XANTENNA__08625__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08910_ top.hTree.write_HT_fin net470 _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__and3_1
X_08841_ _02813_ _05023_ _05025_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or4_1
XANTENNA__08950__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05764__B1 _02806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ _02546_ _04959_ _04960_ _02545_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a31o_1
X_05984_ top.WB.CPU_DAT_O\[17\] net1391 net346 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
X_07723_ net472 _04300_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout177_A _04616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07654_ _02831_ _02835_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06605_ top.compVal\[23\] top.compVal\[22\] top.compVal\[21\] top.compVal\[20\] vssd1
+ vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08138__B net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ top.cb_syn.max_index\[6\] top.cb_syn.max_index\[5\] _04184_ vssd1 vssd1 vccd1
+ vccd1 _04185_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ net993 net224 net217 _04479_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06536_ net1596 _03353_ _03334_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__o21ba_1
X_09255_ top.cb_syn.zero_count\[4\] _05214_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__or2_1
X_06467_ net1467 _03308_ net300 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05418_ top.cb_syn.cb_length\[3\] vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout609_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08206_ top.cb_syn.char_path_n\[101\] net201 _04665_ vssd1 vssd1 vccd1 vccd1 _01720_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05778__A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06398_ top.hist_data_o\[28\] top.hist_data_o\[27\] _03262_ vssd1 vssd1 vccd1 vccd1
+ _03263_ sky130_fd_sc_hd__and3_1
X_09186_ net1677 _05051_ net254 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08137_ _02535_ _04627_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05349_ top.findLeastValue.val2\[28\] vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__inv_2
X_08068_ _04566_ _04573_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06244__B2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ top.findLeastValue.val2\[18\] top.findLeastValue.val2\[17\] top.findLeastValue.val2\[16\]
+ top.findLeastValue.val2\[15\] vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__and4_1
XANTENNA__08616__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ net785 net620 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__and2_1
XANTENNA__08941__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ clknet_leaf_59_clk _01497_ _00322_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10863_ clknet_leaf_28_clk top.header_synthesis.next_zero_count\[4\] _00253_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[4\] sky130_fd_sc_hd__dfrtp_1
X_10794_ clknet_leaf_113_clk _01400_ _00184_ vssd1 vssd1 vccd1 vccd1 top.path\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10594__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08224__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ clknet_leaf_78_clk _01980_ _00805_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[19\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_117_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ clknet_leaf_76_clk _01911_ _00736_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05994__A0 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ clknet_leaf_44_clk _01842_ _00667_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_10228_ net810 net645 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__and2_1
XANTENNA__08932__B1 _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10159_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__and2_1
Xhold2 top.HT_fin_reg vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__B net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06710__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07370_ net272 _04010_ _04011_ net278 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1
+ vccd1 _01898_ sky130_fd_sc_hd__a32o_1
X_06321_ _02603_ _03184_ _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a21o_1
XANTENNA__08999__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06252_ _03119_ _03123_ net459 vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__o21a_1
X_09040_ top.WB.CPU_DAT_O\[10\] net1311 net315 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
XANTENNA__07671__B1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08215__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 top.histogram.sram_out\[24\] vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
X_06183_ net545 _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold435 _01548_ vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold413 top.histogram.total\[31\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 top.path\[60\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net794 net629 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__and2_1
Xhold457 top.header_synthesis.header\[0\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 net103 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 top.path\[85\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold479 top.header_synthesis.count\[7\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05985__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__and2_1
X_08824_ top.path\[97\] net325 _05012_ net427 net430 vssd1 vssd1 vccd1 vccd1 _05013_
+ sky130_fd_sc_hd__o221a_1
X_08755_ top.path\[22\] top.path\[23\] net512 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__mux2_1
X_07706_ top.hTree.tree_reg\[55\] _04248_ net387 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05780__B net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05967_ top.sram_interface.TRN_counter\[2\] top.sram_interface.TRN_counter\[1\] top.sram_interface.TRN_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__and3b_1
X_08686_ top.cb_syn.i\[2\] _04879_ _04886_ _04891_ vssd1 vssd1 vccd1 vccd1 _01466_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05898_ top.hist_data_o\[0\] top.WB.CPU_DAT_O\[0\] net349 vssd1 vssd1 vccd1 vccd1
+ _02252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07637_ top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\] top.cb_syn.max_index\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout726_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ _04166_ _04167_ net289 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06519_ net1487 _03340_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__xor2_1
X_09307_ top.header_synthesis.bit1 net36 top.header_synthesis.enable _02807_ vssd1
+ vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_101_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07499_ net342 top.dut.bits_in_buf_next\[0\] _04094_ _04099_ vssd1 vssd1 vccd1 vccd1
+ _04100_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ net1064 _05205_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[7\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ top.cb_syn.setup net488 top.cb_syn.curr_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _05168_ sky130_fd_sc_hd__or3b_1
XANTENNA__05301__A top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11200_ clknet_leaf_30_clk _01765_ _00590_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06831__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ clknet_leaf_60_clk _01696_ _00521_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07965__A1 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05976__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ clknet_leaf_61_clk _01627_ _00452_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_10013_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__and2_1
XANTENNA__08758__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold840_A top.findLeastValue.sum\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06940__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ clknet_leaf_5_clk net918 _00305_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11895_ net926 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
X_10846_ clknet_leaf_2_clk _01440_ _00236_ vssd1 vssd1 vccd1 vccd1 top.translation.totalEn
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06456__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ clknet_leaf_113_clk _01383_ _00167_ vssd1 vssd1 vccd1 vccd1 top.path\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07405__A0 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07248__B1_N net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ clknet_leaf_88_clk _01894_ _00719_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07708__A1 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_105_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11883__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ top.findLeastValue.val2\[19\] net128 net117 _03640_ vssd1 vssd1 vccd1 vccd1
+ _02027_ sky130_fd_sc_hd__o22a_1
XANTENNA__07572__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05821_ top.findLeastValue.least2\[8\] top.findLeastValue.least1\[8\] _02842_ vssd1
+ vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or3b_1
X_08540_ net1228 top.cb_syn.char_path_n\[19\] net246 vssd1 vssd1 vccd1 vccd1 _01502_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09072__B _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05752_ net442 _02793_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__or2_1
X_08471_ net1186 top.cb_syn.char_path_n\[88\] net236 vssd1 vssd1 vccd1 vccd1 _01571_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07567__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05683_ net1397 net169 _02742_ net211 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09800__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ top.findLeastValue.least1\[6\] net141 _03660_ net482 vssd1 vssd1 vccd1 vccd1
+ _01875_ sky130_fd_sc_hd__a22o_1
XANTENNA__05498__A2 _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07353_ _03798_ _03852_ _03797_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06304_ top.cb_syn.char_index\[2\] top.cb_syn.char_index\[1\] _02588_ net309 vssd1
+ vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__o22a_1
X_07284_ net270 _03948_ _03949_ net276 top.findLeastValue.sum\[35\] vssd1 vssd1 vccd1
+ vccd1 _01922_ sky130_fd_sc_hd__a32o_1
XANTENNA__06998__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06235_ top.TRN_char_index\[4\] _03050_ top.TRN_char_index\[5\] vssd1 vssd1 vccd1
+ vccd1 _03108_ sky130_fd_sc_hd__a21oi_1
X_09023_ top.WB.CPU_DAT_O\[27\] net1223 net314 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
Xhold210 top.cb_syn.char_path\[116\] vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05670__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06166_ top.cb_syn.char_index\[6\] top.cb_syn.char_index\[5\] _02607_ _03035_ _03040_
+ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__a41o_1
Xhold221 top.path\[57\] vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 top.path\[103\] vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 top.path\[121\] vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08151__B net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06097_ net523 net463 _02969_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__and3_2
Xhold287 top.cb_syn.char_path\[104\] vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 top.cb_syn.char_path\[102\] vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 top.path\[55\] vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 top.path\[119\] vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__and2_1
Xfanout701 net702 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_2
Xhold298 top.hTree.nulls\[60\] vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 net44 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_4
Xfanout723 net726 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_2
X_11939__902 vssd1 vssd1 vccd1 vccd1 _11939__902/HI net902 sky130_fd_sc_hd__conb_1
X_09856_ net871 net706 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__and2_1
Xfanout767 net768 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_2
Xfanout745 net748 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_2
Xfanout734 net735 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_2
Xfanout789 net794 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_2
Xfanout778 net780 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_2
X_08807_ net427 _04994_ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__o21a_1
X_09787_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout843_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ _02511_ net126 net123 _03684_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06922__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ top.path\[126\] top.path\[127\] net511 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__mux2_1
X_08669_ _04605_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__or2_2
XANTENNA__06135__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10700_ clknet_leaf_7_clk _01331_ _00090_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11680_ clknet_leaf_94_clk _02230_ _01070_ vssd1 vssd1 vccd1 vccd1 top.compVal\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_10631_ clknet_leaf_66_clk _01262_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ net860 net695 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__and2_1
XANTENNA__06127__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05661__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ net753 net588 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07938__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05949__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ clknet_leaf_38_clk _01679_ _00504_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_11045_ clknet_leaf_39_clk _01610_ _00435_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_11947_ net910 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__06126__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11878_ net881 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__07421__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10829_ clknet_leaf_97_clk _01423_ _00219_ vssd1 vssd1 vccd1 vccd1 top.path\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09379__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06020_ top.sram_interface.init_counter\[9\] _02931_ vssd1 vssd1 vccd1 vccd1 _02932_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__05652__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ top.findLeastValue.sum\[3\] _04502_ net391 vssd1 vssd1 vccd1 vccd1 _04503_
+ sky130_fd_sc_hd__mux2_1
X_09710_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__and2_1
X_06922_ top.findLeastValue.val1\[35\] net137 net114 top.compVal\[35\] vssd1 vssd1
+ vccd1 vccd1 _01996_ sky130_fd_sc_hd__o22a_1
X_09641_ net762 net597 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__and2_1
X_06853_ top.compVal\[27\] top.findLeastValue.val1\[27\] net151 vssd1 vssd1 vccd1
+ vccd1 _03632_ sky130_fd_sc_hd__mux2_1
X_09572_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__and2_1
XANTENNA__06904__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06784_ top.compVal\[28\] _02466_ _03566_ _03574_ vssd1 vssd1 vccd1 vccd1 _03582_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10022__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05804_ top.sram_interface.write_counter_FLV\[0\] net455 _02823_ vssd1 vssd1 vccd1
+ vccd1 _02828_ sky130_fd_sc_hd__nand3_1
X_08523_ net1141 top.cb_syn.char_path_n\[36\] net237 vssd1 vssd1 vccd1 vccd1 _01519_
+ sky130_fd_sc_hd__mux2_1
X_05735_ top.TRN_char_index\[3\] net41 net715 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
X_05666_ top.cb_syn.char_path\[74\] net540 net529 top.cb_syn.char_path\[42\] vssd1
+ vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
X_08454_ net1115 top.cb_syn.char_path_n\[105\] net240 vssd1 vssd1 vccd1 vccd1 _01588_
+ sky130_fd_sc_hd__mux2_1
X_08385_ top.cb_syn.char_path_n\[12\] net383 net340 top.cb_syn.char_path_n\[10\] net187
+ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a221o_1
X_05597_ top.hTree.node_reg\[22\] net410 _02669_ _02670_ vssd1 vssd1 vccd1 vccd1 _02671_
+ sky130_fd_sc_hd__a211o_1
X_07405_ net482 top.findLeastValue.least1\[6\] net150 vssd1 vssd1 vccd1 vccd1 _04033_
+ sky130_fd_sc_hd__mux2_1
X_07336_ net269 _03986_ _03987_ net275 net1680 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a32o_1
XANTENNA__08814__C1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09006_ top.WB.CPU_DAT_O\[14\] net1270 net365 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
X_07267_ _03721_ _03935_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout793_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06218_ net483 net484 _03089_ _02787_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a31o_1
X_07198_ _03872_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__and2_1
X_06149_ top.sram_interface.init_counter\[10\] _03025_ _03018_ vssd1 vssd1 vccd1 vccd1
+ _03026_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08593__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 top.cb_syn.char_path_n\[0\] vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_2
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
X_09908_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__and2_1
XANTENNA__08345__A1 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout553 net571 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_2
Xfanout575 net584 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_2
Xfanout564 net571 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_2
X_09839_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__and2_1
Xfanout597 net612 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_2
Xfanout586 net588 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11801_ clknet_leaf_7_clk _02334_ _01173_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_57_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ clknet_leaf_40_clk _02282_ _01122_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11663_ clknet_leaf_113_clk _02213_ _01053_ vssd1 vssd1 vccd1 vccd1 top.path\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10614_ net719 net554 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ clknet_leaf_5_clk top.dut.bit_buf_next\[1\] _00984_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ net736 net571 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__and2_1
X_10476_ net856 net691 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08584__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ clknet_leaf_57_clk _01593_ _00418_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06958__C net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07850__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05520_ net461 net545 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__nand2_1
X_05451_ top.WB.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__and2_1
X_08170_ net1738 net195 _04647_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__o21a_1
XANTENNA_16 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05382_ top.findLeastValue.wipe_the_char_2 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07121_ top.findLeastValue.val2\[12\] top.findLeastValue.val1\[12\] vssd1 vssd1 vccd1
+ vccd1 _03797_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
X_07052_ top.findLeastValue.val2\[37\] top.findLeastValue.val1\[37\] vssd1 vssd1 vccd1
+ vccd1 _03728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06003_ net542 net452 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nand2_1
X_07954_ net436 net1603 net249 net1800 _04489_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a221o_1
X_07885_ top.hTree.tree_reg\[20\] top.findLeastValue.sum\[20\] net283 vssd1 vssd1
+ vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
X_06905_ top.compVal\[1\] top.findLeastValue.val1\[1\] net154 vssd1 vssd1 vccd1 vccd1
+ _03658_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout374_A _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ net770 net605 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__and2_1
X_06836_ top.findLeastValue.val2\[36\] net128 net118 _03623_ vssd1 vssd1 vccd1 vccd1
+ _02044_ sky130_fd_sc_hd__o22a_1
XANTENNA__07760__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A top.sram_interface.word_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06767_ top.compVal\[29\] _02465_ _02466_ top.compVal\[28\] vssd1 vssd1 vccd1 vccd1
+ _03565_ sky130_fd_sc_hd__a22o_1
X_09555_ net734 net569 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__and2_1
X_08506_ net1071 top.cb_syn.char_path_n\[53\] net232 vssd1 vssd1 vccd1 vccd1 _01536_
+ sky130_fd_sc_hd__mux2_1
X_09486_ net765 net600 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05718_ top.histogram.sram_out\[2\] net357 net408 top.hTree.node_reg\[2\] _02771_
+ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__a221o_1
X_06698_ _02413_ top.findLeastValue.val1\[34\] _02489_ top.compVal\[32\] _03480_ vssd1
+ vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__o221a_1
X_05649_ _02712_ _02713_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ net1280 top.cb_syn.char_path_n\[122\] net234 vssd1 vssd1 vccd1 vccd1 _01605_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout806_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ top.cb_syn.char_path_n\[20\] net198 _04746_ vssd1 vssd1 vccd1 vccd1 _01639_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08299_ top.cb_syn.char_path_n\[55\] net372 net329 top.cb_syn.char_path_n\[53\] net175
+ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a221o_1
X_07319_ _03866_ _03973_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nand2_1
XANTENNA__08802__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05616__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08566__A1 _02538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__and2_1
Xfanout350 net352 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout383 net385 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_2
Xfanout372 net374 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06329__B1 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout361 _02578_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_2
Xfanout394 net397 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_4
XFILLER_0_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ clknet_leaf_69_clk _02265_ _01105_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11646_ clknet_leaf_108_clk _02196_ _01036_ vssd1 vssd1 vccd1 vccd1 top.path\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_11577_ clknet_leaf_27_clk _02142_ _00967_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_103_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput36 gpio_in[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xhold809 top.hist_data_o\[20\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
X_10528_ net804 net639 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__and2_1
XANTENNA__08557__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ net735 net570 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__and2_1
XANTENNA__07845__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07670_ _04259_ _04260_ net474 vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__mux2_1
XANTENNA__05543__A1 top.hTree.node_reg\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ _03415_ _03416_ _03417_ _03418_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__or4b_1
X_09340_ net983 net221 net219 _04415_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__a22o_1
X_06552_ _03329_ _03359_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05503_ net537 net528 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_51_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ _04044_ _04095_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__nor2_1
X_08222_ top.cb_syn.char_path_n\[93\] net191 _04673_ vssd1 vssd1 vccd1 vccd1 _01712_
+ sky130_fd_sc_hd__o21a_1
X_06483_ top.hist_data_o\[2\] _03245_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05434_ net550 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__inv_2
XANTENNA__08245__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ top.cb_syn.curr_path\[127\] net369 net326 top.cb_syn.char_path_n\[126\] net172
+ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_99_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05365_ top.findLeastValue.val1\[41\] vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08084_ top.cb_syn.check_right _04552_ _02896_ net412 vssd1 vssd1 vccd1 vccd1 _04586_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06256__C1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ _03778_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08796__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05296_ top.compVal\[34\] vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__inv_2
X_07035_ top.findLeastValue.val1\[34\] top.findLeastValue.val1\[33\] top.findLeastValue.val1\[32\]
+ top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07755__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ top.WB.CPU_DAT_O\[15\] top.cb_syn.h_element\[47\] net368 vssd1 vssd1 vccd1
+ vccd1 _01352_ sky130_fd_sc_hd__mux2_1
X_07937_ net477 _04474_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07868_ net422 _04419_ _04420_ net259 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o211a_1
X_07799_ net435 net1607 net252 top.findLeastValue.sum\[38\] _04365_ vssd1 vssd1 vccd1
+ vccd1 _01827_ sky130_fd_sc_hd__a221o_1
X_09607_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__and2_1
X_06819_ top.compVal\[44\] top.findLeastValue.val1\[44\] net153 vssd1 vssd1 vccd1
+ vccd1 _03615_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09538_ net737 net572 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__and2_1
X_09469_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__and2_1
X_11500_ clknet_leaf_120_clk _02065_ _00890_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ clknet_leaf_96_clk _01996_ _00821_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[35\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_59_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11362_ clknet_leaf_81_clk _01927_ _00752_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_10313_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__and2_1
X_11293_ clknet_leaf_24_clk _01858_ _00683_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10244_ net817 net652 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__and2_1
X_10175_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__and2_1
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
Xfanout180 net189 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
XANTENNA__05773__B2 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11629_ clknet_leaf_28_clk _02179_ _01019_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08778__B2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 _01805_ vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold606 top.hTree.tree_reg\[22\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold639 _01799_ vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold628 top.hTree.tree_reg\[5\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08625__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08840_ net513 top.translation.totalEn net466 _05028_ vssd1 vssd1 vccd1 vccd1 _05029_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06961__B1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05764__B2 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08771_ _04948_ _04949_ _04950_ net429 net502 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a221o_1
X_05983_ top.WB.CPU_DAT_O\[18\] net1117 net346 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ net472 _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__nand2_1
X_07653_ net1556 _04246_ _04212_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__mux2_1
X_06604_ top.compVal\[31\] top.compVal\[30\] top.compVal\[29\] top.compVal\[28\] vssd1
+ vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09323_ net1003 net226 net217 _04483_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__a22o_1
X_07584_ top.cb_syn.max_index\[4\] _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__or2_1
X_06535_ top.histogram.total\[15\] top.histogram.total\[14\] _03333_ vssd1 vssd1 vccd1
+ vccd1 _03353_ sky130_fd_sc_hd__and3_1
X_09254_ top.cb_syn.zero_count\[4\] _05214_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nand2_1
X_06466_ _03250_ _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05417_ top.cb_syn.cb_length\[4\] vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__inv_2
X_08205_ top.cb_syn.char_path_n\[102\] net380 net336 top.cb_syn.char_path_n\[100\]
+ net183 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ top.hTree.state\[4\] net255 _05121_ net1522 vssd1 vssd1 vccd1 vccd1 _00023_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__05778__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _04617_ _04619_ net190 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__o21a_1
X_06397_ top.hist_data_o\[26\] _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08769__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05348_ top.findLeastValue.val2\[29\] vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__inv_2
X_08067_ top.cb_syn.zeroes\[7\] _04575_ _04576_ _04577_ vssd1 vssd1 vccd1 vccd1 _01771_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07018_ top.findLeastValue.val2\[22\] top.findLeastValue.val2\[21\] top.findLeastValue.val2\[20\]
+ top.findLeastValue.val2\[19\] vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__and4_1
XANTENNA__08616__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A1 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net465 top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__nand2_1
XANTENNA__06829__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ clknet_leaf_59_clk _01496_ _00321_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05733__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10862_ clknet_leaf_29_clk top.header_synthesis.next_zero_count\[3\] _00252_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[3\] sky130_fd_sc_hd__dfrtp_1
X_10793_ clknet_leaf_113_clk _01399_ _00183_ vssd1 vssd1 vccd1 vccd1 top.path\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05969__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05691__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ clknet_leaf_79_clk _01979_ _00804_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[18\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11345_ clknet_leaf_76_clk _01910_ _00735_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11276_ clknet_leaf_43_clk _01841_ _00666_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08607__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ net812 net647 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 top.cb_syn.finished vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
X_10158_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__and2_1
XANTENNA__06943__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ net832 net667 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__and2_1
X_11891__922 vssd1 vssd1 vccd1 vccd1 net922 _11891__922/LO sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06320_ top.findLeastValue.histo_index\[2\] net361 _02600_ _03188_ _03187_ vssd1
+ vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__a221o_1
X_06251_ net483 net361 _03122_ net534 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a22o_1
XANTENNA__05682__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07671__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06182_ top.TRN_char_index\[5\] top.TRN_char_index\[4\] _03055_ vssd1 vssd1 vccd1
+ vccd1 _03057_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold436 top.cb_syn.char_path\[59\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 top.cb_syn.char_path\[34\] vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 net83 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 top.histogram.sram_out\[6\] vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ net788 net623 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold458 top.cb_syn.char_path\[2\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 top.cb_syn.char_path\[5\] vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 top.path\[78\] vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
X_09872_ net790 net625 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__and2_1
XANTENNA__05737__A1 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06934__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08823_ top.path\[98\] top.path\[99\] net510 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__mux2_1
X_05966_ _02902_ _02912_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout287_A _03394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08754_ top.path\[28\] net405 _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__o21a_1
X_07705_ net257 _04288_ _04289_ net1191 net432 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a32o_1
XANTENNA__08149__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ top.cb_syn.i\[2\] _04880_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_49_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_92_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout454_A top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05897_ top.hist_data_o\[1\] top.WB.CPU_DAT_O\[1\] net349 vssd1 vssd1 vccd1 vccd1
+ _02253_ sky130_fd_sc_hd__mux2_1
X_07636_ net518 top.cb_syn.h_element\[48\] net525 top.cb_syn.h_element\[57\] _04180_
+ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__a221o_1
X_07567_ top.cb_syn.char_path_n\[58\] top.cb_syn.char_path_n\[57\] top.cb_syn.char_path_n\[60\]
+ top.cb_syn.char_path_n\[59\] net394 net292 vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout621_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06518_ _03341_ net1507 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__nor2_1
X_09306_ net513 _05249_ net423 vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout719_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09237_ top.header_synthesis.header\[7\] top.cb_syn.char_index\[7\] net490 vssd1
+ vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07498_ top.dut.bits_in_buf_next\[1\] _04091_ _04095_ _04098_ _04046_ vssd1 vssd1
+ vccd1 vccd1 _04099_ sky130_fd_sc_hd__a221o_1
X_06449_ net1013 net298 vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__nand2_1
XANTENNA__05673__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ net519 _05165_ _05166_ _05167_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a211o_1
XANTENNA__09403__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ _04178_ net370 vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nor2_1
X_09099_ net462 net534 _02582_ _03038_ _02575_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a32o_1
X_11130_ clknet_leaf_59_clk _01695_ _00520_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[76\]
+ sky130_fd_sc_hd__dfrtp_2
X_11061_ clknet_leaf_56_clk _01626_ _00451_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10012_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__and2_1
XANTENNA__06925__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__B net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
X_11894_ net925 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
X_11916__947 vssd1 vssd1 vccd1 vccd1 net947 _11916__947/LO sky130_fd_sc_hd__conb_1
X_10914_ clknet_leaf_4_clk net952 _00304_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10845_ clknet_leaf_108_clk _01439_ _00235_ vssd1 vssd1 vccd1 vccd1 top.path\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10776_ clknet_leaf_109_clk _01382_ _00166_ vssd1 vssd1 vccd1 vccd1 top.path\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__B1 top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05664__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06208__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11328_ clknet_leaf_88_clk _01893_ _00718_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11259_ clknet_leaf_80_clk _01824_ _00649_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07708__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05820_ top.sram_interface.counter_HTREE\[0\] _02841_ top.sram_interface.counter_HTREE\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_74_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
X_05751_ net444 _02562_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__nor2_1
X_08470_ net1554 net1808 net234 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__mux2_1
XANTENNA__07567__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05682_ top.histogram.sram_out\[8\] net358 net409 top.hTree.node_reg\[8\] _02741_
+ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07421_ net287 _04040_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07352_ net269 _03977_ _03998_ net275 net1707 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06303_ _03019_ _03171_ _03172_ top.histogram.init net454 vssd1 vssd1 vccd1 vccd1
+ _03173_ sky130_fd_sc_hd__o221a_1
XANTENNA__09094__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07283_ _03880_ _03947_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__nand2_1
XANTENNA__05655__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06234_ top.TRN_char_index\[5\] _03056_ _03106_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o21a_1
X_09022_ top.WB.CPU_DAT_O\[28\] net1372 net313 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
Xhold200 top.cb_syn.char_path\[55\] vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06165_ _02787_ _03037_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a21oi_1
Xhold211 top.path\[16\] vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold233 top.cb_syn.char_path\[83\] vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 top.header_synthesis.header\[3\] vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 top.hTree.tree_reg\[59\] vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 top.cb_syn.char_path\[19\] vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
X_06096_ _02554_ net423 _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__or3_4
Xhold255 top.hTree.nulls\[62\] vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09149__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05958__B2 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold266 top.path\[76\] vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__and2_1
Xfanout702 net711 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_2
Xhold299 top.path\[67\] vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_2
Xhold288 top.path\[0\] vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout713 net714 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08357__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__and2_1
Xfanout746 net747 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09544__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_2
Xfanout757 net796 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout768 net771 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_2
Xfanout779 net780 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout571_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ top.path\[44\] net404 net324 top.path\[45\] net505 vssd1 vssd1 vccd1 vccd1
+ _04995_ sky130_fd_sc_hd__o221a_1
X_09786_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__and2_1
XANTENNA__09158__A_N top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06998_ top.cw1\[1\] net148 _03662_ net487 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_65_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout836_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ top.path\[52\] top.path\[53\] top.path\[54\] top.path\[55\] net511 net507
+ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__mux4_1
X_05949_ top.compVal\[12\] net161 net146 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 _02229_ sky130_fd_sc_hd__a22o_1
X_08668_ net522 net523 _04189_ _04190_ _04561_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o221ai_2
X_07619_ net521 _04214_ _04217_ net516 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__a22o_1
X_08599_ top.cb_syn.char_path_n\[121\] top.cb_syn.char_path_n\[122\] top.cb_syn.char_path_n\[125\]
+ top.cb_syn.char_path_n\[126\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__mux4_1
X_10630_ clknet_leaf_67_clk _01261_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10561_ net862 net697 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__and2_1
XANTENNA__08832__B1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10492_ net780 net615 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07399__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05949__B2 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ clknet_leaf_37_clk _01678_ _00503_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ clknet_leaf_39_clk _01609_ _00434_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08363__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
X_11946_ net909 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__07874__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ net880 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828_ clknet_leaf_96_clk _01422_ _00218_ vssd1 vssd1 vccd1 vccd1 top.path\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ clknet_leaf_8_clk net1041 _00149_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05637__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ top.hTree.tree_reg\[3\] top.findLeastValue.sum\[3\] net284 vssd1 vssd1 vccd1
+ vccd1 _04502_ sky130_fd_sc_hd__mux2_1
XANTENNA__09000__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ top.findLeastValue.val1\[36\] net137 net114 top.compVal\[36\] vssd1 vssd1
+ vccd1 vccd1 _01997_ sky130_fd_sc_hd__o22a_1
XANTENNA__08354__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ net760 net595 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__and2_1
X_06852_ top.findLeastValue.val2\[28\] net127 net118 _03631_ vssd1 vssd1 vccd1 vccd1
+ _02036_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09571_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__and2_1
X_06783_ top.compVal\[20\] top.findLeastValue.val2\[20\] vssd1 vssd1 vccd1 vccd1 _03581_
+ sky130_fd_sc_hd__xnor2_1
X_05803_ net1631 _02824_ _02825_ _02827_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a22o_1
XANTENNA__10022__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
X_08522_ net1271 top.cb_syn.char_path_n\[37\] net239 vssd1 vssd1 vccd1 vccd1 _01520_
+ sky130_fd_sc_hd__mux2_1
X_05734_ top.TRN_char_index\[4\] net42 net715 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XANTENNA__08737__S0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ net1358 top.cb_syn.char_path_n\[106\] net241 vssd1 vssd1 vccd1 vccd1 _01589_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07314__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09303__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05665_ net1307 net168 _02727_ net210 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a22o_1
X_07404_ top.findLeastValue.least2\[7\] net127 net117 _04032_ vssd1 vssd1 vccd1 vccd1
+ _01885_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout152_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08384_ top.cb_syn.char_path_n\[12\] net204 _04754_ vssd1 vssd1 vccd1 vccd1 _01631_
+ sky130_fd_sc_hd__o21a_1
X_05596_ top.histogram.sram_out\[22\] net359 net354 top.hTree.node_reg\[54\] vssd1
+ vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
X_07335_ _03780_ _03985_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09539__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ _03721_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout417_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ top.WB.CPU_DAT_O\[15\] net1331 net366 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
X_06217_ net484 _03089_ _02787_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__a21oi_1
X_07197_ _03855_ _03858_ _03863_ _03870_ _03750_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06840__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06148_ top.sram_interface.init_counter\[9\] _03024_ vssd1 vssd1 vccd1 vccd1 _03025_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06079_ _02977_ _02978_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout786_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__and2_1
Xfanout521 top.cb_syn.curr_state\[4\] vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_2
Xfanout532 top.sram_interface.word_cnt\[10\] vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout510 net512 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08345__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_1
Xfanout565 net567 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_2
Xfanout554 net571 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_2
X_09838_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__and2_1
XANTENNA__06356__A1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout598 net601 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_2
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_2
Xfanout576 net584 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_2
X_09769_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
X_11800_ clknet_leaf_6_clk _02333_ _01172_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__A _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold629_A top.hTree.node_reg\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ clknet_leaf_40_clk _02281_ _01121_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11662_ clknet_leaf_114_clk _02212_ _01052_ vssd1 vssd1 vccd1 vccd1 top.path\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_11593_ clknet_leaf_0_clk top.dut.bit_buf_next\[0\] _00983_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[0\] sky130_fd_sc_hd__dfrtp_1
X_10613_ net719 net554 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__and2_1
XANTENNA__05619__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__S _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ net728 net563 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10475_ net855 net690 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ clknet_leaf_60_clk _01592_ _00417_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06898__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05570__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929_ net892 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_86_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09049__A0 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05450_ net1 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__inv_2
XANTENNA_28 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05381_ top.findLeastValue.val1\[5\] vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ _03790_ _03791_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06822__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07051_ top.findLeastValue.val2\[37\] top.findLeastValue.val1\[37\] vssd1 vssd1 vccd1
+ vccd1 _03727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06002_ net439 _02913_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__nand2_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07953_ net418 _04487_ _04488_ net261 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__o211a_1
X_07884_ net438 net1552 net248 top.findLeastValue.sum\[21\] _04433_ vssd1 vssd1 vccd1
+ vccd1 _01810_ sky130_fd_sc_hd__a221o_1
XANTENNA__06338__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ top.findLeastValue.val2\[2\] net129 net120 _03657_ vssd1 vssd1 vccd1 vccd1
+ _02010_ sky130_fd_sc_hd__o22a_1
X_09623_ net769 net604 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__and2_1
XANTENNA__09822__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06835_ top.compVal\[36\] top.findLeastValue.val1\[36\] net152 vssd1 vssd1 vccd1
+ vccd1 _03623_ sky130_fd_sc_hd__mux2_1
XANTENNA__05561__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ net729 net564 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__and2_1
X_06766_ top.findLeastValue.val2\[21\] top.compVal\[21\] vssd1 vssd1 vccd1 vccd1 _03564_
+ sky130_fd_sc_hd__nand2b_1
X_08505_ net1221 top.cb_syn.char_path_n\[54\] net232 vssd1 vssd1 vccd1 vccd1 _01537_
+ sky130_fd_sc_hd__mux2_1
X_09485_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout534_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07838__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05717_ top.hTree.node_reg\[34\] net307 _02770_ net469 vssd1 vssd1 vccd1 vccd1 _02771_
+ sky130_fd_sc_hd__a22o_1
X_06697_ _03477_ _03482_ _03493_ _03494_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__or4_1
X_08436_ net1333 top.cb_syn.char_path_n\[123\] net234 vssd1 vssd1 vccd1 vccd1 _01606_
+ sky130_fd_sc_hd__mux2_1
X_05648_ top.cb_syn.char_path\[45\] net531 net310 top.cb_syn.char_path\[109\] vssd1
+ vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08367_ top.cb_syn.char_path_n\[21\] net377 net330 top.cb_syn.char_path_n\[19\] net180
+ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout701_A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05579_ top.hTree.node_reg\[25\] net410 _02654_ _02655_ vssd1 vssd1 vccd1 vccd1 _02656_
+ sky130_fd_sc_hd__a211o_1
X_07318_ _03866_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__or2_1
XANTENNA__05797__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ top.cb_syn.char_path_n\[55\] net193 _04711_ vssd1 vssd1 vccd1 vccd1 _01674_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06813__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ _03918_ _03923_ top.findLeastValue.sum\[44\] net277 vssd1 vssd1 vccd1 vccd1
+ _01931_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09716__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05736__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__and2_1
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_2
XANTENNA__05963__C _02898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_2
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_4
XANTENNA__07951__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05552__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11714_ clknet_leaf_69_clk _02264_ _01104_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11645_ clknet_leaf_109_clk _02195_ _01035_ vssd1 vssd1 vccd1 vccd1 top.path\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_11576_ clknet_leaf_27_clk _02141_ _00966_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
Xinput37 gpio_in[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_10527_ net804 net639 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__and2_1
XANTENNA__09907__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ net735 net570 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__and2_1
X_10389_ net770 net605 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__and2_1
X_11924__887 vssd1 vssd1 vccd1 vccd1 _11924__887/HI net887 sky130_fd_sc_hd__conb_1
XANTENNA__07517__A0 top.cb_syn.char_path_n\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07861__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06620_ top.compVal\[19\] top.findLeastValue.val1\[19\] vssd1 vssd1 vccd1 vccd1 _03418_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__05543__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ _03325_ _03328_ net1583 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05502_ net537 net527 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__nor2_1
X_06482_ net1346 net297 _03317_ _03318_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a22o_1
X_09270_ _04046_ _04086_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[3\] sky130_fd_sc_hd__and2_1
X_08221_ top.cb_syn.char_path_n\[94\] net370 net326 top.cb_syn.char_path_n\[92\] net172
+ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a221o_1
X_05433_ net513 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__inv_2
X_08152_ net1555 net172 _04638_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_99_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05364_ top.findLeastValue.val1\[42\] vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08083_ _04203_ _04551_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_9_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
X_07103_ top.findLeastValue.val2\[21\] top.findLeastValue.val1\[21\] vssd1 vssd1 vccd1
+ vccd1 _03779_ sky130_fd_sc_hd__nor2_1
X_05295_ top.compVal\[35\] vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout115_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ top.findLeastValue.val1\[38\] top.findLeastValue.val1\[37\] top.findLeastValue.val1\[36\]
+ top.findLeastValue.val1\[35\] vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__and4_1
XANTENNA__08721__A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ top.WB.CPU_DAT_O\[16\] top.cb_syn.h_element\[48\] net367 vssd1 vssd1 vccd1
+ vccd1 _01353_ sky130_fd_sc_hd__mux2_1
X_07936_ top.hTree.tree_reg\[10\] top.findLeastValue.sum\[10\] net266 vssd1 vssd1
+ vccd1 vccd1 _04475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07771__S _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ net471 _04418_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout651_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07798_ net421 _04363_ _04364_ net260 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__o211a_1
X_09606_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__and2_1
X_06818_ top.findLeastValue.val2\[45\] net131 net119 _03614_ vssd1 vssd1 vccd1 vccd1
+ _02053_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09537_ net744 net579 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__and2_1
XANTENNA__06731__B2 top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06749_ _03531_ _03546_ _03544_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__a21o_1
X_09468_ net840 net675 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__and2_1
X_08419_ top.cb_syn.h_element\[60\] top.cb_syn.h_element\[51\] net518 vssd1 vssd1
+ vccd1 vccd1 _04775_ sky130_fd_sc_hd__mux2_1
X_09399_ top.hTree.nulls\[59\] net400 net228 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o21a_1
X_11430_ clknet_leaf_96_clk _01995_ _00820_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_11361_ clknet_leaf_94_clk _01926_ _00751_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[39\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07946__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ net785 net620 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ clknet_leaf_24_clk _01857_ _00682_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10243_ net818 net653 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__and2_1
XANTENNA__05470__B2 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__and2_1
Xfanout192 _04615_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
Xfanout181 net189 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
XANTENNA__05773__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ clknet_leaf_28_clk _02178_ _01018_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ clknet_leaf_21_clk _02124_ _00949_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
Xhold618 top.hTree.tree_reg\[42\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07856__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 top.hTree.tree_reg\[27\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07986__A0 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold629 top.hTree.node_reg\[63\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05461__B2 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06961__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ _02547_ _04953_ _04956_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__or3_1
X_05982_ top.WB.CPU_DAT_O\[19\] net1189 net346 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
X_07721_ _02515_ net387 _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07604__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ net521 _04243_ _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__a21o_1
X_07583_ top.cb_syn.max_index\[3\] top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_36_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06603_ top.compVal\[27\] top.compVal\[26\] top.compVal\[25\] top.compVal\[24\] vssd1
+ vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09322_ net996 net224 net216 _04487_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__a22o_1
X_06534_ net1563 _03334_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__xor2_1
X_09253_ _05207_ _05213_ _05215_ _05208_ net1561 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[3\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout232_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06465_ top.hist_data_o\[8\] _03249_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__nor2_1
X_05416_ top.cb_syn.zeroes\[0\] vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__inv_2
X_08204_ top.cb_syn.char_path_n\[102\] net201 _04664_ vssd1 vssd1 vccd1 vccd1 _01721_
+ sky130_fd_sc_hd__o21a_1
X_06396_ top.hist_data_o\[25\] top.hist_data_o\[24\] _03260_ vssd1 vssd1 vccd1 vccd1
+ _03261_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05778__C net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09184_ net1004 net254 _05175_ net470 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a22o_1
X_08135_ _02534_ _04626_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__xnor2_1
X_05347_ top.findLeastValue.val2\[33\] vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07766__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08066_ top.cb_syn.zeroes\[7\] _04574_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09547__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ top.findLeastValue.val2\[30\] top.findLeastValue.val2\[29\] top.findLeastValue.val2\[28\]
+ top.findLeastValue.val2\[27\] vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__and4_1
X_08968_ top.WB.CPU_DAT_O\[0\] net1401 net320 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__mux2_1
X_07919_ net437 net1584 net251 top.findLeastValue.sum\[14\] _04461_ vssd1 vssd1 vccd1
+ vccd1 _01803_ sky130_fd_sc_hd__a221o_1
X_08899_ net1054 top.WB.CPU_DAT_O\[3\] net305 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__mux2_1
X_10930_ clknet_leaf_60_clk _01495_ _00320_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10861_ clknet_leaf_29_clk top.header_synthesis.next_zero_count\[2\] _00251_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10792_ clknet_leaf_114_clk _01398_ _00182_ vssd1 vssd1 vccd1 vccd1 top.path\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06845__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05969__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08209__B2 top.cb_syn.char_path_n\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ clknet_leaf_101_clk _01978_ _00803_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[17\]
+ sky130_fd_sc_hd__dfstp_2
X_11344_ clknet_leaf_76_clk _01909_ _00734_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11275_ clknet_leaf_42_clk _01840_ _00665_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10226_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__and2_1
XANTENNA__09904__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__and2_1
Xhold4 top.controller.fin_FLV vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10088_ net824 net659 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__and2_1
X_06250_ _02502_ _03091_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06181_ top.TRN_char_index\[4\] _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 _01517_ vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 top.histogram.sram_out\[11\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 top.path\[65\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09940_ net788 net623 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__and2_1
Xhold437 top.hist_data_o\[23\] vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 top.histogram.sram_out\[1\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 top.path\[63\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__and2_1
X_08822_ net427 _05009_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__o21a_1
X_05965_ _02899_ _02910_ top.CB_write_complete vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a21oi_1
X_08753_ top.path\[29\] net325 _04941_ net427 net502 vssd1 vssd1 vccd1 vccd1 _04942_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__08136__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ net473 _04286_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08684_ _04882_ _04886_ _04890_ _04879_ net1714 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_49_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05896_ top.hist_data_o\[2\] top.WB.CPU_DAT_O\[2\] net349 vssd1 vssd1 vccd1 vccd1
+ _02254_ sky130_fd_sc_hd__mux2_1
X_07635_ top.cb_syn.h_element\[57\] top.cb_syn.h_element\[48\] _04176_ vssd1 vssd1
+ vccd1 vccd1 _04231_ sky130_fd_sc_hd__mux2_1
X_07566_ top.cb_syn.char_path_n\[62\] top.cb_syn.char_path_n\[61\] top.cb_syn.char_path_n\[64\]
+ top.cb_syn.char_path_n\[63\] net394 net292 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06517_ top.histogram.total\[26\] _03340_ net1506 vssd1 vssd1 vccd1 vccd1 _03346_
+ sky130_fd_sc_hd__a21oi_1
X_09305_ top.translation.totalEn _05248_ _05227_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ net1247 _05204_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[6\]
+ sky130_fd_sc_hd__mux2_1
X_07497_ top.dut.bit_buf\[0\] net38 net714 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__mux2_1
X_06448_ top.hist_data_o\[14\] _03255_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09167_ _02969_ _02993_ top.cb_syn.curr_state\[2\] net464 vssd1 vssd1 vccd1 vccd1
+ _05167_ sky130_fd_sc_hd__and4b_1
X_06379_ _02594_ net444 top.histogram.state\[3\] vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__or3b_4
XANTENNA__06870__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08118_ net515 net523 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or2_2
X_09098_ net546 _02839_ _05118_ top.sram_interface.word_cnt\[14\] vssd1 vssd1 vccd1
+ vccd1 _05119_ sky130_fd_sc_hd__a22o_1
X_08049_ net523 _02969_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__and2_1
X_11060_ clknet_leaf_48_clk _01625_ _00450_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10011_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold826_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ net924 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
X_10913_ clknet_leaf_107_clk net955 _00303_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ clknet_leaf_108_clk _01438_ _00234_ vssd1 vssd1 vccd1 vccd1 top.path\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10775_ clknet_leaf_109_clk _01381_ _00165_ vssd1 vssd1 vccd1 vccd1 top.path\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__A1 top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11327_ clknet_leaf_88_clk _01892_ _00717_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11258_ clknet_leaf_79_clk _01823_ _00648_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_11189_ clknet_leaf_33_clk _01754_ _00579_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10209_ net824 net659 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__and2_1
XANTENNA__05719__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05750_ _02783_ _02793_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_19_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09330__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05681_ top.hTree.node_reg\[40\] net308 _02740_ net468 vssd1 vssd1 vccd1 vccd1 _02741_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07420_ _03412_ net149 _02523_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_46_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07351_ _03855_ _03858_ _03862_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nand3_1
X_06302_ top.hist_addr\[4\] _03098_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__xor2_1
X_07282_ _03880_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or2_1
X_06233_ _02585_ _03057_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__nor2_1
XANTENNA__06852__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09021_ top.WB.CPU_DAT_O\[29\] net1328 net314 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold201 top.cb_syn.char_path\[30\] vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09397__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06164_ net459 net361 _03038_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a21oi_1
Xhold212 top.cb_syn.char_path\[77\] vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 net64 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 top.path\[59\] vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
X_06095_ net550 _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__and2_1
Xhold245 net81 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 top.path\[14\] vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 top.path\[20\] vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 top.hTree.tree_reg\[3\] vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08357__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout703 net711 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_2
X_09923_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__and2_1
Xhold289 top.path\[1\] vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 net715 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
X_09854_ net867 net702 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__and2_1
X_11898__929 vssd1 vssd1 vccd1 vccd1 net929 _11898__929/LO sky130_fd_sc_hd__conb_1
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_2
Xfanout736 net796 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_0_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_2
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_2
X_08805_ top.path\[46\] top.path\[47\] net510 vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09785_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__and2_1
X_06997_ _02510_ net125 net123 _03683_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout564_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05591__B1 _02664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ top.path\[48\] net404 net324 top.path\[49\] net429 vssd1 vssd1 vccd1 vccd1
+ _04925_ sky130_fd_sc_hd__o221a_1
X_05948_ top.compVal\[13\] net161 net146 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 _02230_ sky130_fd_sc_hd__a22o_1
X_08667_ net1621 _04866_ _04877_ _04861_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a22o_1
XANTENNA__06135__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05879_ net1718 top.WB.CPU_DAT_O\[19\] net350 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
X_07618_ _04185_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ top.cb_syn.char_path_n\[123\] top.cb_syn.char_path_n\[124\] top.cb_syn.char_path_n\[127\]
+ top.cb_syn.curr_path\[127\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__mux4_1
XANTENNA__05894__A1 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _04147_ _04148_ net290 vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08293__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net862 net697 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__and2_1
XANTENNA__08832__A1 top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09719__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ top.header_synthesis.write_num_lefts _03375_ _05196_ vssd1 vssd1 vccd1 vccd1
+ top.header_synthesis.next_enable sky130_fd_sc_hd__a21bo_1
X_10491_ net779 net614 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__and2_1
XANTENNA__09388__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold776_A top.findLeastValue.sum\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05949__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold790 top.cb_syn.char_path_n\[76\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ clknet_leaf_50_clk _01677_ _00502_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_11043_ clknet_leaf_38_clk _01608_ _00433_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08899__A1 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06374__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05582__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11945_ net908 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__07323__A1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05885__A1 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05503__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ net879 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
X_10827_ clknet_leaf_113_clk _01421_ _00217_ vssd1 vssd1 vccd1 vccd1 top.path\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10758_ clknet_leaf_12_clk _00039_ _00148_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06834__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ clknet_leaf_107_clk _01320_ _00079_ vssd1 vssd1 vccd1 vccd1 top.path\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06920_ top.findLeastValue.val1\[37\] net137 net114 top.compVal\[37\] vssd1 vssd1
+ vccd1 vccd1 _01998_ sky130_fd_sc_hd__o22a_1
X_06851_ top.compVal\[28\] top.findLeastValue.val1\[28\] net151 vssd1 vssd1 vccd1
+ vccd1 _03631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ net788 net623 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__and2_1
XANTENNA__05573__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06782_ _03575_ _03576_ _03577_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__and3_1
X_05802_ top.sram_interface.write_counter_FLV\[2\] _02826_ vssd1 vssd1 vccd1 vccd1
+ _02827_ sky130_fd_sc_hd__xnor2_1
X_08521_ net1298 top.cb_syn.char_path_n\[38\] net239 vssd1 vssd1 vccd1 vccd1 _01521_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08737__S1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05733_ top.TRN_char_index\[5\] net43 net715 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
X_08452_ net1370 top.cb_syn.char_path_n\[107\] net244 vssd1 vssd1 vccd1 vccd1 _01590_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07314__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05876__A1 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05664_ top.histogram.sram_out\[11\] net357 net408 top.hTree.node_reg\[11\] _02726_
+ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a221o_1
X_07403_ _03662_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nor2_1
X_08383_ top.cb_syn.char_path_n\[13\] net383 net340 top.cb_syn.char_path_n\[11\] net187
+ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a221o_1
X_05595_ _02667_ _02668_ net467 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout145_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _03780_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07265_ _03724_ _03934_ _03722_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ top.WB.CPU_DAT_O\[16\] net1222 net365 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
X_06216_ net486 _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__or2_2
XFILLER_0_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ _03750_ _03762_ _03871_ _03760_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o211a_1
X_06147_ top.sram_interface.init_counter\[8\] top.sram_interface.init_counter\[7\]
+ _03023_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06078_ _02534_ top.cb_syn.i\[4\] vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__or2_1
X_09906_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__and2_1
Xfanout522 top.cb_syn.curr_state\[4\] vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_2
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_4
XANTENNA_fanout681_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout533 net535 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_4
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_1
Xfanout544 top.sram_interface.word_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_2
Xfanout555 net571 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_1
X_09837_ net849 net684 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__and2_1
Xfanout599 net601 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_2
Xfanout577 net584 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_2
Xfanout588 net631 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_2
X_09768_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__and2_1
XANTENNA__05564__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ net431 _04255_ net980 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__o21a_1
X_09699_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__and2_1
X_11730_ clknet_leaf_41_clk _02280_ _01120_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05867__A1 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11661_ clknet_leaf_115_clk _02211_ _01051_ vssd1 vssd1 vccd1 vccd1 top.path\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_10612_ net771 net606 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__and2_1
X_11592_ clknet_leaf_4_clk top.dut.out_valid_next _00982_ vssd1 vssd1 vccd1 vccd1
+ top.dut.out_valid sky130_fd_sc_hd__dfrtp_1
XANTENNA__06853__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ net730 net565 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__and2_1
XANTENNA__06816__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06292__A1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10474_ net855 net690 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11026_ clknet_leaf_60_clk _01591_ _00416_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09404__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ net891 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11859_ clknet_leaf_96_clk _02392_ _01231_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05380_ top.findLeastValue.val1\[8\] vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07050_ _02460_ _02486_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06001_ top.WB.CPU_DAT_O\[0\] net1343 net348 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_81_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XANTENNA__08980__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ net477 _04486_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__or2_1
X_07883_ net421 _04431_ _04432_ net263 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o211a_1
X_06903_ top.compVal\[2\] top.findLeastValue.val1\[2\] net153 vssd1 vssd1 vccd1 vccd1
+ _03657_ sky130_fd_sc_hd__mux2_1
X_09622_ net769 net604 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__and2_1
XANTENNA__09822__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05546__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06834_ top.findLeastValue.val2\[37\] net128 net118 _03622_ vssd1 vssd1 vccd1 vccd1
+ _02045_ sky130_fd_sc_hd__o22a_1
XANTENNA__08732__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09553_ net738 net573 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__and2_1
X_08504_ net1151 top.cb_syn.char_path_n\[55\] net232 vssd1 vssd1 vccd1 vccd1 _01538_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout262_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06765_ _02432_ top.findLeastValue.val2\[17\] _02471_ top.compVal\[16\] _03562_ vssd1
+ vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a221o_1
X_09484_ net765 net600 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__and2_1
X_05716_ _02768_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06239__A top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ _02409_ top.findLeastValue.val1\[38\] top.findLeastValue.val1\[33\] _02414_
+ _03492_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a221o_1
X_05647_ top.cb_syn.char_path\[13\] net547 net540 top.cb_syn.char_path\[77\] vssd1
+ vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a22o_1
X_08435_ net1303 top.cb_syn.char_path_n\[124\] net230 vssd1 vssd1 vccd1 vccd1 _01607_
+ sky130_fd_sc_hd__mux2_1
X_08366_ top.cb_syn.char_path_n\[21\] net194 _04745_ vssd1 vssd1 vccd1 vccd1 _01640_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05578_ top.histogram.sram_out\[25\] net359 net354 top.hTree.node_reg\[57\] vssd1
+ vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a22o_1
X_07317_ _03737_ _03955_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__nand2_1
X_08297_ top.cb_syn.char_path_n\[56\] net372 net329 top.cb_syn.char_path_n\[54\] net175
+ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a221o_1
XANTENNA__05797__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ _03915_ _03917_ net271 vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a21bo_1
X_07179_ _03848_ _03854_ _03853_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a21oi_4
X_10190_ net804 net639 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__and2_1
XANTENNA__08971__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__B2 top.findLeastValue.sum\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout341 _04637_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout374 _04612_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout363 _02571_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_2
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_4
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
XFILLER_0_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ clknet_leaf_69_clk _02263_ _01103_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11644_ clknet_leaf_109_clk _02194_ _01034_ vssd1 vssd1 vccd1 vccd1 top.path\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11575_ clknet_leaf_31_clk _02140_ _00965_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ net799 net634 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__and2_1
Xinput38 gpio_in[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
XANTENNA__09907__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ net803 net638 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07418__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05927__S _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ net769 net604 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__and2_1
XANTENNA__07765__A1 top.findLeastValue.sum\[44\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__A0 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05776__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__A1 top.cb_syn.char_path_n\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ clknet_leaf_35_clk net1440 _00399_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ net1105 _03329_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__xor2_1
X_05501_ net526 net527 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06481_ net297 _03246_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__nor2_1
X_08220_ net1794 net191 _04672_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05432_ net507 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08151_ top.cb_syn.char_path_n\[127\] net190 net326 vssd1 vssd1 vccd1 vccd1 _04638_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_99_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05363_ top.findLeastValue.val1\[44\] vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08082_ _04541_ _04548_ _04583_ _04584_ net1085 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__o32a_1
X_07102_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__inv_2
X_05294_ top.compVal\[36\] vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__inv_2
X_07033_ top.findLeastValue.val1\[46\] top.findLeastValue.val1\[45\] top.findLeastValue.val1\[44\]
+ top.findLeastValue.val1\[43\] vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07756__A1 top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ top.WB.CPU_DAT_O\[17\] top.cb_syn.h_element\[49\] net367 vssd1 vssd1 vccd1
+ vccd1 _01354_ sky130_fd_sc_hd__mux2_1
XANTENNA__05767__B1 _02806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ top.hTree.tree_reg\[10\] top.findLeastValue.sum\[10\] net283 vssd1 vssd1
+ vccd1 vccd1 _04474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout477_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ top.findLeastValue.sum\[24\] _04418_ net390 vssd1 vssd1 vccd1 vccd1 _04419_
+ sky130_fd_sc_hd__mux2_1
X_09605_ net725 net560 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07797_ net476 _04362_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__or2_1
X_06817_ top.compVal\[45\] top.findLeastValue.val1\[45\] net152 vssd1 vssd1 vccd1
+ vccd1 _03614_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09536_ net744 net579 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__and2_1
X_06748_ _03542_ _03543_ _03545_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21oi_1
X_09467_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__and2_1
X_08418_ top.cb_syn.char_index\[6\] _04774_ _04772_ vssd1 vssd1 vccd1 vccd1 _01617_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06679_ top.compVal\[41\] _02482_ _02483_ top.compVal\[40\] vssd1 vssd1 vccd1 vccd1
+ _03477_ sky130_fd_sc_hd__a22o_1
X_09398_ net400 _04272_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__nand2_1
X_08349_ top.cb_syn.char_path_n\[30\] net373 net327 top.cb_syn.char_path_n\[28\] net172
+ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11360_ clknet_leaf_94_clk _01925_ _00750_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[38\]
+ sky130_fd_sc_hd__dfrtp_2
X_10311_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08619__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ clknet_leaf_22_clk _01856_ _00681_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08944__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ net818 net653 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__and2_1
X_10173_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__and2_1
XANTENNA_input38_A gpio_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 net185 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout171 _02621_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
Xfanout193 net195 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XFILLER_0_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05930__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09121__B1 _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11627_ clknet_leaf_23_clk _02177_ _01017_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11558_ clknet_leaf_21_clk _02123_ _00948_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06238__A1 top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10509_ net754 net589 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold619 top.hTree.tree_reg\[18\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ clknet_leaf_94_clk _02054_ _00879_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[46\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05997__A0 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05461__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05749__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07720_ net387 _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__nand2_1
XANTENNA__06961__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05981_ top.WB.CPU_DAT_O\[20\] net1219 net345 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XANTENNA__09360__B1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ top.cb_syn.h_element\[55\] net525 _04180_ top.cb_syn.max_index\[1\] _04244_
+ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a221o_1
X_07582_ net517 top.cb_syn.h_element\[52\] net525 top.cb_syn.h_element\[61\] _04180_
+ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a221o_1
XANTENNA__07910__A1 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ _03396_ _03397_ _03398_ _03399_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09321_ net1035 net224 net216 _04491_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__a22o_1
X_06533_ _03335_ _03352_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__inv_2
X_06464_ net1278 _03306_ net300 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05415_ top.cb_syn.zeroes\[1\] vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__inv_2
XANTENNA__08218__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05421__A top.cb_syn.char_path_n\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08203_ top.cb_syn.char_path_n\[103\] net380 net337 top.cb_syn.char_path_n\[101\]
+ net183 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a221o_1
X_06395_ top.hist_data_o\[23\] _03259_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__and2_1
X_09183_ net248 _05058_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08134_ _04618_ _04620_ net172 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07426__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05346_ top.findLeastValue.val2\[34\] vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__inv_2
XANTENNA__07521__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08065_ _04566_ _04179_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__and2b_2
XANTENNA__05988__A0 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ top.findLeastValue.val2\[26\] top.findLeastValue.val2\[25\] top.findLeastValue.val2\[24\]
+ top.findLeastValue.val2\[23\] vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout594_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06952__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ top.WB.CPU_DAT_O\[1\] net1377 net320 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__mux2_1
X_07918_ net420 _04459_ _04460_ net262 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o211a_1
X_08898_ net1148 top.WB.CPU_DAT_O\[4\] net306 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__mux2_1
X_07849_ net434 net1495 net248 net1801 _04405_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a221o_1
XANTENNA__09351__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ clknet_leaf_28_clk top.header_synthesis.next_zero_count\[1\] _00250_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[1\] sky130_fd_sc_hd__dfrtp_1
X_09519_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__and2_1
X_10791_ clknet_leaf_114_clk _01397_ _00181_ vssd1 vssd1 vccd1 vccd1 top.path\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05691__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ clknet_leaf_101_clk _01977_ _00802_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[16\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06861__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ clknet_leaf_77_clk _01908_ _00733_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05979__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ clknet_leaf_44_clk _01839_ _00664_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08393__A1 top.cb_syn.char_path_n\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__and2_1
XANTENNA__06943__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__A1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 top.sram_interface.CB_read_counter vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__and2_1
XANTENNA__09342__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ clknet_leaf_65_clk net1348 _00379_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05682__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06180_ top.TRN_char_index\[3\] net445 _03053_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__and3_1
Xhold416 top.cb_syn.char_path\[75\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08620__A2 top.cb_syn.char_path_n\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 top.WB.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 top.hTree.tree_reg\[32\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 top.path\[88\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 top.path\[61\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_09870_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__and2_1
X_08821_ top.path\[100\] net405 net325 top.path\[101\] net505 vssd1 vssd1 vccd1 vccd1
+ _05010_ sky130_fd_sc_hd__o221a_1
XANTENNA__06934__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05964_ top.CB_read_complete _02911_ _02902_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__o21ba_1
X_08752_ top.path\[30\] top.path\[31\] net511 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__mux2_1
X_08683_ top.cb_syn.i\[2\] top.cb_syn.i\[1\] top.cb_syn.i\[0\] top.cb_syn.i\[3\] vssd1
+ vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a31o_1
X_07703_ net473 _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XANTENNA__09333__B1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ net1500 _04230_ _04212_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05895_ net1577 top.WB.CPU_DAT_O\[3\] net349 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ _04161_ _04164_ _04110_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06516_ net1505 _03341_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__xor2_1
X_09304_ _05247_ _05238_ top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 _05248_
+ sky130_fd_sc_hd__mux2_1
X_07496_ net1620 top.dut.out_valid_next _04061_ _04078_ _04097_ vssd1 vssd1 vccd1
+ vccd1 _01862_ sky130_fd_sc_hd__o221a_1
X_09235_ top.header_synthesis.header\[6\] top.cb_syn.char_index\[6\] net490 vssd1
+ vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__mux2_1
X_06447_ net1125 _03295_ net300 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XANTENNA__05673__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ top.cb_syn.char_path_n\[1\] net515 net464 _04201_ vssd1 vssd1 vccd1 vccd1
+ _05166_ sky130_fd_sc_hd__and4b_1
X_06378_ net439 top.histogram.state\[3\] net360 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__and3_4
X_08117_ net515 top.cb_syn.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09097_ net443 net462 net451 _05107_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a211o_1
X_05329_ top.compVal\[0\] vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08048_ _04558_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__inv_2
X_10010_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__and2_1
X_09999_ net855 net690 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__and2_1
XANTENNA__06925__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06138__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ clknet_leaf_106_clk net953 _00302_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06153__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net923 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_80_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10843_ clknet_leaf_108_clk _01437_ _00233_ vssd1 vssd1 vccd1 vccd1 top.path\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10774_ clknet_leaf_113_clk _01380_ _00164_ vssd1 vssd1 vccd1 vccd1 top.path\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05664__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11326_ clknet_leaf_88_clk _01891_ _00716_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11257_ clknet_leaf_80_clk net1586 _00647_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_11188_ clknet_leaf_33_clk _01753_ _00578_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09407__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ net824 net659 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__and2_1
X_10139_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__and2_1
XANTENNA__10142__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05680_ _02738_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ net269 _03996_ _03997_ net275 net1709 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a32o_1
XANTENNA__08826__C1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06301_ top.sram_interface.init_counter\[4\] _03020_ vssd1 vssd1 vccd1 vccd1 _03171_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09094__A2 top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07281_ _03875_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__nand2_1
X_09020_ top.WB.CPU_DAT_O\[30\] net1135 net314 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
XANTENNA__05655__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06232_ top.cb_syn.max_index\[7\] _03102_ _03104_ top.hTree.nullSumIndex\[6\] vssd1
+ vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold202 top.cb_syn.char_path\[0\] vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
X_06163_ net459 net534 _02787_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__and3_1
Xhold235 top.cb_syn.char_path\[88\] vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 top.hTree.tree_reg\[55\] vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 top.hTree.nulls\[59\] vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 top.cb_syn.char_path\[79\] vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
X_06094_ _02969_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__nor2_1
Xhold268 top.path\[52\] vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 top.path\[44\] vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 top.cb_syn.char_path\[24\] vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout704 net711 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_2
X_09922_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__and2_1
Xfanout715 net37 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_2
X_09853_ net867 net702 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__and2_1
Xfanout726 net736 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_2
Xfanout737 net740 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_2
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_2
X_09784_ net871 net706 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout292_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net777 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_1
X_08804_ _04990_ _04991_ _04992_ net503 top.translation.index\[2\] vssd1 vssd1 vccd1
+ vccd1 _04993_ sky130_fd_sc_hd__a221o_1
X_06996_ top.cw1\[2\] net148 _03662_ top.findLeastValue.histo_index\[2\] vssd1 vssd1
+ vccd1 vccd1 _03683_ sky130_fd_sc_hd__a22o_1
X_08735_ net426 _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__or2_1
XANTENNA__09306__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05947_ top.compVal\[14\] net161 net146 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 _02231_ sky130_fd_sc_hd__a22o_1
X_08666_ top.cb_syn.cb_enable _04792_ _04868_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05878_ net1760 top.WB.CPU_DAT_O\[20\] net350 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
X_08597_ _04811_ _04813_ _04816_ top.cb_syn.end_cnt\[3\] _02540_ vssd1 vssd1 vccd1
+ vccd1 _04817_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07617_ top.cb_syn.max_index\[5\] _04184_ top.cb_syn.max_index\[6\] vssd1 vssd1 vccd1
+ vccd1 _04216_ sky130_fd_sc_hd__o21ai_1
X_07548_ top.cb_syn.char_path_n\[2\] top.cb_syn.char_path_n\[1\] top.cb_syn.char_path_n\[4\]
+ top.cb_syn.char_path_n\[3\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08817__C1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08904__B net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ _04048_ _04069_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__or2_1
XANTENNA__05646__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11946__909 vssd1 vssd1 vccd1 vccd1 _11946__909/HI net909 sky130_fd_sc_hd__conb_1
X_09218_ _03371_ _03388_ _05195_ net291 top.header_synthesis.write_num_lefts vssd1
+ vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a311o_1
X_10490_ net779 net614 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09149_ net537 _05108_ _05154_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07399__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ clknet_leaf_50_clk _01676_ _00501_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[57\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold791 top.cw1\[7\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold780 top.compVal\[11\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
X_11042_ clknet_leaf_38_clk _01607_ _00432_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_110_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09751__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ net907 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA__07859__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ clknet_leaf_120_clk net878 _01247_ vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07323__A2 _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05503__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ clknet_leaf_112_clk _01420_ _00216_ vssd1 vssd1 vccd1 vccd1 top.path\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10757_ clknet_leaf_13_clk _00052_ _00147_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ clknet_leaf_11_clk _01319_ _00078_ vssd1 vssd1 vccd1 vccd1 top.path\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ clknet_leaf_14_clk _01874_ _00699_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08339__B2 top.cb_syn.char_path_n\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ top.findLeastValue.val2\[29\] net127 net118 _03630_ vssd1 vssd1 vccd1 vccd1
+ _02037_ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07880__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05801_ top.sram_interface.write_counter_FLV\[1\] top.sram_interface.write_counter_FLV\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06781_ top.compVal\[24\] _02468_ _03567_ _03570_ _03571_ vssd1 vssd1 vccd1 vccd1
+ _03579_ sky130_fd_sc_hd__o2111a_1
X_08520_ net1349 top.cb_syn.char_path_n\[39\] net239 vssd1 vssd1 vccd1 vccd1 _01522_
+ sky130_fd_sc_hd__mux2_1
X_05732_ top.TRN_char_index\[6\] net35 net714 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
X_08451_ net1210 top.cb_syn.char_path_n\[108\] net244 vssd1 vssd1 vccd1 vccd1 _01591_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05663_ top.hTree.node_reg\[43\] net308 _02725_ net469 vssd1 vssd1 vccd1 vccd1 _02726_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ top.findLeastValue.histo_index\[7\] _02523_ net148 vssd1 vssd1 vccd1 vccd1
+ _04031_ sky130_fd_sc_hd__mux2_1
X_08382_ top.cb_syn.char_path_n\[13\] net204 _04753_ vssd1 vssd1 vccd1 vccd1 _01632_
+ sky130_fd_sc_hd__o21a_1
X_05594_ top.cb_syn.char_path\[54\] net530 net311 top.cb_syn.char_path\[118\] vssd1
+ vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ _03781_ _03979_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08814__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ _03727_ _03730_ _03933_ _03728_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06215_ top.findLeastValue.histo_index\[2\] net487 top.findLeastValue.histo_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__and3_1
X_09003_ top.WB.CPU_DAT_O\[17\] net1260 net365 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
X_07195_ _03750_ _03870_ _03789_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__or3b_1
X_06146_ top.sram_interface.init_counter\[6\] top.sram_interface.init_counter\[5\]
+ _03021_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__and3_1
X_06077_ _02534_ top.cb_syn.i\[4\] vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__nand2_1
X_11906__937 vssd1 vssd1 vccd1 vccd1 net937 _11906__937/LO sky130_fd_sc_hd__conb_1
X_09905_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__and2_1
Xfanout501 top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_4
Xfanout523 top.cb_syn.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
XANTENNA__05800__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout512 top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout674_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_2
Xfanout556 net558 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_2
X_09836_ net849 net684 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__and2_1
XANTENNA__07790__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout567 net571 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_2
Xfanout578 net583 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_2
X_09767_ net792 net627 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout841_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ top.findLeastValue.histo_index\[5\] _03670_ _03668_ vssd1 vssd1 vccd1 vccd1
+ _03677_ sky130_fd_sc_hd__a21bo_1
X_09698_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__and2_1
X_08718_ _04896_ _04907_ _04911_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_29_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _02538_ _04791_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ clknet_leaf_114_clk _02210_ _01050_ vssd1 vssd1 vccd1 vccd1 top.path\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_11591_ clknet_leaf_31_clk _02156_ _00981_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10611_ net743 net578 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_115_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ net731 net566 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__and2_1
XANTENNA__06816__B2 top.findLeastValue.val1\[46\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ net855 net690 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11025_ clknet_leaf_61_clk _01590_ _00415_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_11927_ net890 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_86_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ clknet_leaf_113_clk _02391_ _01230_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_10809_ clknet_leaf_32_clk _00007_ _00199_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11789_ clknet_leaf_95_clk _02323_ _01161_ vssd1 vssd1 vccd1 vccd1 top.compVal\[38\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_19 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_106_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06000_ top.WB.CPU_DAT_O\[1\] net1339 net347 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
X_07951_ top.hTree.tree_reg\[7\] top.findLeastValue.sum\[7\] net266 vssd1 vssd1 vccd1
+ vccd1 _04487_ sky130_fd_sc_hd__mux2_1
XANTENNA__06991__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06902_ top.findLeastValue.val2\[3\] net130 net120 _03656_ vssd1 vssd1 vccd1 vccd1
+ _02011_ sky130_fd_sc_hd__o22a_1
X_07882_ net478 _04430_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ net770 net605 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__and2_1
XANTENNA__07535__A2 top.cb_syn.char_path_n\[96\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ top.compVal\[37\] top.findLeastValue.val1\[37\] net152 vssd1 vssd1 vccd1
+ vccd1 _03622_ sky130_fd_sc_hd__mux2_1
X_09552_ net738 net573 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__and2_1
X_06764_ top.findLeastValue.val2\[17\] _02432_ top.compVal\[18\] _02470_ vssd1 vssd1
+ vccd1 vccd1 _03562_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__05424__A top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ net1087 top.cb_syn.char_path_n\[56\] net233 vssd1 vssd1 vccd1 vccd1 _01539_
+ sky130_fd_sc_hd__mux2_1
X_05715_ top.cb_syn.char_path\[34\] net530 net311 top.cb_syn.char_path\[98\] vssd1
+ vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09483_ net765 net600 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__and2_1
X_06695_ _03479_ _03491_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__nand2b_1
X_08434_ net1413 top.cb_syn.char_path_n\[125\] net230 vssd1 vssd1 vccd1 vccd1 _01608_
+ sky130_fd_sc_hd__mux2_1
X_05646_ net1316 net171 _02711_ net211 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a22o_1
XANTENNA__08735__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ top.cb_syn.char_path_n\[22\] net377 net330 top.cb_syn.char_path_n\[20\] net177
+ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a221o_1
X_05577_ _02652_ _02653_ net466 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ net1648 net274 net268 _03972_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08296_ top.cb_syn.char_path_n\[56\] net195 _04710_ vssd1 vssd1 vccd1 vccd1 _01675_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07247_ _03920_ _03921_ net271 net277 net1732 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a32o_1
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ _03803_ _03811_ _03849_ _03851_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__and4b_1
XANTENNA__08420__A0 top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06129_ net1226 net164 _03016_ net207 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a22o_1
Xfanout331 net341 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout320 net322 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout353 _02881_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_4
Xfanout364 _02570_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_2
Xfanout342 _04048_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout397 _02981_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_4
Xfanout386 _04612_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_2
X_09819_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_70_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ clknet_leaf_81_clk _02262_ _01102_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11643_ clknet_leaf_109_clk _02193_ _01033_ vssd1 vssd1 vccd1 vccd1 top.path\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ clknet_leaf_27_clk _02139_ _00964_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
X_10525_ net799 net634 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__and2_1
X_10456_ net802 net637 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__and2_1
X_10387_ net769 net604 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__and2_1
XANTENNA__05776__B2 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ clknet_leaf_36_clk _01573_ _00398_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08573__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05500_ net451 net545 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__nand2_2
XFILLER_0_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06480_ top.hist_data_o\[2\] top.hist_data_o\[1\] top.hist_data_o\[0\] top.hist_data_o\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a31o_1
X_05431_ net504 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__inv_2
X_08150_ _02538_ net371 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07101_ top.findLeastValue.val2\[21\] top.findLeastValue.val1\[21\] vssd1 vssd1 vccd1
+ vccd1 _03777_ sky130_fd_sc_hd__nand2_1
X_05362_ top.findLeastValue.val2\[0\] vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08081_ _04549_ _04552_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__nor2_1
X_05293_ top.compVal\[37\] vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__inv_2
X_07032_ top.findLeastValue.val1\[42\] top.findLeastValue.val1\[41\] top.findLeastValue.val1\[40\]
+ top.findLeastValue.val1\[39\] vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ top.WB.CPU_DAT_O\[18\] top.cb_syn.h_element\[50\] net367 vssd1 vssd1 vccd1
+ vccd1 _01355_ sky130_fd_sc_hd__mux2_1
XANTENNA__05767__B2 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ net437 net1600 net251 top.findLeastValue.sum\[11\] _04473_ vssd1 vssd1 vccd1
+ vccd1 _01800_ sky130_fd_sc_hd__a221o_1
X_07865_ top.hTree.tree_reg\[24\] top.findLeastValue.sum\[24\] net282 vssd1 vssd1
+ vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout372_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ net749 net584 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__and2_1
X_07796_ top.hTree.tree_reg\[38\] top.findLeastValue.sum\[38\] net266 vssd1 vssd1
+ vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
X_06816_ top.findLeastValue.val2\[46\] net128 net119 top.findLeastValue.val1\[46\]
+ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__and2_1
X_06747_ _02438_ top.findLeastValue.val2\[8\] top.findLeastValue.val2\[7\] _02439_
+ _03532_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a221o_1
X_09466_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__and2_1
X_06678_ _03458_ _03463_ _03470_ _03475_ _03465_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05629_ top.cb_syn.char_path\[16\] net547 net540 top.cb_syn.char_path\[80\] vssd1
+ vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a22o_1
X_08417_ top.cb_syn.h_element\[61\] top.cb_syn.h_element\[52\] net517 vssd1 vssd1
+ vccd1 vccd1 _04774_ sky130_fd_sc_hd__mux2_1
X_09397_ net990 net221 _05277_ _05278_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout804_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ top.cb_syn.char_path_n\[30\] net191 _04736_ vssd1 vssd1 vccd1 vccd1 _01649_
+ sky130_fd_sc_hd__o21a_1
X_08279_ top.cb_syn.char_path_n\[65\] net372 net329 top.cb_syn.char_path_n\[63\] net175
+ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__a221o_1
X_10310_ net839 net674 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__and2_1
X_11290_ clknet_leaf_20_clk _01855_ _00680_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09296__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ net805 net640 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__and2_1
X_10172_ net807 net642 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__and2_1
XANTENNA__06859__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout172 net174 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net185 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
XANTENNA__08157__C1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout161 _02908_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_4
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05930__B2 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11930__893 vssd1 vssd1 vccd1 vccd1 _11930__893/HI net893 sky130_fd_sc_hd__conb_1
X_11626_ clknet_leaf_23_clk _02176_ _01016_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05694__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ clknet_leaf_7_clk _02122_ _00947_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
Xhold609 _01802_ vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10508_ net754 net589 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__and2_1
X_11488_ clknet_leaf_94_clk _02053_ _00878_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[45\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10439_ net819 net654 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__and2_1
XANTENNA__06946__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05980_ top.WB.CPU_DAT_O\[21\] net1051 net345 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XANTENNA__06961__A3 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ _02543_ top.cb_syn.max_index\[1\] top.cb_syn.h_element\[46\] net517 vssd1
+ vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__a2bb2o_1
X_07581_ _04178_ _04179_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__or2_2
X_06601_ top.compVal\[3\] top.compVal\[2\] top.compVal\[1\] top.compVal\[0\] vssd1
+ vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09320_ net1049 net224 net216 _04495_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a22o_1
X_06532_ net1798 _03334_ net1502 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__a21oi_1
X_09251_ _02557_ _05212_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__nor2_1
X_08202_ top.cb_syn.char_path_n\[103\] net201 _04663_ vssd1 vssd1 vccd1 vccd1 _01722_
+ sky130_fd_sc_hd__o21a_1
X_06463_ top.hist_data_o\[9\] _03250_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_16_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05414_ top.cb_syn.zeroes\[2\] vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__inv_2
XANTENNA__05685__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06394_ top.hist_data_o\[22\] top.hist_data_o\[21\] _03258_ vssd1 vssd1 vccd1 vccd1
+ _03259_ sky130_fd_sc_hd__and3_1
X_09182_ net287 _05050_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__and3_1
X_08133_ net1723 _04622_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07426__B2 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05345_ top.findLeastValue.val2\[35\] vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout120_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07521__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _04179_ _04574_ _04566_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout218_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _03687_ _03688_ _03689_ _03690_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout587_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06937__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ top.WB.CPU_DAT_O\[2\] net1258 net320 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__mux2_1
XANTENNA__08154__A2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ net479 _04458_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_95_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
X_08897_ net1110 top.WB.CPU_DAT_O\[5\] net305 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__mux2_1
X_07848_ net417 _04403_ _04404_ net256 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__o211a_1
X_07779_ net437 net1569 net251 top.findLeastValue.sum\[42\] _04349_ vssd1 vssd1 vccd1
+ vccd1 _01831_ sky130_fd_sc_hd__a221o_1
XANTENNA__08907__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ net734 net569 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__and2_1
X_10790_ clknet_leaf_117_clk _01396_ _00180_ vssd1 vssd1 vccd1 vccd1 top.path\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ net750 net585 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__and2_1
XANTENNA__05676__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07417__A1 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ clknet_leaf_86_clk _01976_ _00801_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[15\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__08642__B _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11342_ clknet_leaf_77_clk _01907_ _00732_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11273_ clknet_leaf_44_clk _01838_ _00663_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06162__B top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__and2_1
X_10155_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__and2_1
XANTENNA__06928__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05600__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 _02251_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ net823 net658 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_86_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10988_ clknet_leaf_70_clk net1178 _00378_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05667__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11609_ clknet_leaf_21_clk _02159_ _00999_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08620__A3 top.cb_syn.char_path_n\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 top.cb_syn.char_path\[41\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 top.cb_syn.char_path\[9\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 net71 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 top.sram_interface.zero_cnt\[2\] vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09030__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06919__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ top.path\[102\] top.path\[103\] net512 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__mux2_1
X_05963_ _02910_ _02899_ _02898_ top.sram_interface.CB_read_counter vssd1 vssd1 vccd1
+ vccd1 _02911_ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_77_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
X_08751_ net425 _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__or2_1
X_08682_ _04883_ _04886_ _04889_ _04879_ net1783 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a32o_1
X_07702_ top.findLeastValue.least1\[1\] net264 _04285_ vssd1 vssd1 vccd1 vccd1 _04287_
+ sky130_fd_sc_hd__a21oi_1
X_05894_ top.hist_data_o\[4\] top.WB.CPU_DAT_O\[4\] net349 vssd1 vssd1 vccd1 vccd1
+ _02256_ sky130_fd_sc_hd__mux2_1
X_07633_ top.cb_syn.max_index\[4\] _04181_ _04226_ _04229_ vssd1 vssd1 vccd1 vccd1
+ _04230_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout168_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ _04162_ _04163_ net290 vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09303_ _05243_ _05246_ net502 vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__mux2_1
X_06515_ _03342_ net1449 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__nor2_1
XANTENNA__05432__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ top.dut.bits_in_buf_next\[1\] _04087_ _04096_ _04046_ vssd1 vssd1 vccd1 vccd1
+ _04097_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout335_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05658__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09234_ net1083 _05203_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[5\]
+ sky130_fd_sc_hd__mux2_1
X_06446_ top.hist_data_o\[15\] _03256_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09165_ net424 _02890_ _05084_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__or3b_1
X_08116_ _02539_ _02886_ _04606_ _04608_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a311o_1
X_06377_ net1174 net164 _03242_ net208 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a22o_1
XANTENNA__06870__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09096_ net447 net1581 net527 _02795_ _05117_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__a221o_1
X_05328_ top.compVal\[1\] vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__inv_2
X_08047_ net523 _02995_ _04204_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_116_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09574__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09021__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net861 net696 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__and2_1
X_08949_ top.WB.CPU_DAT_O\[19\] net1124 net318 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__mux2_1
XANTENNA__08780__C1 top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07822__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ clknet_leaf_11_clk net977 _00301_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ net922 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XANTENNA_hold714_A top.hTree.node_reg\[47\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ clknet_leaf_108_clk _01436_ _00232_ vssd1 vssd1 vccd1 vccd1 top.path\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10773_ clknet_leaf_113_clk _01379_ _00163_ vssd1 vssd1 vccd1 vccd1 top.path\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11325_ clknet_leaf_89_clk _01890_ _00715_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07810__A1 top.findLeastValue.sum\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ clknet_leaf_79_clk _01821_ _00646_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08366__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11187_ clknet_leaf_33_clk _01752_ _00577_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06377__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ net825 net660 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__and2_1
X_10138_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__and2_1
XANTENNA__10142__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__C1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
X_10069_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06129__B2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06300_ _03167_ _03169_ net459 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__o21a_1
X_07280_ _03877_ _03884_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_100_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06231_ net526 top.sram_interface.word_cnt\[13\] _03103_ vssd1 vssd1 vccd1 vccd1
+ _03104_ sky130_fd_sc_hd__or3_4
XANTENNA__06852__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06162_ top.findLeastValue.histo_index\[8\] top.findLeastValue.histo_index\[7\] vssd1
+ vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06093_ _02979_ net394 _02984_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__and4b_1
Xhold225 top.cb_syn.char_path\[73\] vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A1 top.findLeastValue.sum\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 top.path\[56\] vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 top.path\[82\] vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 top.cb_syn.char_path\[17\] vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__and2_1
Xhold269 top.cb_syn.char_path\[20\] vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 top.cb_syn.char_path\[60\] vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09003__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07907__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 top.path\[2\] vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08357__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 net710 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_2
X_09852_ net863 net698 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__and2_1
Xfanout716 net718 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_2
Xfanout738 net740 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_2
Xfanout749 net796 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_2
Xfanout727 net729 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_2
X_09783_ net870 net705 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__and2_1
X_08803_ top.path\[72\] top.path\[73\] top.path\[74\] top.path\[75\] net511 net507
+ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__mux4_1
X_06995_ _02509_ net125 net123 _03682_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a2bb2o_1
X_08734_ top.path\[50\] top.path\[51\] net511 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__mux2_1
XANTENNA__05591__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05946_ top.compVal\[15\] net161 net146 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 _02232_ sky130_fd_sc_hd__a22o_1
X_08665_ net499 _04868_ _04876_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a21bo_1
X_05877_ net1625 top.WB.CPU_DAT_O\[21\] net350 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XANTENNA__07868__A1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_A top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ _04814_ _04815_ net497 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__mux2_1
X_07616_ net518 top.cb_syn.h_element\[51\] net525 top.cb_syn.h_element\[60\] _04180_
+ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ top.cb_syn.char_path_n\[6\] top.cb_syn.char_path_n\[5\] top.cb_syn.char_path_n\[8\]
+ top.cb_syn.char_path_n\[7\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ _04073_ _04082_ net342 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ top.header_synthesis.write_zeroes _05193_ net491 _02565_ vssd1 vssd1 vccd1
+ vccd1 _05195_ sky130_fd_sc_hd__a211o_1
X_06429_ _03260_ _03285_ net301 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__and3b_1
XANTENNA__09242__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ top.sram_interface.CB_write_counter\[1\] top.sram_interface.CB_write_counter\[0\]
+ _05098_ _05153_ net317 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ net442 net451 _05096_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ clknet_leaf_49_clk _01675_ _00500_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold770 top.cb_syn.char_path_n\[91\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 top.findLeastValue.sum\[45\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07817__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ clknet_leaf_37_clk _01606_ _00431_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[123\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold792 top.findLeastValue.sum\[8\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08753__C1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05582__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06867__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ net906 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11874_ clknet_leaf_1_clk top.dut.bits_in_buf_next\[2\] _01246_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bits_in_buf\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_43_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ clknet_leaf_97_clk _01419_ _00215_ vssd1 vssd1 vccd1 vccd1 top.path\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10756_ clknet_leaf_10_clk _00051_ _00146_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06834__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687_ clknet_leaf_11_clk _01318_ _00077_ vssd1 vssd1 vccd1 vccd1 top.path\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ clknet_leaf_14_clk _01873_ _00698_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11239_ clknet_leaf_67_clk net1437 _00629_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10153__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05800_ net533 net527 _02823_ net455 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__o211a_1
XANTENNA__05573__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06780_ top.compVal\[21\] top.findLeastValue.val2\[21\] vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__nand2b_1
X_05731_ net1473 net170 _02782_ net209 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__a22o_1
X_05662_ _02723_ _02724_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__or2_1
X_08450_ net1266 top.cb_syn.char_path_n\[109\] net244 vssd1 vssd1 vccd1 vccd1 _01592_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08381_ top.cb_syn.char_path_n\[14\] net384 net340 top.cb_syn.char_path_n\[12\] net187
+ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a221o_1
X_07401_ top.findLeastValue.least2\[8\] _03611_ net117 _04030_ vssd1 vssd1 vccd1 vccd1
+ _01886_ sky130_fd_sc_hd__o22a_1
X_05593_ top.cb_syn.char_path\[22\] net548 net539 top.cb_syn.char_path\[86\] vssd1
+ vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
X_07332_ net1733 net275 net269 _03984_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08275__B2 top.cb_syn.char_path_n\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07263_ _03890_ _03893_ _03732_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__a21o_1
X_09002_ top.WB.CPU_DAT_O\[18\] net1445 net365 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
X_06214_ net487 top.findLeastValue.histo_index\[0\] vssd1 vssd1 vccd1 vccd1 _03087_
+ sky130_fd_sc_hd__nand2_1
X_07194_ _03757_ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06145_ top.sram_interface.init_counter\[5\] _03021_ vssd1 vssd1 vccd1 vccd1 _03022_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06076_ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__and2_1
Xfanout524 net525 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_2
Xfanout502 top.translation.index\[3\] vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
Xfanout513 top.translation.resEn vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_2
X_09835_ net849 net684 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__and2_1
Xfanout546 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_4
Xfanout535 top.sram_interface.word_cnt\[8\] vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_2
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 net583 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_1
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_2
X_09766_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__and2_1
XANTENNA__05564__A2 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06978_ net1617 _03671_ _03676_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__o21ba_1
X_09697_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__and2_1
X_08717_ _02544_ _03389_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__nand2_1
X_05929_ _02906_ net158 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _02888_ _04863_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_1_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ net496 _04798_ _02541_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__a21o_1
X_11590_ clknet_leaf_32_clk _02155_ _00980_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10610_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net730 net565 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__and2_1
XANTENNA__06816__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ net830 net665 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__and2_1
XANTENNA__08650__B _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold781_A top.findLeastValue.sum\[45\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11024_ clknet_leaf_61_clk _01589_ _00414_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07981__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05555__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11926_ net889 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_86_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ clknet_leaf_112_clk _02390_ _01229_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_10808_ clknet_leaf_26_clk _00006_ _00198_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.finished
+ sky130_fd_sc_hd__dfrtp_1
X_11788_ clknet_leaf_95_clk _02322_ _01160_ vssd1 vssd1 vccd1 vccd1 top.compVal\[37\]
+ sky130_fd_sc_hd__dfrtp_4
X_10739_ clknet_leaf_4_clk _00029_ _00129_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__09301__S0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ top.hTree.tree_reg\[7\] top.findLeastValue.sum\[7\] net284 vssd1 vssd1 vccd1
+ vccd1 _04486_ sky130_fd_sc_hd__mux2_1
XANTENNA__07891__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ top.compVal\[3\] top.findLeastValue.val1\[3\] net153 vssd1 vssd1 vccd1 vccd1
+ _03656_ sky130_fd_sc_hd__mux2_1
X_07881_ top.hTree.tree_reg\[21\] top.findLeastValue.sum\[21\] net264 vssd1 vssd1
+ vccd1 vccd1 _04431_ sky130_fd_sc_hd__mux2_1
X_09620_ net770 net605 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__and2_1
XANTENNA__05546__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ top.findLeastValue.val2\[38\] net128 net119 _03621_ vssd1 vssd1 vccd1 vccd1
+ _02046_ sky130_fd_sc_hd__o22a_1
X_09551_ net737 net572 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__and2_1
X_06763_ _02432_ top.findLeastValue.val2\[17\] vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nand2_1
X_08502_ net1336 top.cb_syn.char_path_n\[57\] net231 vssd1 vssd1 vccd1 vccd1 _01540_
+ sky130_fd_sc_hd__mux2_1
X_05714_ top.cb_syn.char_path\[2\] net548 net539 top.cb_syn.char_path\[66\] vssd1
+ vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a22o_1
X_09482_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__and2_1
X_06694_ _02412_ top.findLeastValue.val1\[35\] top.findLeastValue.val1\[34\] _02413_
+ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__a22o_1
X_08433_ net1139 top.cb_syn.char_path_n\[126\] net230 vssd1 vssd1 vccd1 vccd1 _01609_
+ sky130_fd_sc_hd__mux2_1
X_05645_ top.hTree.node_reg\[46\] net355 _02709_ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout150_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ net1766 net195 _04744_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__o21a_1
X_05576_ top.cb_syn.char_path\[25\] net546 net312 top.cb_syn.char_path\[121\] vssd1
+ vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _03753_ _03956_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08799__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08295_ top.cb_syn.char_path_n\[57\] net371 net329 top.cb_syn.char_path_n\[55\] net175
+ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08751__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ _03393_ _03718_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_1
XANTENNA__05482__B2 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07177_ _03803_ _03816_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__and2b_1
X_06128_ net533 net527 _03013_ _03015_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06059_ top.cb_syn.zeroes\[3\] _02557_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__nor2_1
Xfanout332 net335 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
Xfanout310 net311 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09582__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout354 net356 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
Xfanout343 _04042_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_2
Xfanout376 net386 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
X_09818_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__and2_1
Xfanout387 net389 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_2
Xfanout398 net399 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_2
X_09749_ net863 net698 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__and2_1
XANTENNA__08926__A _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11711_ clknet_leaf_81_clk _02261_ _01101_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11642_ clknet_leaf_110_clk _02192_ _01032_ vssd1 vssd1 vccd1 vccd1 top.path\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11573_ clknet_leaf_31_clk _02138_ _00963_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07976__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ net800 net635 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__and2_1
XANTENNA__05473__B2 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ net802 net637 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__and2_1
X_10386_ net762 net597 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__and2_1
XANTENNA__06973__A1 top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05776__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__S _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ clknet_leaf_36_clk _01572_ _00397_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08573__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ net940 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05430_ net503 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__inv_2
X_05361_ top.findLeastValue.val2\[3\] vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__inv_2
XANTENNA__05700__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07886__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07100_ top.findLeastValue.val2\[19\] top.findLeastValue.val1\[19\] _03774_ _03775_
+ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a211o_1
X_08080_ net550 _02890_ net524 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05292_ top.compVal\[38\] vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__inv_2
XANTENNA__05464__B2 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _03703_ _03704_ _03705_ _03706_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06413__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ top.WB.CPU_DAT_O\[19\] top.cb_syn.h_element\[51\] net367 vssd1 vssd1 vccd1
+ vccd1 _01356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07933_ net420 _04471_ _04472_ net262 vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout198_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ net432 net1565 net253 top.findLeastValue.sum\[25\] _04417_ vssd1 vssd1 vccd1
+ vccd1 _01814_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06815_ _03394_ net126 vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__nand2_1
X_09603_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout365_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07795_ top.hTree.tree_reg\[38\] top.findLeastValue.sum\[38\] net283 vssd1 vssd1
+ vccd1 vccd1 _04362_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ net746 net581 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__and2_1
X_06746_ _03528_ _03529_ _03531_ _03532_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a22o_1
X_09465_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__and2_1
X_06677_ _03462_ _03474_ _03464_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08416_ net1050 _04773_ _04772_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__mux2_1
X_05628_ net1196 net169 _02696_ net210 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09396_ top.hTree.nulls\[58\] net400 net228 vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08347_ top.cb_syn.char_path_n\[31\] net369 net327 top.cb_syn.char_path_n\[29\] net173
+ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a221o_1
X_05559_ _02637_ _02638_ net465 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07796__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08641__A1 top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ top.cb_syn.char_path_n\[65\] net195 _04701_ vssd1 vssd1 vccd1 vccd1 _01684_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_59_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05455__B2 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07229_ top.findLeastValue.val2\[43\] top.findLeastValue.val1\[43\] vssd1 vssd1 vccd1
+ vccd1 _03905_ sky130_fd_sc_hd__nand2_1
X_10240_ net805 net640 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__and2_1
X_10171_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08420__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 net142 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_4
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
Xfanout151 _03506_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_4
Xfanout162 _02805_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_4
Xfanout195 _04615_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07904__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08656__A _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05930__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06875__S net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08880__A1 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ clknet_leaf_23_clk _02175_ _01015_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ clknet_leaf_40_clk _02121_ _00946_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10507_ net754 net589 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11487_ clknet_leaf_93_clk _02052_ _00877_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10438_ net820 net655 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ net758 net593 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07580_ _04178_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nor2_2
X_06600_ top.compVal\[7\] top.compVal\[6\] top.compVal\[5\] top.compVal\[4\] vssd1
+ vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06531_ net1512 _03335_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__xor2_1
X_09250_ _02557_ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nand2_1
X_08201_ top.cb_syn.char_path_n\[104\] net380 net337 top.cb_syn.char_path_n\[102\]
+ net183 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06462_ net1576 net299 _03304_ _03305_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08871__A1 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05413_ top.cb_syn.zeroes\[3\] vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06393_ top.hist_data_o\[20\] top.hist_data_o\[19\] top.hist_data_o\[18\] _03257_
+ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09181_ _02514_ _02835_ top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06882__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__A1 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ net1470 _04625_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__xor2_1
XANTENNA__06814__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05344_ top.findLeastValue.val2\[36\] vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08063_ top.cb_syn.zeroes\[6\] _04572_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__nand2_1
X_07014_ top.findLeastValue.val2\[2\] top.findLeastValue.val2\[1\] top.findLeastValue.val2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout113_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08965_ top.WB.CPU_DAT_O\[3\] net1250 net320 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__mux2_1
X_07916_ top.hTree.tree_reg\[14\] top.findLeastValue.sum\[14\] net267 vssd1 vssd1
+ vccd1 vccd1 _04459_ sky130_fd_sc_hd__mux2_1
X_08896_ net1091 top.WB.CPU_DAT_O\[6\] net305 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__mux2_1
XANTENNA__07898__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ net471 _04402_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ net420 _04347_ _04348_ net262 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__and2_1
X_06729_ top.findLeastValue.val2\[38\] _02409_ top.compVal\[39\] _02459_ vssd1 vssd1
+ vccd1 vccd1 _03527_ sky130_fd_sc_hd__a2bb2o_1
X_09448_ net750 net585 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__and2_1
X_09379_ top.hTree.nulls\[52\] net399 net228 vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08614__A1 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ clknet_leaf_85_clk _01975_ _00800_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ clknet_leaf_77_clk _01906_ _00731_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ clknet_leaf_42_clk _01837_ _00662_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_10223_ net813 net648 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__and2_1
X_10154_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__and2_1
XANTENNA_input43_A gpio_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 top.sram_interface.init_counter\[22\] vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net822 net657 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__and2_1
X_10987_ clknet_leaf_70_clk _01552_ _00377_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06864__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08605__A1 _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ clknet_leaf_22_clk _02158_ _00998_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_96_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold407 top.cb_syn.char_path\[106\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
X_11539_ clknet_leaf_70_clk _02104_ _00929_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold418 top.path\[100\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07813__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold429 top.path\[69\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05962_ top.sram_interface.CB_write_counter\[0\] top.sram_interface.CB_write_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__and2b_1
X_08750_ top.path\[18\] top.path\[19\] net508 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__mux2_1
X_08681_ top.cb_syn.i\[4\] _04881_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__or2_1
X_07701_ top.hTree.tree_reg\[56\] top.findLeastValue.least1\[1\] net281 vssd1 vssd1
+ vccd1 vccd1 _04286_ sky130_fd_sc_hd__mux2_1
XANTENNA__09333__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05893_ net1528 top.WB.CPU_DAT_O\[5\] net349 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XANTENNA__07344__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ net521 _04225_ _04228_ net516 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07563_ top.cb_syn.char_path_n\[34\] top.cb_syn.char_path_n\[33\] top.cb_syn.char_path_n\[36\]
+ top.cb_syn.char_path_n\[35\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux4_1
X_09302_ _05244_ _05245_ net504 vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06514_ top.histogram.total\[28\] _03341_ net1448 vssd1 vssd1 vccd1 vccd1 _03345_
+ sky130_fd_sc_hd__a21oi_1
X_07494_ net342 top.dut.bits_in_buf_next\[0\] _04090_ _04094_ _04095_ vssd1 vssd1
+ vccd1 vccd1 _04096_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout230_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09233_ top.header_synthesis.header\[5\] top.cb_syn.char_index\[5\] net490 vssd1
+ vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__mux2_1
X_06445_ net298 _03267_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout328_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09164_ _04547_ _05162_ _05164_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__or3_1
X_08115_ net412 _02887_ _04178_ net489 _04585_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a221o_1
X_06376_ _03241_ _03240_ _03239_ _03238_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__or4bb_1
X_09095_ _03013_ _05093_ top.sram_interface.word_cnt\[13\] vssd1 vssd1 vccd1 vccd1
+ _05117_ sky130_fd_sc_hd__o21a_1
X_05327_ top.compVal\[2\] vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08046_ _04190_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout697_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ net861 net696 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__and2_1
XANTENNA__05594__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ top.WB.CPU_DAT_O\[20\] net1435 net318 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__mux2_1
X_08879_ net1055 top.WB.CPU_DAT_O\[23\] net303 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__mux2_1
XANTENNA__06138__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ clknet_leaf_25_clk net954 _00300_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ net921 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XANTENNA__05897__A1 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09088__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ clknet_leaf_116_clk _01435_ _00231_ vssd1 vssd1 vccd1 vccd1 top.path\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10772_ clknet_leaf_113_clk _01378_ _00162_ vssd1 vssd1 vccd1 vccd1 top.path\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09749__B net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06846__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11324_ clknet_leaf_89_clk _01889_ _00714_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11255_ clknet_leaf_105_clk _01820_ _00645_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ net822 net657 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__and2_1
X_11186_ clknet_leaf_34_clk _01751_ _00576_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10137_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__and2_1
X_10068_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05888__A1 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08287__C1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06230_ top.hTree.write_HT_fin top.WorR net533 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06161_ top.cb_syn.char_index\[5\] _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__nand2_1
X_06092_ _02972_ _02976_ _02987_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__nor4_1
Xhold226 top.cb_syn.char_path\[70\] vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 top.histogram.sram_out\[4\] vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 top.path\[36\] vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 _01500_ vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 top.cb_syn.char_path\[108\] vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ net871 net706 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__and2_1
Xhold237 top.histogram.sram_out\[22\] vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_1
XANTENNA__07416__A2_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ net864 net699 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__and2_1
Xfanout717 net718 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_2
Xfanout739 net740 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_1
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_1
XANTENNA__05576__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09782_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__and2_1
X_06994_ top.cw1\[3\] net148 _03662_ net486 vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a22o_1
X_08802_ top.path\[64\] net404 net324 top.path\[65\] _02547_ vssd1 vssd1 vccd1 vccd1
+ _04991_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08733_ net430 _04918_ _04920_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__a22o_1
X_05945_ top.compVal\[16\] net161 net146 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout180_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ net496 _04876_ _04874_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a21o_1
X_05876_ net1536 top.WB.CPU_DAT_O\[22\] net350 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
X_08595_ top.cb_syn.char_path_n\[99\] top.cb_syn.char_path_n\[100\] top.cb_syn.char_path_n\[103\]
+ top.cb_syn.char_path_n\[104\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__mux4_1
X_07615_ top.cb_syn.h_element\[60\] top.cb_syn.h_element\[51\] _04176_ vssd1 vssd1
+ vccd1 vccd1 _04214_ sky130_fd_sc_hd__mux2_1
XANTENNA__05879__A1 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ _04144_ _04145_ net290 vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__mux2_1
XANTENNA__06828__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout612_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ _04076_ _04081_ net393 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06428_ top.hist_data_o\[23\] _03259_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06359_ top.cw2\[1\] top.cw2\[0\] vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__or2_1
X_09147_ net457 net361 _02596_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a21oi_1
X_09078_ net455 top.sram_interface.word_cnt\[7\] _02797_ _05104_ vssd1 vssd1 vccd1
+ vccd1 _05105_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_15_Left_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08029_ top.CB_write_complete _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nor2_1
Xhold771 top.cb_syn.zeroes\[3\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 top.findLeastValue.sum\[22\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 top.findLeastValue.wipe_the_char_1 vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 top.cb_syn.char_path_n\[111\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ clknet_leaf_37_clk _01605_ _00430_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05567__B1 _02644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07308__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ net905 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_11873_ clknet_leaf_1_clk top.dut.bits_in_buf_next\[1\] _01245_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bits_in_buf\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_43_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ clknet_leaf_97_clk _01418_ _00214_ vssd1 vssd1 vccd1 vccd1 top.path\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06883__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08284__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ clknet_leaf_10_clk _00050_ _00145_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10686_ clknet_leaf_108_clk _01317_ _00076_ vssd1 vssd1 vccd1 vccd1 top.path\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__A1 top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08992__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ clknet_leaf_43_clk _01872_ _00697_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07795__A1 top.findLeastValue.sum\[38\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11238_ clknet_leaf_67_clk _01803_ _00628_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10153__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05528__A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ clknet_leaf_55_clk _01734_ _00559_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05558__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_42_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05730_ top.histogram.sram_out\[0\] net357 net408 top.hTree.node_reg\[0\] _02781_
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a221o_1
X_05661_ top.cb_syn.char_path\[43\] net529 net310 top.cb_syn.char_path\[107\] vssd1
+ vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
X_08380_ top.cb_syn.char_path_n\[14\] net204 _04752_ vssd1 vssd1 vccd1 vccd1 _01633_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ _02522_ net150 _03662_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a21oi_1
X_05592_ net1211 net168 _02666_ net210 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a22o_1
X_07331_ _03766_ _03980_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__xor2_1
XANTENNA__05730__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07262_ top.findLeastValue.sum\[40\] net278 net272 _03932_ vssd1 vssd1 vccd1 vccd1
+ _01927_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_51_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ top.WB.CPU_DAT_O\[19\] net1486 net365 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
X_06213_ top.cw1\[7\] _03073_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__xor2_1
X_07193_ _03737_ _03866_ _03867_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nand3_1
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08578__A3 top.cb_syn.char_path_n\[96\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06144_ top.sram_interface.init_counter\[3\] _02926_ top.sram_interface.init_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08983__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06075_ _02973_ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nor2_2
X_09903_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__and2_1
Xfanout514 top.cb_syn.curr_state\[8\] vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_2
Xfanout503 top.translation.index\[3\] vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XANTENNA__09852__B net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ net849 net684 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout525 top.cb_syn.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_2
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_60_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout536 top.sram_interface.word_cnt\[5\] vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_2
XANTENNA__05872__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net561 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08749__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 net570 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
X_09765_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__and2_1
X_06977_ top.findLeastValue.histo_index\[6\] _03671_ _03668_ vssd1 vssd1 vccd1 vccd1
+ _03676_ sky130_fd_sc_hd__a21bo_1
X_09696_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__and2_1
X_08716_ _04898_ _04910_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__nor2_1
X_05928_ _02803_ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__or2_2
X_11952__915 vssd1 vssd1 vccd1 vccd1 _11952__915/HI net915 sky130_fd_sc_hd__conb_1
X_08647_ net519 net1037 _04865_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__mux2_1
X_05859_ top.sram_interface.init_counter\[11\] _02876_ vssd1 vssd1 vccd1 vccd1 _02877_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout827_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ top.cb_syn.char_path_n\[91\] top.cb_syn.char_path_n\[92\] top.cb_syn.char_path_n\[95\]
+ top.cb_syn.char_path_n\[96\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__mux4_1
XANTENNA__05721__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07529_ top.cb_syn.char_path_n\[74\] top.cb_syn.char_path_n\[73\] top.cb_syn.char_path_n\[76\]
+ top.cb_syn.char_path_n\[75\] net397 net295 vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__mux4_1
X_10540_ net731 net566 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__and2_1
X_10471_ net830 net665 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__and2_1
XANTENNA__08974__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold590 top.cb_syn.left_check vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11023_ clknet_leaf_62_clk _01588_ _00413_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_11925_ net888 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ clknet_leaf_112_clk _02389_ _01228_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05712__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ clknet_leaf_31_clk _00005_ _00197_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11787_ clknet_leaf_95_clk _02321_ _01159_ vssd1 vssd1 vccd1 vccd1 top.compVal\[36\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06268__B2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ clknet_leaf_5_clk _00028_ _00128_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07560__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ clknet_leaf_98_clk _01300_ _00059_ vssd1 vssd1 vccd1 vccd1 top.path\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08965__A0 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09301__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09953__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ top.findLeastValue.val2\[4\] net129 net120 _03655_ vssd1 vssd1 vccd1 vccd1
+ _02012_ sky130_fd_sc_hd__o22a_1
XANTENNA__09390__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ top.hTree.tree_reg\[21\] top.findLeastValue.sum\[21\] net281 vssd1 vssd1
+ vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
X_06831_ top.compVal\[38\] top.findLeastValue.val1\[38\] net152 vssd1 vssd1 vccd1
+ vccd1 _03621_ sky130_fd_sc_hd__mux2_1
X_09550_ net737 net572 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__and2_1
X_06762_ top.compVal\[19\] _02469_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__and2_1
XANTENNA__07940__A1 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ net1291 top.cb_syn.char_path_n\[58\] net231 vssd1 vssd1 vccd1 vccd1 _01541_
+ sky130_fd_sc_hd__mux2_1
X_09481_ net765 net600 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__and2_1
X_05713_ net1248 net170 _02767_ net209 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__a22o_1
X_08432_ net1119 top.cb_syn.char_path_n\[127\] net230 vssd1 vssd1 vccd1 vccd1 _01610_
+ sky130_fd_sc_hd__mux2_1
X_06693_ _02411_ top.findLeastValue.val1\[36\] top.findLeastValue.val1\[35\] _02412_
+ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__o22a_1
XANTENNA__05703__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05644_ top.histogram.sram_out\[14\] net358 net409 top.hTree.node_reg\[14\] vssd1
+ vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a22o_1
XANTENNA__08248__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ top.cb_syn.char_path_n\[23\] net373 net330 top.cb_syn.char_path_n\[21\] net176
+ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a221o_1
X_05575_ top.cb_syn.char_path\[89\] net537 net532 top.cb_syn.char_path\[57\] vssd1
+ vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a22o_1
X_11912__943 vssd1 vssd1 vccd1 vccd1 net943 _11912__943/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout143_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ top.cb_syn.char_path_n\[57\] net193 _04709_ vssd1 vssd1 vccd1 vccd1 _01676_
+ sky130_fd_sc_hd__o21a_1
X_07314_ net268 _03970_ _03971_ net274 net1676 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__S0 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ _03720_ _03918_ _03919_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout310_A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05867__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__A1 top.findLeastValue.sum\[45\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__A0 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05482__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _03811_ _03850_ _03851_ _03816_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a31oi_2
X_06127_ net444 net453 net447 _03014_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__or4_1
X_06058_ _02530_ top.cb_syn.zero_count\[3\] top.cb_syn.zero_count\[2\] _02531_ vssd1
+ vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__o22a_1
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout777_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout300 _03243_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_4
Xfanout322 _05075_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout333 net335 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
Xfanout366 _05078_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08803__S0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 _04042_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_2
Xfanout377 net386 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_2
X_09817_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__and2_1
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dlymetal6s2s_1
X_09748_ net863 net698 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__and2_1
XANTENNA__07931__A1 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876__879 vssd1 vssd1 vccd1 vccd1 _11876__879/HI net879 sky130_fd_sc_hd__conb_1
XANTENNA__05942__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11710_ clknet_leaf_81_clk _02260_ _01100_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08418__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10249__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ clknet_leaf_109_clk _02191_ _01031_ vssd1 vssd1 vccd1 vccd1 top.path\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_11572_ clknet_leaf_5_clk _02137_ _00962_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ net725 net560 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__and2_1
X_10454_ net803 net638 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__and2_1
XANTENNA__08947__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10385_ net762 net597 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__and2_1
X_11006_ clknet_leaf_52_clk _01571_ _00396_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05933__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ net939 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ clknet_leaf_96_clk _02372_ _01211_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05360_ top.findLeastValue.val2\[5\] vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07989__B2 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05291_ top.compVal\[43\] vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06372__A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05464__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07030_ top.findLeastValue.val1\[2\] top.findLeastValue.val1\[1\] top.findLeastValue.val1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__and3_1
XANTENNA__08938__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ top.WB.CPU_DAT_O\[20\] top.cb_syn.h_element\[52\] net368 vssd1 vssd1 vccd1
+ vccd1 _01357_ sky130_fd_sc_hd__mux2_1
X_07932_ net479 _04470_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__or2_1
XANTENNA__07407__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ net417 _04415_ _04416_ net258 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o211a_1
X_06814_ net287 net125 vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__and2_1
X_09602_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__and2_1
X_07794_ net435 net1610 net249 top.findLeastValue.sum\[39\] _04361_ vssd1 vssd1 vccd1
+ vccd1 _01828_ sky130_fd_sc_hd__a221o_1
X_09533_ net744 net579 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout260_A _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06745_ _02439_ top.findLeastValue.val2\[7\] top.findLeastValue.val2\[6\] _02440_
+ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ net840 net675 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__and2_1
X_06676_ _03459_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__nor2_1
X_08415_ top.cb_syn.h_element\[62\] top.cb_syn.h_element\[53\] net518 vssd1 vssd1
+ vccd1 vccd1 _04773_ sky130_fd_sc_hd__mux2_1
X_05627_ top.hTree.node_reg\[17\] net409 _02694_ _02695_ vssd1 vssd1 vccd1 vccd1 _02696_
+ sky130_fd_sc_hd__a211o_1
X_09395_ net400 _04277_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__nand2_1
XANTENNA__05451__A top.WB.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ top.cb_syn.char_path_n\[31\] net194 _04735_ vssd1 vssd1 vccd1 vccd1 _01650_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07524__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05558_ top.cb_syn.char_path\[60\] net528 net309 top.cb_syn.char_path\[124\] vssd1
+ vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a22o_1
X_08277_ top.cb_syn.char_path_n\[66\] net372 net329 top.cb_syn.char_path_n\[64\] net177
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a221o_1
X_05489_ net487 top.findLeastValue.histo_index\[0\] vssd1 vssd1 vccd1 vccd1 _02574_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05455__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07228_ top.findLeastValue.val2\[43\] top.findLeastValue.val1\[43\] vssd1 vssd1 vccd1
+ vccd1 _03904_ sky130_fd_sc_hd__and2_1
X_07159_ top.findLeastValue.val2\[3\] top.findLeastValue.val1\[3\] vssd1 vssd1 vccd1
+ vccd1 _03835_ sky130_fd_sc_hd__or2_1
XANTENNA__06955__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ net827 net662 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__and2_1
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
Xfanout174 _04616_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout152 net155 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_4
Xfanout163 _02805_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout185 net189 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_1
Xfanout196 net197 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XANTENNA__07904__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08148__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11624_ clknet_leaf_23_clk _02174_ _01014_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06891__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05694__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11555_ clknet_leaf_41_clk _02120_ _00945_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ clknet_leaf_92_clk _02051_ _00876_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[43\]
+ sky130_fd_sc_hd__dfstp_1
X_10506_ net750 net585 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10437_ net820 net655 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__and2_1
XANTENNA__06946__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10299_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__and2_1
XANTENNA__09345__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06530_ _03336_ net1521 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06461_ net299 _03251_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nor2_1
X_05412_ top.cb_syn.zeroes\[4\] vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__inv_2
X_08200_ top.cb_syn.char_path_n\[104\] net201 _04662_ vssd1 vssd1 vccd1 vccd1 _01723_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_16_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08582__A _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05685__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06392_ top.hist_data_o\[17\] top.hist_data_o\[16\] top.hist_data_o\[15\] _03256_
+ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__and4_1
X_09180_ net1699 top.hTree.state\[2\] net254 _05091_ top.hTree.state\[6\] vssd1 vssd1
+ vccd1 vccd1 _00024_ sky130_fd_sc_hd__a32o_1
X_08131_ _04623_ _04624_ _04622_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a21oi_1
X_05343_ top.findLeastValue.val2\[37\] vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__inv_2
X_08062_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__inv_2
XANTENNA__06814__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07013_ top.findLeastValue.val2\[6\] top.findLeastValue.val2\[5\] top.findLeastValue.val2\[4\]
+ top.findLeastValue.val2\[3\] vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08964_ top.WB.CPU_DAT_O\[4\] net1352 net321 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__mux2_1
XANTENNA__06937__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__B1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ top.hTree.tree_reg\[14\] top.findLeastValue.sum\[14\] net285 vssd1 vssd1
+ vccd1 vccd1 _04458_ sky130_fd_sc_hd__mux2_1
XANTENNA__05446__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ net1078 top.WB.CPU_DAT_O\[7\] net305 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__mux2_1
XANTENNA__05880__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ top.findLeastValue.sum\[28\] _04402_ net390 vssd1 vssd1 vccd1 vccd1 _04403_
+ sky130_fd_sc_hd__mux2_1
X_07777_ net479 _04346_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout642_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ net735 net570 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__and2_1
X_06728_ _03523_ _03525_ _03517_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o21a_1
X_09447_ net750 net585 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06659_ _02431_ top.findLeastValue.val1\[20\] _03414_ _03419_ _03456_ vssd1 vssd1
+ vccd1 vccd1 _03457_ sky130_fd_sc_hd__a2111o_1
X_09378_ net398 _04302_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__nand2_1
XANTENNA__05676__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ top.cb_syn.char_path_n\[40\] net380 net337 top.cb_syn.char_path_n\[38\] net183
+ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ clknet_leaf_77_clk _01905_ _00730_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11271_ clknet_leaf_43_clk _01836_ _00661_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10222_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__and2_1
X_10153_ net753 net588 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__and2_1
XANTENNA__06928__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05600__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__B1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 top.sram_interface.init_counter\[13\] vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
X_10084_ net822 net657 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__and2_1
XANTENNA_input36_A gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ clknet_leaf_71_clk _01551_ _00376_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05667__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ clknet_leaf_7_clk _02157_ _00997_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.check
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold408 net79 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
X_11538_ clknet_leaf_69_clk _02103_ _00928_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold419 top.cb_syn.char_path\[107\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ clknet_leaf_103_clk _02034_ _00859_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[26\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06919__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07700_ top.hTree.tree_reg\[56\] _04248_ net388 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__and3_1
X_05961_ top.compVal\[0\] net160 net143 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ _02217_ sky130_fd_sc_hd__a22o_1
XANTENNA__08577__A _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ net1622 _04888_ _04885_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__o21a_1
XANTENNA__07001__A2_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05892_ top.hist_data_o\[6\] top.WB.CPU_DAT_O\[6\] net349 vssd1 vssd1 vccd1 vccd1
+ _02258_ sky130_fd_sc_hd__mux2_1
X_07631_ _04184_ _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07562_ top.cb_syn.char_path_n\[38\] top.cb_syn.char_path_n\[37\] top.cb_syn.char_path_n\[40\]
+ top.cb_syn.char_path_n\[39\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_49_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09097__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ top.histogram.total\[12\] top.histogram.total\[13\] top.histogram.total\[14\]
+ top.histogram.total\[15\] net509 net506 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__mux4_1
X_06513_ net1501 _03342_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07493_ top.dut.bits_in_buf\[1\] top.dut.bits_in_buf_next\[0\] vssd1 vssd1 vccd1
+ vccd1 _04095_ sky130_fd_sc_hd__nor2_1
XANTENNA__05658__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09232_ net1173 _05202_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[4\]
+ sky130_fd_sc_hd__mux2_1
X_06444_ net1058 net298 vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__nand2_1
X_09163_ _04206_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__nor2_1
X_06375_ net460 top.sram_interface.word_cnt\[9\] _02586_ net451 _02862_ vssd1 vssd1
+ vccd1 vccd1 _03241_ sky130_fd_sc_hd__a221o_1
X_08114_ net464 _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout223_A _05253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05326_ top.compVal\[3\] vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__inv_2
X_09094_ net456 top.sram_interface.word_cnt\[2\] net527 net447 _05116_ vssd1 vssd1
+ vccd1 vccd1 _00041_ sky130_fd_sc_hd__a221o_1
XANTENNA__07804__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ net550 _04189_ _04188_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_116_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05875__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout592_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ net861 net696 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__and2_1
X_08947_ top.WB.CPU_DAT_O\[21\] net1419 net318 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__mux2_1
X_08878_ net1190 top.WB.CPU_DAT_O\[24\] net302 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ net435 net1356 net249 top.findLeastValue.sum\[32\] _04389_ vssd1 vssd1 vccd1
+ vccd1 _01821_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_88_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ clknet_leaf_116_clk _01434_ _00230_ vssd1 vssd1 vccd1 vccd1 top.path\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ clknet_leaf_111_clk _01377_ _00161_ vssd1 vssd1 vccd1 vccd1 top.path\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08426__S _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__B _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11323_ clknet_leaf_90_clk _01888_ _00713_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07271__A1 top.findLeastValue.sum\[38\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ clknet_leaf_103_clk net1491 _00644_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10205_ net825 net660 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__and2_1
X_11185_ clknet_leaf_34_clk _01750_ _00575_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10136_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__and2_1
XANTENNA__08771__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10969_ clknet_leaf_55_clk net1122 _00359_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06160_ top.cb_syn.char_index\[4\] top.cb_syn.char_index\[3\] top.cb_syn.char_index\[2\]
+ top.cb_syn.char_index\[1\] vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__and4_1
XANTENNA__07798__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06091_ _02989_ _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__or2_2
XANTENNA__09675__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 top.histogram.sram_out\[20\] vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 top.path\[28\] vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07262__B2 _03932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold227 _01553_ vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 top.path\[15\] vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 top.path\[51\] vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout707 net710 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_2
X_09850_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__and2_1
Xfanout718 net736 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_2
Xfanout729 net736 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_2
X_09781_ net863 net698 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__and2_1
X_06993_ _02508_ net125 net123 _03681_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a2bb2o_1
X_08801_ net426 _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or2_1
X_08732_ top.path\[60\] net404 net324 top.path\[61\] net505 vssd1 vssd1 vccd1 vccd1
+ _04921_ sky130_fd_sc_hd__o221a_1
X_05944_ top.compVal\[17\] net161 net146 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 _02234_ sky130_fd_sc_hd__a22o_1
X_08663_ net499 _04866_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__or2_1
XANTENNA__07415__S net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05875_ net1388 top.WB.CPU_DAT_O\[23\] net350 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__mux2_1
X_08594_ top.cb_syn.char_path_n\[97\] top.cb_syn.char_path_n\[98\] top.cb_syn.char_path_n\[101\]
+ top.cb_syn.char_path_n\[102\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__mux4_1
X_07614_ net1499 _04213_ _04212_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
X_07545_ top.cb_syn.char_path_n\[10\] top.cb_syn.char_path_n\[9\] top.cb_syn.char_path_n\[12\]
+ top.cb_syn.char_path_n\[11\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout340_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06258__C _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08817__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07476_ top.dut.bit_buf\[4\] net42 net713 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__mux2_1
X_09215_ _02963_ _02968_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or3_1
X_06427_ net1353 _03284_ net301 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06358_ _02602_ _03224_ _03223_ net535 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__o211a_1
X_09146_ _05150_ _05152_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__or2_1
XANTENNA__08770__A _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06289_ net545 _03045_ _03159_ _02583_ top.cb_syn.curr_index\[5\] vssd1 vssd1 vccd1
+ vccd1 _03160_ sky130_fd_sc_hd__a32o_1
X_09077_ net458 net545 top.sram_interface.word_cnt\[2\] net446 _02590_ vssd1 vssd1
+ vccd1 vccd1 _05104_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05309_ top.compVal\[26\] vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__inv_2
X_08028_ net514 net463 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nand2_1
Xhold772 top.cb_syn.cb_length\[5\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold750 top.compVal\[21\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 top.compVal\[1\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 top.cb_syn.char_path_n\[63\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 top.compVal\[28\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
X_09979_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__and2_1
XANTENNA__08929__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ net904 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XANTENNA__06449__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11872_ clknet_leaf_1_clk top.dut.bits_in_buf_next\[0\] _01244_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bits_in_buf\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ clknet_leaf_97_clk _01417_ _00213_ vssd1 vssd1 vccd1 vccd1 top.path\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_118_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ clknet_leaf_8_clk _00049_ _00144_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10685_ clknet_leaf_108_clk _01316_ _00075_ vssd1 vssd1 vccd1 vccd1 top.path\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07492__A1 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ clknet_leaf_43_clk _01871_ _00696_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11237_ clknet_leaf_67_clk net1560 _00627_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05528__B net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ clknet_leaf_54_clk _01733_ _00558_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[114\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07547__A2 top.cb_syn.char_path_n\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__and2_1
X_11099_ clknet_leaf_62_clk _01664_ _00489_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_05660_ top.cb_syn.char_path\[11\] net547 net539 top.cb_syn.char_path\[75\] vssd1
+ vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
X_05591_ top.hTree.node_reg\[23\] net410 _02664_ _02665_ vssd1 vssd1 vccd1 vccd1 _02666_
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_109_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07330_ net268 _03982_ _03983_ net274 net1616 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09000_ top.WB.CPU_DAT_O\[20\] net1425 net365 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
X_07261_ _03895_ _03898_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__xor2_2
XANTENNA__09686__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06212_ net1691 net164 _03085_ net208 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a22o_1
X_07192_ _03737_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nand2_1
X_06143_ top.sram_interface.init_counter\[3\] _02926_ vssd1 vssd1 vccd1 vccd1 _03020_
+ sky130_fd_sc_hd__nor2_1
X_06074_ top.cb_syn.i\[2\] top.cb_syn.cb_length\[2\] vssd1 vssd1 vccd1 vccd1 _02974_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_113_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06994__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ net793 net628 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__and2_1
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_2
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07538__A2 top.cb_syn.char_path_n\[88\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09833_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__and2_1
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
Xfanout537 top.sram_interface.word_cnt\[3\] vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_4
Xfanout526 top.sram_interface.word_cnt\[12\] vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
XANTENNA_fanout290_A _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07943__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net849 net684 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__and2_1
X_06976_ top.findLeastValue.histo_index\[7\] _03672_ _03674_ vssd1 vssd1 vccd1 vccd1
+ _01956_ sky130_fd_sc_hd__o21a_1
XANTENNA__05454__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__and2_1
X_08715_ top.header_synthesis.count\[1\] _04896_ _04907_ vssd1 vssd1 vccd1 vccd1 _04910_
+ sky130_fd_sc_hd__o21ai_1
X_05927_ net443 _02553_ _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout555_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ _04196_ _04768_ _04769_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05858_ _02873_ _02874_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _02542_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout722_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05789_ top.sram_interface.zero_cnt\[0\] net456 top.sram_interface.word_cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ top.cb_syn.char_path_n\[78\] top.cb_syn.char_path_n\[77\] top.cb_syn.char_path_n\[80\]
+ top.cb_syn.char_path_n\[79\] net397 net294 vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ _04045_ _04056_ _04066_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a21o_1
X_10470_ net829 net664 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__and2_1
X_09129_ net360 _05122_ _05138_ net1574 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold580 top.histogram.init_edge vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11022_ clknet_leaf_65_clk _01587_ _00412_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[104\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold591 top.hTree.state\[9\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10270__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11924_ net887 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__08585__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__B2 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11855_ clknet_leaf_96_clk _02388_ _01227_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_10806_ clknet_leaf_39_clk _00004_ _00196_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11786_ clknet_leaf_96_clk _02320_ _01158_ vssd1 vssd1 vccd1 vccd1 top.compVal\[35\]
+ sky130_fd_sc_hd__dfrtp_4
X_10737_ clknet_leaf_40_clk _01368_ _00127_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07560__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ clknet_leaf_110_clk _01299_ _00058_ vssd1 vssd1 vccd1 vccd1 top.path\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_10599_ net738 net573 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__and2_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__08569__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ top.findLeastValue.val2\[39\] net128 net119 _03620_ vssd1 vssd1 vccd1 vccd1
+ _02047_ sky130_fd_sc_hd__o22a_1
XANTENNA__05951__A1 top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ _03547_ _03552_ _03554_ _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__a31o_1
XANTENNA__08576__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ net1387 top.cb_syn.char_path_n\[59\] net231 vssd1 vssd1 vccd1 vccd1 _01542_
+ sky130_fd_sc_hd__mux2_1
X_09480_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__and2_1
X_05712_ top.histogram.sram_out\[3\] net357 net408 top.hTree.node_reg\[3\] _02766_
+ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a221o_1
X_06692_ _02408_ top.findLeastValue.val1\[43\] _02481_ top.compVal\[42\] vssd1 vssd1
+ vccd1 vccd1 _03490_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__05951__B2 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05643_ _02707_ _02708_ net468 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__o21a_1
X_08431_ _04586_ _04610_ _04178_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__nor3b_1
XANTENNA__06150__C_N net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06900__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ top.cb_syn.char_path_n\[23\] net195 _04743_ vssd1 vssd1 vccd1 vccd1 _01642_
+ sky130_fd_sc_hd__o21a_1
X_05574_ net1421 net168 _02651_ net210 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a22o_1
X_08293_ top.cb_syn.char_path_n\[58\] net371 net329 top.cb_syn.char_path_n\[56\] net177
+ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a221o_1
X_07313_ _03756_ _03969_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ _03720_ _03918_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout136_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08405__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ _03812_ _03813_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__and2_1
X_06126_ net542 net526 net406 vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__o21ai_1
X_06057_ _02527_ top.cb_syn.zero_count\[6\] _02559_ top.cb_syn.zeroes\[5\] vssd1 vssd1
+ vccd1 vccd1 _02957_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08169__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _03243_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
Xfanout312 _02606_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_4
XANTENNA__07664__A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 _04917_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_4
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
Xfanout356 _02609_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout672_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08803__S1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
Xfanout378 net386 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_2
X_09816_ net843 net678 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__and2_1
Xfanout367 _05077_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_2
XANTENNA__06195__B2 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__and2_1
X_06959_ top.findLeastValue.wipe_the_char_1 net149 _03662_ vssd1 vssd1 vccd1 vccd1
+ _03663_ sky130_fd_sc_hd__a21o_1
XANTENNA__05942__B2 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ net850 net685 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08629_ _04847_ _04848_ net496 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ clknet_leaf_110_clk _02190_ _01030_ vssd1 vssd1 vccd1 vccd1 top.path\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_11571_ clknet_leaf_27_clk _02136_ _00961_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10249__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ net733 net568 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ net809 net644 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__and2_1
X_10384_ net760 net595 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05630__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06889__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ clknet_leaf_52_clk _01570_ _00395_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06186__B2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11894__925 vssd1 vssd1 vccd1 vccd1 net925 _11894__925/LO sky130_fd_sc_hd__conb_1
XANTENNA__05933__B2 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ net938 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XANTENNA__05697__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ clknet_leaf_65_clk _02371_ _01210_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08635__A0 top.cb_syn.char_path_n\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
X_11769_ clknet_leaf_45_clk _02308_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05290_ top.compVal\[44\] vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06949__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ top.WB.CPU_DAT_O\[21\] net1485 net367 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__mux2_1
X_07931_ top.hTree.tree_reg\[11\] top.findLeastValue.sum\[11\] net267 vssd1 vssd1
+ vccd1 vccd1 _04471_ sky130_fd_sc_hd__mux2_1
XANTENNA__08166__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ net475 _04414_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or2_1
X_06813_ _03412_ net149 _03610_ net288 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a211o_1
X_09601_ net741 net576 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__and2_1
X_07793_ net418 _04359_ _04360_ net260 vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__o211a_1
X_09532_ net744 net579 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06744_ _03539_ _03540_ _03541_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__o21bai_1
X_09463_ net836 net671 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__and2_1
X_06675_ _02424_ top.findLeastValue.val1\[28\] top.findLeastValue.val1\[27\] _02425_
+ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__o221a_1
X_08414_ _04769_ _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__nor2_4
X_09394_ net978 net221 _05275_ _05276_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a22o_1
X_05626_ top.histogram.sram_out\[17\] net358 net355 top.hTree.node_reg\[49\] vssd1
+ vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a22o_1
X_05557_ top.cb_syn.char_path\[28\] net546 net537 top.cb_syn.char_path\[92\] vssd1
+ vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
X_08345_ top.cb_syn.char_path_n\[32\] net373 net327 top.cb_syn.char_path_n\[30\] net176
+ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_50_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07524__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05878__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08276_ top.cb_syn.char_path_n\[66\] net196 _04700_ vssd1 vssd1 vccd1 vccd1 _01685_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07659__A _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05488_ net483 net485 net486 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1
+ vccd1 _02573_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07227_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__inv_2
XANTENNA__07378__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__inv_2
X_06109_ _02997_ _03005_ _03007_ _02996_ net1641 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a32o_1
XANTENNA__05612__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07089_ top.findLeastValue.val2\[22\] top.findLeastValue.val1\[22\] vssd1 vssd1 vccd1
+ vccd1 _03765_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_98_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
Xfanout120 net121 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08157__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 _03507_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08788__S0 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_4
Xfanout164 net167 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_2
Xfanout186 net188 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_2
Xfanout175 net177 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_2
Xfanout197 net206 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XANTENNA__07365__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05679__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11623_ clknet_leaf_28_clk _02173_ _01013_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
X_11554_ clknet_leaf_41_clk _02119_ _00944_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11485_ clknet_leaf_91_clk _02050_ _00875_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[42\]
+ sky130_fd_sc_hd__dfstp_1
X_10505_ net750 net585 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10436_ net818 net653 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__and2_1
XANTENNA__09042__A0 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ net758 net593 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__and2_1
X_10298_ net859 net694 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09345__A1 top.hTree.node_reg\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_108_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06460_ top.hist_data_o\[9\] top.hist_data_o\[8\] _03249_ top.hist_data_o\[10\] vssd1
+ vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a31o_1
X_05411_ top.cb_syn.zeroes\[5\] vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_117_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08130_ top.cb_syn.cb_length\[5\] _04611_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_103_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06391_ top.hist_data_o\[14\] _03249_ _03252_ _03254_ vssd1 vssd1 vccd1 vccd1 _03256_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06882__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05342_ top.findLeastValue.val2\[39\] vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08061_ _02528_ _04571_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09033__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07012_ top.findLeastValue.val2\[14\] top.findLeastValue.val2\[13\] top.findLeastValue.val2\[12\]
+ top.findLeastValue.val2\[11\] vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ top.WB.CPU_DAT_O\[5\] net1380 net321 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
X_07914_ net437 net1436 net251 top.findLeastValue.sum\[15\] _04457_ vssd1 vssd1 vccd1
+ vccd1 _01804_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08894_ net1044 top.WB.CPU_DAT_O\[8\] net306 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__mux2_1
XANTENNA__07942__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ top.hTree.tree_reg\[28\] top.findLeastValue.sum\[28\] net282 vssd1 vssd1
+ vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
X_07776_ top.hTree.tree_reg\[42\] top.findLeastValue.sum\[42\] net266 vssd1 vssd1
+ vccd1 vccd1 _04347_ sky130_fd_sc_hd__mux2_1
X_06727_ top.compVal\[37\] _02460_ _03521_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_
+ sky130_fd_sc_hd__a22o_1
X_09515_ net733 net568 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09446_ net750 net585 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__and2_1
X_06658_ _02432_ top.findLeastValue.val1\[17\] top.findLeastValue.val1\[16\] _02433_
+ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a221o_1
X_06589_ top.header_synthesis.write_num_lefts top.header_synthesis.write_char_path
+ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__nor2_1
X_09377_ net1030 net221 _05264_ _05265_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
X_05609_ top.hTree.node_reg\[52\] net354 _02679_ _02680_ vssd1 vssd1 vccd1 vccd1 _02681_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_65_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout802_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ top.cb_syn.char_path_n\[40\] net200 _04726_ vssd1 vssd1 vccd1 vccd1 _01659_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ top.cb_syn.char_path_n\[75\] net383 net341 top.cb_syn.char_path_n\[73\] net186
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09024__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ clknet_leaf_45_clk _01835_ _00660_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_10221_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__and2_1
XANTENNA__08783__C1 top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ net751 net586 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__and2_1
X_10083_ net822 net657 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__and2_1
Xhold9 top.hTree.node_reg\[53\] vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07889__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ clknet_leaf_71_clk _01550_ _00375_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06313__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06313__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ clknet_leaf_0_clk top.dut.bit_buf_next\[13\] _00996_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11537_ clknet_leaf_69_clk _02102_ _00927_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07813__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold409 top.cb_syn.char_path\[42\] vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output97_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ clknet_leaf_103_clk _02033_ _00858_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[25\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ clknet_leaf_90_clk _01964_ _00789_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_10419_ net740 net575 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__and2_1
X_05960_ top.compVal\[1\] net160 net143 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ _02218_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05891_ net1549 top.WB.CPU_DAT_O\[7\] net349 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XANTENNA__06001__A0 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ top.cb_syn.max_index\[4\] _04183_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nand2_1
XANTENNA__06378__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07561_ _04159_ _04160_ net290 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08829__B1 top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09300_ top.histogram.total\[8\] top.histogram.total\[9\] top.histogram.total\[10\]
+ top.histogram.total\[11\] net509 net506 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__mux4_1
X_06512_ net1364 _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__a21o_1
XANTENNA__07701__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06304__B2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07492_ top.dut.bit_buf\[1\] net39 net714 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ top.header_synthesis.header\[4\] top.cb_syn.char_index\[4\] net490 vssd1
+ vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__mux2_1
X_06443_ top.hist_data_o\[16\] _03266_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09162_ net525 _04551_ _04606_ net520 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a22oi_1
X_06374_ net528 net309 net461 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09201__B top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08113_ net489 _04195_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__or3_1
XANTENNA__07804__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05325_ top.compVal\[4\] vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__inv_2
XANTENNA__09006__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07804__B2 top.findLeastValue.sum\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ net526 _05113_ _05115_ net536 vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout216_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08532__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net488 _04555_ _04550_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09995_ net860 net695 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout585_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05594__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ top.WB.CPU_DAT_O\[22\] net1215 net318 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__mux2_1
XANTENNA__08768__A _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ net1337 top.WB.CPU_DAT_O\[25\] net302 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__mux2_1
X_07828_ net418 _04387_ _04388_ net260 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ top.hTree.tree_reg\[45\] top.findLeastValue.sum\[45\] net286 vssd1 vssd1
+ vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
X_10770_ clknet_leaf_111_clk _01376_ _00160_ vssd1 vssd1 vccd1 vccd1 top.path\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06846__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ net801 net636 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__and2_1
XANTENNA__08442__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11322_ clknet_leaf_90_clk _01887_ _00712_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07271__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10273__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11253_ clknet_leaf_106_clk net1494 _00643_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10204_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__and2_1
XANTENNA__08756__C1 _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ clknet_leaf_34_clk _01749_ _00574_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09781__B net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05585__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ net778 net613 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__and2_1
XANTENNA__06897__S net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08617__S _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ clknet_leaf_55_clk net1130 _00358_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10899_ clknet_leaf_33_clk _01471_ _00289_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_enable
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06090_ _02535_ top.cb_syn.i\[3\] vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 top.cb_syn.char_path\[47\] vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 top.hTree.nulls\[53\] vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold228 top.cb_syn.char_path\[14\] vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 top.path\[24\] vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08211__B2 top.cb_syn.char_path_n\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_2
X_08800_ top.path\[66\] top.path\[67\] net510 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__mux2_1
Xfanout719 net736 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05576__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ net862 net697 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__and2_1
X_06992_ top.cw1\[4\] net148 _03662_ net484 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08731_ net426 _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__or2_1
X_05943_ top.compVal\[18\] net158 net145 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 _02235_ sky130_fd_sc_hd__a22o_1
X_08662_ net492 _04874_ _04875_ _04868_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__o22a_1
X_05874_ top.hist_data_o\[24\] top.WB.CPU_DAT_O\[24\] net350 vssd1 vssd1 vccd1 vccd1
+ _02276_ sky130_fd_sc_hd__mux2_1
X_07613_ top.cb_syn.max_index\[7\] _04181_ _04182_ _04187_ vssd1 vssd1 vccd1 vccd1
+ _04213_ sky130_fd_sc_hd__o22a_1
X_08593_ net497 _04812_ _02541_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout166_A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07544_ top.cb_syn.char_path_n\[14\] top.cb_syn.char_path_n\[13\] top.cb_syn.char_path_n\[16\]
+ top.cb_syn.char_path_n\[15\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__mux4_1
XANTENNA__08278__A1 top.cb_syn.char_path_n\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06828__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ net1325 net344 _04045_ _04078_ _04080_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout333_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _02955_ _05191_ _02962_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06426_ top.hist_data_o\[24\] _03260_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_62_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout500_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06357_ top.cw1\[1\] top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__xor2_1
X_09145_ net448 _02860_ _05149_ net544 _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a221o_1
X_06288_ top.cb_syn.char_index\[2\] _03042_ top.cb_syn.char_index\[3\] vssd1 vssd1
+ vccd1 vccd1 _03159_ sky130_fd_sc_hd__a21o_1
X_09076_ _02794_ _05101_ _05102_ net542 vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05308_ top.compVal\[27\] vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__inv_2
X_08027_ top.findLeastValue.alternator_timer\[0\] _03665_ _04540_ _03395_ vssd1 vssd1
+ vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
Xhold762 top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 top.sram_interface.init_counter\[3\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 net45 vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 top.cb_syn.char_path_n\[89\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 top.findLeastValue.sum\[42\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__and2_1
XANTENNA__05567__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _04240_ _04255_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__nand2_1
X_11940_ net903 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__07713__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ clknet_leaf_26_clk top.header_synthesis.next_write_num_lefts _01243_ vssd1
+ vssd1 vccd1 vccd1 top.header_synthesis.write_num_lefts sky130_fd_sc_hd__dfrtp_4
XANTENNA__08437__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ clknet_leaf_111_clk _01416_ _00212_ vssd1 vssd1 vccd1 vccd1 top.path\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10753_ clknet_leaf_12_clk _00048_ _00143_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10684_ clknet_leaf_3_clk _01315_ _00074_ vssd1 vssd1 vccd1 vccd1 top.path\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11305_ clknet_leaf_43_clk _01870_ _00695_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ clknet_leaf_66_clk _01801_ _00626_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11167_ clknet_leaf_54_clk _01732_ _00557_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[113\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05558__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__A3 top.cb_syn.char_path_n\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__and2_1
X_11098_ clknet_leaf_61_clk _01663_ _00488_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[44\]
+ sky130_fd_sc_hd__dfrtp_2
X_10049_ net759 net594 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__and2_1
X_05590_ top.histogram.sram_out\[23\] net359 net354 top.hTree.node_reg\[55\] vssd1
+ vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
XANTENNA__05730__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07260_ net271 _03930_ _03931_ net277 net1791 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a32o_1
XANTENNA__09686__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06211_ _03064_ _03066_ _03069_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__or4_1
X_07191_ top.findLeastValue.val2\[24\] top.findLeastValue.val1\[24\] vssd1 vssd1 vccd1
+ vccd1 _03867_ sky130_fd_sc_hd__or2_1
XANTENNA__05494__B2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06142_ net481 _02877_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06073_ top.cb_syn.cb_length\[2\] top.cb_syn.i\[2\] vssd1 vssd1 vccd1 vccd1 _02973_
+ sky130_fd_sc_hd__and2b_1
X_09901_ net848 net683 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_113_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout505 top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__and2_1
Xfanout516 top.cb_syn.pulse_first_n vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_2
Xfanout538 top.sram_interface.word_cnt\[3\] vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XANTENNA__05549__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_2
X_09763_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__and2_1
Xfanout549 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_2
X_08714_ _04899_ _04909_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A _04249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ top.findLeastValue.histo_index\[8\] _03674_ _03675_ _03673_ vssd1 vssd1 vccd1
+ vccd1 _01957_ sky130_fd_sc_hd__a22o_1
X_09694_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__and2_1
X_05926_ net536 net537 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__nor2_1
XANTENNA__08594__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05857_ top.sram_interface.init_counter\[23\] top.sram_interface.init_counter\[22\]
+ top.sram_interface.init_counter\[21\] top.sram_interface.init_counter\[20\] vssd1
+ vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__or4_1
X_08645_ net519 _04770_ _04864_ net1647 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ top.cb_syn.char_path_n\[89\] top.cb_syn.char_path_n\[90\] top.cb_syn.char_path_n\[93\]
+ top.cb_syn.char_path_n\[94\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ _04119_ _04126_ _04109_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__mux2_1
XANTENNA__05721__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05788_ net456 top.sram_interface.word_cnt\[5\] vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ top.dut.out_valid_next _04057_ _04058_ _04059_ _04065_ vssd1 vssd1 vccd1
+ vccd1 _04066_ sky130_fd_sc_hd__a311o_1
X_06409_ top.hist_data_o\[21\] top.hist_data_o\[20\] _03272_ vssd1 vssd1 vccd1 vccd1
+ _03273_ sky130_fd_sc_hd__and3_1
XANTENNA__05485__B2 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07389_ net272 _04023_ _04024_ net278 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1
+ vccd1 _01892_ sky130_fd_sc_hd__a32o_1
X_09128_ _02417_ _05127_ _05131_ _05137_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_75_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09059_ _02859_ _04257_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold570 _03351_ vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 top.histogram.total\[22\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ clknet_leaf_64_clk _01586_ _00411_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[103\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold592 _00027_ vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10551__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10270__B net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net886 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__08585__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ clknet_leaf_97_clk _02387_ _01226_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_10805_ clknet_leaf_25_clk _00003_ _00195_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05712__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ clknet_leaf_96_clk _02319_ _01157_ vssd1 vssd1 vccd1 vccd1 top.compVal\[34\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08662__B2 _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10736_ clknet_leaf_40_clk _01367_ _00126_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05476__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05476__B2 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ clknet_leaf_110_clk _01298_ _00057_ vssd1 vssd1 vccd1 vccd1 top.path\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_10598_ net743 net578 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__and2_1
XANTENNA__06976__A1 top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__08630__S _02541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ clknet_leaf_43_clk _01784_ _00609_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
X_06760_ top.compVal\[14\] _03557_ _03556_ _03548_ vssd1 vssd1 vccd1 vccd1 _03558_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08576__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05711_ top.hTree.node_reg\[35\] net307 _02765_ net469 vssd1 vssd1 vccd1 vccd1 _02766_
+ sky130_fd_sc_hd__a22o_1
X_06691_ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__inv_2
X_05642_ top.cb_syn.char_path\[14\] net547 net312 top.cb_syn.char_path\[110\] vssd1
+ vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
X_08430_ top.cb_syn.char_index\[0\] _04780_ _04772_ vssd1 vssd1 vccd1 vccd1 _01611_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05703__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ top.cb_syn.char_path_n\[24\] net373 net330 top.cb_syn.char_path_n\[22\] net176
+ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a221o_1
X_05573_ top.hTree.node_reg\[58\] net354 net410 top.hTree.node_reg\[26\] _02650_ vssd1
+ vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a221o_1
X_08292_ top.cb_syn.char_path_n\[58\] net193 _04708_ vssd1 vssd1 vccd1 vccd1 _01677_
+ sky130_fd_sc_hd__o21a_1
X_07312_ _03756_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__or2_1
XANTENNA__08805__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05467__B2 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07243_ top.findLeastValue.val2\[45\] top.findLeastValue.val1\[45\] vssd1 vssd1 vccd1
+ vccd1 _03919_ sky130_fd_sc_hd__xor2_1
XANTENNA__08405__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ _03848_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06125_ net461 top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__or2_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08540__S net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06056_ _02533_ top.cb_syn.zero_count\[0\] top.cb_syn.zero_count\[1\] _02532_ vssd1
+ vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08169__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07664__B _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 net304 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
Xfanout313 net317 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
Xfanout335 net341 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
X_09815_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__and2_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout324 _04917_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
Xfanout346 net348 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
Xfanout379 net382 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_2
Xfanout368 _05077_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout665_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__and2_1
X_06958_ net149 _03609_ net406 vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__and3b_4
X_05909_ net521 _02889_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__nand2_1
X_09677_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__and2_1
XANTENNA__05942__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ top.cb_syn.char_path_n\[51\] top.cb_syn.char_path_n\[52\] top.cb_syn.char_path_n\[55\]
+ top.cb_syn.char_path_n\[56\] net499 net493 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__mux4_1
X_06889_ top.compVal\[9\] top.findLeastValue.val1\[9\] net154 vssd1 vssd1 vccd1 vccd1
+ _03650_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08892__A1 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ net1153 top.cb_syn.char_path_n\[0\] net232 vssd1 vssd1 vccd1 vccd1 _01483_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ clknet_leaf_27_clk _02135_ _00960_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05458__B2 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ net733 net568 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__and2_1
X_10452_ net809 net644 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__and2_1
XANTENNA__08016__A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10383_ net762 net597 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__and2_1
X_11004_ clknet_leaf_52_clk _01569_ _00394_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05933__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ net937 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08883__A1 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06894__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ clknet_leaf_5_clk _02370_ _01209_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_2
X_11768_ clknet_leaf_74_clk _02307_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_10719_ clknet_leaf_104_clk _01350_ _00109_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11699_ clknet_leaf_9_clk _02249_ _01089_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.CB_write_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11942__905 vssd1 vssd1 vccd1 vccd1 _11942__905/HI net905 sky130_fd_sc_hd__conb_1
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ top.hTree.tree_reg\[11\] top.findLeastValue.sum\[11\] net285 vssd1 vssd1
+ vccd1 vccd1 _04470_ sky130_fd_sc_hd__mux2_1
X_07861_ top.hTree.tree_reg\[25\] top.findLeastValue.sum\[25\] net264 vssd1 vssd1
+ vccd1 vccd1 _04415_ sky130_fd_sc_hd__mux2_1
X_07792_ net476 _04358_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__or2_1
X_06812_ _03412_ _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__and2_1
X_09600_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__and2_1
X_09531_ net743 net578 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__and2_1
X_06743_ _02440_ top.findLeastValue.val2\[6\] top.findLeastValue.val2\[5\] _02441_
+ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09462_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__and2_1
XANTENNA__08874__A1 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06674_ _03463_ _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__or2_1
X_05625_ _02692_ _02693_ net468 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__o21a_1
X_08413_ _04767_ _04768_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__or2_1
X_09393_ top.hTree.nulls\[57\] net399 net229 vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08535__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08344_ top.cb_syn.char_path_n\[32\] net193 _04734_ vssd1 vssd1 vccd1 vccd1 _01651_
+ sky130_fd_sc_hd__o21a_1
X_05556_ net1777 net167 _02636_ net213 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08275_ top.cb_syn.char_path_n\[67\] net375 net333 top.cb_syn.char_path_n\[65\] net178
+ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout413_A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05487_ top.WB.curr_state\[2\] top.WB.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _02572_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07226_ _03898_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__nand2_1
X_07157_ _03827_ _03830_ _03832_ _03825_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__o211a_1
X_06108_ top.cb_syn.count\[6\] _03003_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__or2_1
X_07088_ top.findLeastValue.val2\[22\] top.findLeastValue.val1\[22\] vssd1 vssd1 vccd1
+ vccd1 _03764_ sky130_fd_sc_hd__nand2_1
XANTENNA__07414__A2_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06039_ top.sram_interface.init_counter\[5\] top.sram_interface.init_counter\[4\]
+ top.sram_interface.init_counter\[3\] top.sram_interface.init_counter\[2\] vssd1
+ vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__or4_1
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
Xfanout165 net167 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_1
Xfanout132 _03611_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08788__S1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_4
Xfanout143 net144 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
XANTENNA__09354__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout176 net177 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
Xfanout198 net206 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
X_09729_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__and2_1
XANTENNA__07614__S _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06876__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ clknet_leaf_28_clk _02172_ _01012_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11553_ clknet_leaf_42_clk _02118_ _00943_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10504_ net750 net585 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__and2_1
X_11484_ clknet_leaf_92_clk _02049_ _00874_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[41\]
+ sky130_fd_sc_hd__dfstp_1
X_10435_ net820 net655 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10366_ net732 net567 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__and2_1
X_10297_ net859 net694 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__and2_1
XANTENNA__05817__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11902__933 vssd1 vssd1 vccd1 vccd1 net933 _11902__933/LO sky130_fd_sc_hd__conb_1
XFILLER_0_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05410_ top.cb_syn.zeroes\[6\] vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06390_ _03249_ _03252_ _03254_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05341_ top.findLeastValue.val2\[40\] vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__inv_2
X_08060_ top.cb_syn.zeroes\[4\] _04569_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07011_ top.findLeastValue.val2\[10\] top.findLeastValue.val2\[9\] top.findLeastValue.val2\[8\]
+ top.findLeastValue.val2\[7\] vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__and4_1
XANTENNA__08792__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ top.WB.CPU_DAT_O\[6\] net1257 net321 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
X_07913_ net420 _04455_ _04456_ net262 vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o211a_1
XANTENNA__09336__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08893_ net1308 top.WB.CPU_DAT_O\[9\] net305 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout196_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07844_ net434 net1493 net248 top.findLeastValue.sum\[29\] _04401_ vssd1 vssd1 vccd1
+ vccd1 _01818_ sky130_fd_sc_hd__a221o_1
X_07775_ top.hTree.tree_reg\[42\] top.findLeastValue.sum\[42\] net285 vssd1 vssd1
+ vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
X_09514_ net734 net569 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__and2_1
X_06726_ top.compVal\[36\] _02461_ _02462_ top.compVal\[35\] vssd1 vssd1 vccd1 vccd1
+ _03524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06858__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09445_ net742 net577 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__and2_1
X_06657_ _02434_ top.findLeastValue.val1\[15\] _03413_ _03420_ vssd1 vssd1 vccd1 vccd1
+ _03455_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout530_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05608_ top.histogram.sram_out\[20\] net359 net410 top.hTree.node_reg\[20\] vssd1
+ vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XANTENNA__05889__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06588_ top.cb_syn.state8 _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__nand2_2
X_09376_ top.hTree.nulls\[51\] net399 net228 vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__o21a_1
X_08327_ top.cb_syn.char_path_n\[41\] net379 net336 top.cb_syn.char_path_n\[39\] net182
+ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a221o_1
X_05539_ top.cb_syn.char_path\[31\] net546 net538 top.cb_syn.char_path\[95\] vssd1
+ vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ net1792 net203 _04691_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__o21a_1
XANTENNA__09885__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07209_ _03882_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor2_1
X_08189_ top.cb_syn.char_path_n\[110\] net383 net339 top.cb_syn.char_path_n\[108\]
+ net186 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a221o_1
X_10220_ net815 net650 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__and2_1
XANTENNA__05597__B1 _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ net753 net588 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__and2_1
XANTENNA__08783__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ net822 net657 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ clknet_leaf_47_clk net1424 _00374_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ clknet_leaf_120_clk top.dut.bit_buf_next\[12\] _00995_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bit_buf\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ clknet_leaf_68_clk _02101_ _00926_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07519__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07026__B1 _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11467_ clknet_leaf_102_clk _02032_ _00857_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[24\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__08223__C1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11398_ clknet_leaf_90_clk _01963_ _00788_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_10418_ net740 net575 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10349_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__and2_1
XANTENNA__05588__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05890_ top.hist_data_o\[8\] top.WB.CPU_DAT_O\[8\] net352 vssd1 vssd1 vccd1 vccd1
+ _02260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ top.cb_syn.char_path_n\[42\] top.cb_syn.char_path_n\[41\] top.cb_syn.char_path_n\[44\]
+ top.cb_syn.char_path_n\[43\] net395 net293 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_49_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08829__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06511_ top.histogram.total\[31\] top.histogram.total\[30\] _03342_ vssd1 vssd1 vccd1
+ vccd1 _03344_ sky130_fd_sc_hd__and3b_1
X_09230_ net1147 _05201_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[3\]
+ sky130_fd_sc_hd__mux2_1
X_07491_ _04045_ _04092_ _04093_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a21o_1
X_06442_ net1305 _03292_ _03243_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
X_09161_ top.cb_syn.end_check net424 top.cb_syn.curr_state\[5\] vssd1 vssd1 vccd1
+ vccd1 _05162_ sky130_fd_sc_hd__o21a_1
X_06373_ _02416_ top.hist_addr\[0\] _03018_ top.sram_interface.init_counter\[0\] _02417_
+ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a221o_1
X_11948__911 vssd1 vssd1 vccd1 vccd1 _11948__911/HI net911 sky130_fd_sc_hd__conb_1
X_08112_ top.cb_syn.h_element\[54\] net412 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__nor2_1
XANTENNA__07002__B net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05324_ top.compVal\[5\] vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__inv_2
X_09092_ net442 net423 _05114_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__o21ai_1
X_08043_ net515 net514 _02886_ _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout209_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05579__B1 _02654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ net860 net695 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__and2_1
X_08945_ top.WB.CPU_DAT_O\[23\] net1254 net318 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__mux2_1
X_08876_ net1060 top.WB.CPU_DAT_O\[26\] net302 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__mux2_1
X_07827_ net476 _04386_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__or2_1
X_07758_ net433 net1510 net258 _04332_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout745_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06709_ _03412_ net149 net288 vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08296__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ top.hTree.tree_reg\[58\] top.findLeastValue.least1\[3\] net280 vssd1 vssd1
+ vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
X_09428_ net801 net636 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__and2_1
X_09359_ net982 net226 net217 _04339_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07256__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11321_ clknet_leaf_104_clk _01886_ _00711_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[8\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__10554__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11252_ clknet_leaf_103_clk _01817_ _00642_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11183_ clknet_leaf_34_clk _01748_ _00573_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_91_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10203_ net821 net656 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__and2_1
XANTENNA__08756__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A gpio_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__and2_1
X_10065_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__and2_1
XANTENNA__05990__A0 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__B1 top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10967_ clknet_leaf_56_clk _01532_ _00357_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10898_ clknet_leaf_33_clk _01470_ _00288_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07247__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08995__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold207 top.cb_syn.char_path\[96\] vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
X_11519_ clknet_leaf_119_clk _02084_ _00909_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold229 top.histogram.sram_out\[26\] vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 net87 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06222__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ _02507_ net125 net123 _03680_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a2bb2o_1
X_08730_ top.path\[62\] top.path\[63\] net511 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__mux2_1
XANTENNA__05981__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05942_ top.compVal\[19\] net159 net145 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 _02236_ sky130_fd_sc_hd__a22o_1
X_08661_ net492 _04789_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
X_05873_ net1481 top.WB.CPU_DAT_O\[25\] net350 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
X_07612_ _04193_ _04194_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nor3_4
X_08592_ top.cb_syn.char_path_n\[107\] top.cb_syn.char_path_n\[108\] top.cb_syn.char_path_n\[111\]
+ top.cb_syn.char_path_n\[112\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__mux4_1
XANTENNA__08808__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07543_ _04127_ _04142_ _04108_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__mux2_1
XANTENNA__08278__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout159_A _02908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ net342 _04064_ _04079_ _04060_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__o211a_1
X_09213_ _02954_ _05190_ _02957_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__o21bai_1
X_06425_ net1126 _03283_ net301 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06958__A_N net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ net451 _05096_ top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _05151_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08986__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06356_ net406 _03087_ _03203_ _03222_ _02602_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06287_ _02585_ _03055_ _03155_ _03157_ _03154_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__o311a_1
X_09075_ net452 _02916_ _02922_ _02900_ net466 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a32o_1
X_05307_ top.compVal\[28\] vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold730 top.controller.fin_reg\[3\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
X_08026_ top.findLeastValue.alternator_timer\[0\] _02791_ vssd1 vssd1 vccd1 vccd1
+ _04540_ sky130_fd_sc_hd__nor2_1
Xhold752 top.cb_syn.zeroes\[2\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 top.cb_syn.i\[3\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 top.cb_syn.char_path_n\[53\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout695_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 top.cb_syn.char_path_n\[81\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 top.cb_syn.char_path_n\[50\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 top.findLeastValue.sum\[30\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout862_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__and2_1
XANTENNA__07961__A1 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ _05071_ top.cb_syn.max_index\[4\] _05059_ vssd1 vssd1 vccd1 vccd1 _01404_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05972__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08859_ net502 _02811_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11870_ clknet_leaf_112_clk _02403_ _01242_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05724__B1 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ clknet_leaf_97_clk _01415_ _00211_ vssd1 vssd1 vccd1 vccd1 top.path\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10549__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05650__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10752_ clknet_leaf_8_clk _00047_ _00142_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10683_ clknet_leaf_116_clk _01314_ _00073_ vssd1 vssd1 vccd1 vccd1 top.path\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08453__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11304_ clknet_leaf_43_clk _01869_ _00694_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11235_ clknet_leaf_67_clk net1601 _00625_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11166_ clknet_leaf_57_clk _01731_ _00556_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[112\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07401__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ clknet_leaf_61_clk _01662_ _00487_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[43\]
+ sky130_fd_sc_hd__dfrtp_2
X_10117_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__and2_1
X_10048_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 _00040_ vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06002__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05715__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09313__A _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__S0 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06140__B1 _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06210_ _02610_ _03062_ _03083_ net458 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a2bb2o_1
X_07190_ top.findLeastValue.val2\[25\] top.findLeastValue.val1\[25\] vssd1 vssd1 vccd1
+ vccd1 _03866_ sky130_fd_sc_hd__xor2_1
XANTENNA__08968__A0 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06141_ net481 _02877_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__and2_1
X_06072_ _02970_ _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__nand2_1
XANTENNA__09983__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05288__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09900_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_113_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06994__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 top.translation.index\[1\] vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08815__S0 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__and2_1
Xfanout539 net541 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
Xfanout517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
XANTENNA__09393__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout528 net532 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_4
X_09762_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__and2_1
X_06974_ top.findLeastValue.startup _02793_ net288 vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__nor3_2
X_08713_ top.header_synthesis.count\[2\] _04898_ _04907_ vssd1 vssd1 vccd1 vccd1 _04909_
+ sky130_fd_sc_hd__o21ai_1
X_05925_ top.sram_interface.CB_write_counter\[0\] _02903_ _02904_ vssd1 vssd1 vccd1
+ vccd1 _02249_ sky130_fd_sc_hd__o21a_1
X_09693_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout276_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ _04862_ _04863_ top.cb_syn.cb_enable vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or3b_1
X_05856_ top.sram_interface.init_counter\[19\] top.sram_interface.init_counter\[18\]
+ top.sram_interface.init_counter\[17\] top.sram_interface.init_counter\[16\] vssd1
+ vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__or4_1
XANTENNA__05706__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08575_ _04793_ _04794_ net496 vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05751__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05787_ top.sram_interface.zero_cnt\[2\] top.sram_interface.zero_cnt\[1\] vssd1 vssd1
+ vccd1 vccd1 _02816_ sky130_fd_sc_hd__and2b_1
X_07526_ _04122_ _04125_ _04110_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout443_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07457_ _04048_ _04060_ _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__and3_1
XANTENNA__06131__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ top.hist_data_o\[19\] top.hist_data_o\[18\] _03271_ vssd1 vssd1 vccd1 vccd1
+ _03272_ sky130_fd_sc_hd__and3_1
XANTENNA__08959__A0 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07388_ _03840_ _03841_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06339_ top.cw1\[1\] top.cw1\[0\] top.cw1\[2\] vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ _05125_ _05135_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__or3_1
X_09058_ _02859_ _04257_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08009_ top.findLeastValue.least2\[1\] top.findLeastValue.least1\[1\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold560 top.hTree.state\[7\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 top.hTree.state\[5\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ clknet_leaf_64_clk _01585_ _00410_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05926__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold593 top.histogram.total\[24\] vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 top.path\[96\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07934__B2 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05945__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ top.translation.writeBin vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_28_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ clknet_leaf_114_clk _02386_ _01225_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_10804_ clknet_leaf_18_clk _01407_ _00194_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_56_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07545__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05811__D top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11784_ clknet_leaf_96_clk _02318_ _01156_ vssd1 vssd1 vccd1 vccd1 top.compVal\[33\]
+ sky130_fd_sc_hd__dfrtp_2
X_10735_ clknet_leaf_40_clk _01366_ _00125_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06122__B1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ clknet_leaf_106_clk _01297_ _00056_ vssd1 vssd1 vccd1 vccd1 top.path\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ net745 net580 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
X_11218_ clknet_leaf_14_clk _01783_ _00608_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05836__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output72_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ clknet_leaf_35_clk _01714_ _00539_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[95\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__05936__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05710_ _02763_ _02764_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__or2_1
X_06690_ top.compVal\[42\] _02481_ _02482_ top.compVal\[41\] _03487_ vssd1 vssd1 vccd1
+ vccd1 _03488_ sky130_fd_sc_hd__o221a_1
X_05641_ top.cb_syn.char_path\[78\] net540 net531 top.cb_syn.char_path\[46\] vssd1
+ vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
X_08360_ top.cb_syn.char_path_n\[24\] net195 _04742_ vssd1 vssd1 vccd1 vccd1 _01643_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06361__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06900__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08638__C1 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05572_ top.histogram.sram_out\[26\] net359 _02649_ net467 vssd1 vssd1 vccd1 vccd1
+ _02650_ sky130_fd_sc_hd__a22o_1
X_07311_ _03752_ _03956_ _03751_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__a21bo_1
X_08291_ top.cb_syn.char_path_n\[59\] net371 net328 top.cb_syn.char_path_n\[57\] net175
+ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a221o_1
X_07242_ _03915_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09289__S0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07173_ top.findLeastValue.val2\[8\] top.findLeastValue.val1\[8\] vssd1 vssd1 vccd1
+ vccd1 _03849_ sky130_fd_sc_hd__xor2_1
XANTENNA__08405__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06124_ net1018 _02619_ net207 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06967__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06055_ _02527_ top.cb_syn.zero_count\[6\] vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__nand2_1
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
Xfanout314 net317 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
Xfanout336 net338 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
X_09814_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout325 _04917_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_2
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09118__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__and2_1
X_06957_ top.findLeastValue.val1\[0\] net135 net112 net1700 vssd1 vssd1 vccd1 vccd1
+ _01961_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout560_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05908_ net488 net412 vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__or2_1
X_09676_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__and2_1
X_06888_ top.findLeastValue.val2\[10\] net130 net121 _03649_ vssd1 vssd1 vccd1 vccd1
+ _02018_ sky130_fd_sc_hd__o22a_1
X_08627_ top.cb_syn.char_path_n\[49\] top.cb_syn.char_path_n\[50\] top.cb_syn.char_path_n\[53\]
+ top.cb_syn.char_path_n\[54\] net499 net493 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__mux4_1
XANTENNA__08341__B2 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05839_ top.sram_interface.word_cnt\[12\] net533 net536 top.sram_interface.word_cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__or4_2
XANTENNA__09888__A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ net1090 top.cb_syn.char_path_n\[1\] net238 vssd1 vssd1 vccd1 vccd1 _01484_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07509_ _02979_ _04104_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__xnor2_4
X_08489_ net1177 top.cb_syn.char_path_n\[70\] net237 vssd1 vssd1 vccd1 vccd1 _01553_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ net734 net569 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__and2_1
X_10451_ net812 net647 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__and2_1
X_10382_ net769 net604 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__and2_1
XANTENNA__10562__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05630__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 top.path\[80\] vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ clknet_leaf_53_clk _01568_ _00393_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08580__A1 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net875 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_88_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ net936 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XANTENNA__09091__D_N net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05697__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ clknet_leaf_41_clk _02369_ _01208_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11767_ clknet_leaf_76_clk _02306_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10718_ clknet_leaf_41_clk _01349_ _00108_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ clknet_leaf_98_clk _02248_ _01088_ vssd1 vssd1 vccd1 vccd1 top.compVal\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ clknet_leaf_79_clk _01280_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10472__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ top.hTree.tree_reg\[25\] top.findLeastValue.sum\[25\] net281 vssd1 vssd1
+ vccd1 vccd1 _04414_ sky130_fd_sc_hd__mux2_1
X_07791_ top.hTree.tree_reg\[39\] top.findLeastValue.sum\[39\] net266 vssd1 vssd1
+ vccd1 vccd1 _04359_ sky130_fd_sc_hd__mux2_1
X_06811_ _03608_ _03605_ _03516_ top.findLeastValue.val2\[46\] vssd1 vssd1 vccd1 vccd1
+ _03609_ sky130_fd_sc_hd__o2bb2a_2
X_09530_ net744 net579 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__and2_1
X_06742_ top.findLeastValue.val2\[4\] _02442_ top.compVal\[5\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _03540_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_108_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09461_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__and2_1
X_06673_ _03460_ _03461_ _03466_ top.findLeastValue.val1\[26\] _02426_ vssd1 vssd1
+ vccd1 vccd1 _03471_ sky130_fd_sc_hd__o32a_1
X_05624_ top.cb_syn.char_path\[49\] net530 net311 top.cb_syn.char_path\[113\] vssd1
+ vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a22o_1
X_08412_ _04767_ _04768_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__nor2_1
X_09392_ net399 _04282_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05688__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ top.cb_syn.char_path_n\[33\] net371 net328 top.cb_syn.char_path_n\[31\] net175
+ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a221o_1
X_05555_ top.hTree.node_reg\[61\] net356 _02634_ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout141_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08274_ top.cb_syn.char_path_n\[67\] net196 _04699_ vssd1 vssd1 vccd1 vccd1 _01686_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05486_ net2 net414 net362 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 _02372_
+ sky130_fd_sc_hd__o22a_1
X_07225_ _03899_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ top.findLeastValue.val2\[2\] top.findLeastValue.val1\[2\] vssd1 vssd1 vccd1
+ vccd1 _03832_ sky130_fd_sc_hd__or2_1
X_06107_ top.cb_syn.count\[7\] _02996_ _02997_ _03006_ vssd1 vssd1 vccd1 vccd1 _02156_
+ sky130_fd_sc_hd__a22o_1
X_07087_ top.findLeastValue.val2\[23\] top.findLeastValue.val1\[23\] vssd1 vssd1 vccd1
+ vccd1 _03763_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05612__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06038_ top.sram_interface.init_counter\[0\] _02924_ vssd1 vssd1 vccd1 vccd1 _02158_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09339__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__A0 top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout122 _03613_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_4
Xfanout133 net139 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout155 net156 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout144 _02909_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout199 net206 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
Xfanout177 _04616_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout166 net167 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09382__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07365__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__and2_1
X_07989_ net436 net1458 net250 top.findLeastValue.sum\[0\] _04517_ vssd1 vssd1 vccd1
+ vccd1 _01789_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09659_ net846 net681 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__and2_1
XANTENNA__05679__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ clknet_leaf_28_clk _02171_ _01011_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10557__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ clknet_leaf_46_clk _02117_ _00942_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ net730 net565 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__and2_1
X_11483_ clknet_leaf_92_clk _02048_ _00873_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[40\]
+ sky130_fd_sc_hd__dfstp_1
X_10434_ net820 net655 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__and2_1
X_10365_ net720 net555 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05603__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10296_ net859 net694 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07805__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06010__A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07540__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11819_ clknet_leaf_65_clk _02352_ _01191_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05340_ top.findLeastValue.val2\[41\] vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__inv_2
XANTENNA__07816__A0 top.findLeastValue.sum\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ top.cw1\[0\] net140 _03686_ top.findLeastValue.histo_index\[0\] vssd1 vssd1
+ vccd1 vccd1 _01933_ sky130_fd_sc_hd__a22o_1
XANTENNA__09991__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08792__A1 top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08961_ top.WB.CPU_DAT_O\[7\] net1234 net321 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
X_07912_ net479 _04454_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or2_1
X_08892_ net1084 top.WB.CPU_DAT_O\[10\] net306 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__mux2_1
XANTENNA__07715__S _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ net417 _04399_ _04400_ net255 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout189_A _04616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07774_ net437 net1497 net252 top.findLeastValue.sum\[43\] _04345_ vssd1 vssd1 vccd1
+ vccd1 _01832_ sky130_fd_sc_hd__a221o_1
XANTENNA__05743__B top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09513_ net732 net567 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__and2_1
X_06725_ _03520_ _03521_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ net742 net577 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__and2_1
X_06656_ _03452_ _03453_ _03428_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a21oi_1
X_05607_ _02677_ _02678_ net467 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06587_ top.cb_syn.zeroes\[7\] top.cb_syn.zeroes\[6\] _03385_ _03386_ vssd1 vssd1
+ vccd1 vccd1 _03387_ sky130_fd_sc_hd__or4_1
X_09375_ net398 _04307_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__nand2_1
X_08326_ top.cb_syn.char_path_n\[41\] net200 _04725_ vssd1 vssd1 vccd1 vccd1 _01660_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05538_ net441 _02619_ net207 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a21o_1
X_08257_ top.cb_syn.char_path_n\[76\] net383 net339 top.cb_syn.char_path_n\[74\] net186
+ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a221o_1
XANTENNA__09885__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05469_ net10 net416 _02570_ top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 _02389_
+ sky130_fd_sc_hd__a22o_1
X_08188_ top.cb_syn.char_path_n\[110\] net203 _04656_ vssd1 vssd1 vccd1 vccd1 _01729_
+ sky130_fd_sc_hd__o21a_1
X_07208_ top.findLeastValue.val2\[33\] top.findLeastValue.val1\[33\] vssd1 vssd1 vccd1
+ vccd1 _03884_ sky130_fd_sc_hd__nor2_1
X_07139_ _03811_ _03812_ _03814_ _03809_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05918__B _02898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__and2_1
X_10081_ net822 net657 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_58_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10983_ clknet_leaf_47_clk net1386 _00373_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11604_ clknet_leaf_120_clk top.dut.bit_buf_next\[11\] _00994_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bit_buf\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ clknet_leaf_81_clk _02100_ _00925_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11466_ clknet_leaf_76_clk _02031_ _00856_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[23\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__07026__A1 _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417_ net740 net575 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__and2_1
X_11397_ clknet_leaf_90_clk _01962_ _00787_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_10348_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10279_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08526__A1 top.cb_syn.char_path_n\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05844__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06378__C net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06510_ top.histogram.total\[30\] _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__nand2_1
X_07490_ top.dut.out\[2\] net344 _04060_ _04074_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__a22o_1
X_06441_ top.hist_data_o\[17\] _03267_ _03271_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _04557_ _05160_ _05161_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_64_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06372_ net459 _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__nand2_1
X_08111_ net523 _02994_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__and2_1
X_05323_ top.compVal\[6\] vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__inv_2
X_09091_ top.sram_interface.TRN_counter\[2\] top.sram_interface.TRN_counter\[1\] top.sram_interface.TRN_counter\[0\]
+ net452 vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__or4b_1
X_08042_ net524 _02889_ _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_116_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ net832 net667 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__and2_1
X_08944_ top.WB.CPU_DAT_O\[24\] net1389 net322 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__mux2_1
X_08875_ net1114 top.WB.CPU_DAT_O\[27\] net302 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__mux2_1
X_07826_ top.findLeastValue.sum\[32\] _04386_ net391 vssd1 vssd1 vccd1 vccd1 _04387_
+ sky130_fd_sc_hd__mux2_1
X_07757_ _04330_ _04331_ net475 vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout640_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ _03476_ _03498_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__a21oi_1
X_07688_ top.hTree.tree_reg\[58\] _04248_ net389 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06639_ top.compVal\[5\] _02498_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__nor2_1
X_09427_ net747 net582 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__and2_1
X_09358_ net984 net227 net217 _04343_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ top.cb_syn.char_path_n\[50\] net376 net333 top.cb_syn.char_path_n\[48\] net179
+ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07256__B2 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ clknet_leaf_14_clk _01885_ _00710_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05929__A _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ top.histogram.total\[28\] top.histogram.total\[29\] top.histogram.total\[30\]
+ top.histogram.total\[31\] net509 net506 vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10554__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07008__B2 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ clknet_leaf_76_clk _01816_ _00641_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11182_ clknet_leaf_33_clk _01747_ _00572_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_path\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ net825 net660 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_91_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10133_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__and2_1
X_10064_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__and2_1
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10966_ clknet_leaf_56_clk _01531_ _00356_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ clknet_leaf_31_clk _01469_ _00287_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05830__C net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06434__S _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold208 top.path\[11\] vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
X_11518_ clknet_leaf_119_clk _02083_ _00908_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold219 top.cb_syn.char_path\[18\] vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ clknet_leaf_88_clk _02014_ _00839_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06222__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06990_ top.cw1\[5\] net148 _03662_ net483 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__a22o_1
X_05941_ top.compVal\[20\] net159 net145 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 _02237_ sky130_fd_sc_hd__a22o_1
X_08660_ top.cb_syn.char_path_n\[0\] _04789_ _04866_ vssd1 vssd1 vccd1 vccd1 _04874_
+ sky130_fd_sc_hd__o21ba_1
X_05872_ net1509 top.WB.CPU_DAT_O\[26\] net350 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
X_07611_ _04196_ _04197_ _04202_ _04210_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__or4_1
X_08591_ _02542_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_93_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06930__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07542_ _04134_ _04141_ _04109_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__mux2_1
X_07473_ top.dut.bits_in_buf_next\[1\] _04052_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__or2_1
X_09212_ _02529_ top.cb_syn.zero_count\[4\] _02958_ _02959_ _05189_ vssd1 vssd1 vccd1
+ vccd1 _05190_ sky130_fd_sc_hd__o221a_1
X_06424_ _03261_ _03282_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__nor2_1
X_06355_ _02574_ _03087_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__nand2_1
X_09143_ net462 net456 top.sram_interface.word_cnt\[14\] net439 vssd1 vssd1 vccd1
+ vccd1 _05150_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout221_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05306_ top.compVal\[29\] vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06997__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06286_ _02591_ _03050_ _03156_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or3_1
X_09074_ _02796_ _02799_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__nor2_1
Xhold720 top.cw1\[3\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ top.findLeastValue.alternator_timer\[1\] _03665_ _04535_ _04539_ vssd1 vssd1
+ vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
Xhold731 top.cb_syn.num_lefts\[6\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 top.header_synthesis.start vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 top.compVal\[7\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 top.findLeastValue.sum\[33\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 top.cb_syn.char_path_n\[114\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 top.cb_syn.zeroes\[6\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 top.sram_interface.init_counter\[6\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__and2_1
X_08927_ _04228_ _04254_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a21bo_1
X_08858_ net513 _02811_ _05036_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__o21a_1
XANTENNA__07713__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ net435 net1457 net249 top.findLeastValue.sum\[36\] _04373_ vssd1 vssd1 vccd1
+ vccd1 _01825_ sky130_fd_sc_hd__a221o_1
XANTENNA__06921__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ top.path\[2\] top.path\[3\] net510 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ clknet_leaf_97_clk _01414_ _00210_ vssd1 vssd1 vccd1 vccd1 top.path\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10549__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ clknet_leaf_9_clk _00046_ _00141_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08734__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10682_ clknet_leaf_3_clk _01313_ _00072_ vssd1 vssd1 vccd1 vccd1 top.path\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10565__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06988__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ clknet_leaf_0_clk _01868_ _00693_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05660__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ clknet_leaf_82_clk net1590 _00624_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ clknet_leaf_57_clk _01730_ _00555_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[111\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07593__B _04175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11096_ clknet_leaf_62_clk _01661_ _00486_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[42\]
+ sky130_fd_sc_hd__dfrtp_2
X_10116_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__and2_1
X_10047_ net756 net591 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__and2_1
XANTENNA__09154__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__B2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 net53 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold91 net54 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__A1 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ clknet_leaf_41_clk _01514_ _00339_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10459__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__S1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06140_ net1093 net166 _03017_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a21o_1
X_06071_ top.cb_syn.i\[6\] top.cb_syn.cb_length\[6\] vssd1 vssd1 vccd1 vccd1 _02971_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__09983__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05651__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07928__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__S1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09830_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__and2_1
Xfanout518 net520 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
Xfanout507 top.translation.index\[1\] vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_2
X_09761_ net853 net688 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__and2_1
X_06973_ top.findLeastValue.histo_index\[7\] _03672_ _03668_ vssd1 vssd1 vccd1 vccd1
+ _03674_ sky130_fd_sc_hd__a21boi_1
X_08712_ _04900_ _04908_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__nor2_1
X_05924_ top.sram_interface.CB_write_counter\[0\] _02903_ _02905_ _02904_ top.sram_interface.CB_write_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a32o_1
XANTENNA__09145__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05954__B2 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ net869 net704 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__and2_1
XANTENNA__08353__C1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05855_ top.sram_interface.init_counter\[15\] top.sram_interface.init_counter\[14\]
+ top.sram_interface.init_counter\[13\] top.sram_interface.init_counter\[12\] vssd1
+ vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__or4_1
X_08643_ net520 top.cb_syn.curr_state\[5\] _04770_ vssd1 vssd1 vccd1 vccd1 _04863_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout171_A _02621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08574_ top.cb_syn.char_path_n\[83\] top.cb_syn.char_path_n\[84\] top.cb_syn.char_path_n\[87\]
+ top.cb_syn.char_path_n\[88\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05751__B _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05786_ _02815_ _02809_ net1635 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
X_07525_ _04123_ _04124_ net289 vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__mux2_1
XANTENNA__07554__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07456_ _04062_ _04063_ net393 vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__mux2_1
X_06407_ top.hist_data_o\[17\] top.hist_data_o\[16\] _03266_ vssd1 vssd1 vccd1 vccd1
+ _03271_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07387_ _03840_ _03841_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06338_ net407 _03205_ _03203_ _02601_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ top.histogram.eof_n top.histogram.state\[0\] top.histogram.state\[2\] top.histogram.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__or4_1
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06269_ net484 _03089_ net483 vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a21oi_1
X_09057_ _03391_ _04255_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nand2_1
XANTENNA__05642__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08008_ _04528_ net1618 _04522_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold572 _00023_ vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 top.histogram.total\[19\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 top.histogram.total\[30\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap291 _05185_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_1
Xhold583 top.hist_data_o\[11\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05926__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07395__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 _03348_ vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__and2_1
XANTENNA__05945__B2 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ net885 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_87_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ clknet_leaf_112_clk _02385_ _01224_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_10803_ clknet_leaf_18_clk _01406_ _00193_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_56_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07545__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ clknet_leaf_97_clk _02317_ _01155_ vssd1 vssd1 vccd1 vccd1 top.compVal\[32\]
+ sky130_fd_sc_hd__dfrtp_4
X_11933__896 vssd1 vssd1 vccd1 vccd1 _11933__896/HI net896 sky130_fd_sc_hd__conb_1
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08464__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10734_ clknet_leaf_40_clk _01365_ _00124_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_10665_ clknet_leaf_106_clk _01296_ _00055_ vssd1 vssd1 vccd1 vccd1 top.path\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ net797 net632 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__and2_1
XANTENNA__09295__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11217_ clknet_leaf_14_clk _01782_ _00607_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
X_11148_ clknet_leaf_35_clk _01713_ _00538_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[94\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__07386__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05936__B2 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ clknet_leaf_52_clk _01644_ _00469_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08350__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05640_ net1359 net171 _02706_ net211 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a22o_1
X_05571_ _02647_ _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__or2_1
XANTENNA__07536__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_07310_ net268 _03958_ _03968_ net274 net1659 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a32o_1
XANTENNA__08653__A3 _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ top.cb_syn.char_path_n\[59\] net193 _04707_ vssd1 vssd1 vccd1 vccd1 _01678_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07310__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ _03720_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or2_1
XANTENNA__09289__S1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07172_ _03842_ _03846_ _03847_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__o221a_1
XANTENNA__09994__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06123_ net1053 net166 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__and2_1
XANTENNA__05624__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06054_ _02528_ top.cb_syn.zero_count\[5\] top.cb_syn.zero_count\[4\] _02529_ vssd1
+ vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08169__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 _02918_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
X_09813_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__and2_1
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout348 _02915_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_2
Xfanout315 net317 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout386_A _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_4
X_09744_ net856 net691 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__and2_1
X_06956_ top.findLeastValue.val1\[1\] net135 net112 net1712 vssd1 vssd1 vccd1 vccd1
+ _01962_ sky130_fd_sc_hd__o22a_1
X_09675_ net788 net623 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__and2_1
X_05907_ net488 net412 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__nor2_1
XANTENNA__05762__A _02564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ top.compVal\[10\] top.findLeastValue.val1\[10\] net154 vssd1 vssd1 vccd1
+ vccd1 _03649_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout553_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _04844_ _04845_ _02542_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05838_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__inv_2
XANTENNA__09888__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
X_08557_ net1409 top.cb_syn.char_path_n\[2\] net232 vssd1 vssd1 vccd1 vccd1 _01485_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05769_ top.compVal\[39\] net162 net147 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ _02324_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout720_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07508_ _02988_ _04105_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__xnor2_2
X_08488_ net1347 top.cb_syn.char_path_n\[71\] net239 vssd1 vssd1 vccd1 vccd1 _01554_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06593__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07439_ net342 vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf_next\[1\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ net810 net645 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__and2_1
X_09109_ top.histogram.out_of_init top.histogram.eof_n _02561_ _05124_ vssd1 vssd1
+ vccd1 vccd1 _05127_ sky130_fd_sc_hd__and4b_1
X_10381_ net769 net604 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10562__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 top.hTree.nulls\[47\] vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11002_ clknet_leaf_54_clk _01567_ _00392_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[84\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold391 top.cb_syn.char_path\[25\] vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_2
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_88_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11904_ net935 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_25_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
X_11835_ clknet_leaf_41_clk _02368_ _01207_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06894__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ clknet_leaf_72_clk _02305_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10717_ clknet_leaf_41_clk _01348_ _00107_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07843__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09045__A0 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11697_ clknet_leaf_110_clk _02247_ _01087_ vssd1 vssd1 vccd1 vccd1 top.compVal\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10648_ clknet_leaf_103_clk _01279_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10579_ net862 net697 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05606__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06442__S _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ top.hTree.tree_reg\[39\] top.findLeastValue.sum\[39\] net283 vssd1 vssd1
+ vccd1 vccd1 _04358_ sky130_fd_sc_hd__mux2_1
X_06810_ _03510_ _03511_ _03513_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__and4b_1
X_06741_ top.compVal\[3\] _02478_ _03536_ _03537_ _03538_ vssd1 vssd1 vccd1 vccd1
+ _03539_ sky130_fd_sc_hd__o221a_1
X_09460_ net732 net567 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__and2_1
XANTENNA__09989__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08411_ net519 net524 _04583_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__o21bai_2
XANTENNA__06960__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06334__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06672_ _03461_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__nand2_1
X_05623_ top.cb_syn.char_path\[17\] net547 net539 top.cb_syn.char_path\[81\] vssd1
+ vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
X_09391_ net1019 net221 _05273_ _05274_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_16_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_08342_ top.cb_syn.char_path_n\[33\] net195 _04733_ vssd1 vssd1 vccd1 vccd1 _01652_
+ sky130_fd_sc_hd__o21a_1
X_05554_ top.histogram.sram_out\[29\] net360 net411 top.hTree.node_reg\[29\] vssd1
+ vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08273_ top.cb_syn.char_path_n\[68\] net375 net333 top.cb_syn.char_path_n\[66\] net178
+ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a221o_1
XANTENNA__07834__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05485_ net13 net415 net364 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 _02373_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout134_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ top.findLeastValue.val2\[41\] top.findLeastValue.val1\[41\] vssd1 vssd1 vccd1
+ vccd1 _03900_ sky130_fd_sc_hd__nand2_1
XANTENNA__09036__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout301_A _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06106_ top.cb_syn.count\[7\] _03005_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__xnor2_1
X_07086_ _03739_ _03757_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__o21a_1
XANTENNA__08795__C1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06037_ _02925_ _02939_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__nor2_1
Xfanout112 net113 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
XANTENNA__08011__A1 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout123 _03612_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
Xfanout134 net139 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_2
Xfanout156 _03506_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
XANTENNA_fanout670_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
Xfanout189 _04616_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
XANTENNA_fanout768_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ net419 _04515_ _04516_ net261 vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o211a_1
Xfanout167 _02621_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net851 net686 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__and2_1
X_06939_ top.findLeastValue.val1\[18\] net138 net116 top.compVal\[18\] vssd1 vssd1
+ vccd1 vccd1 _01979_ sky130_fd_sc_hd__o22a_1
X_09658_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__and2_1
XANTENNA__07911__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ net496 _04828_ _02541_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_83_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09589_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__and2_1
XANTENNA__06876__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ clknet_leaf_28_clk _02170_ _01010_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11551_ clknet_leaf_46_clk _02116_ _00941_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10557__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09027__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10502_ net734 net569 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__and2_1
X_11482_ clknet_leaf_95_clk _02047_ _00872_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[39\]
+ sky130_fd_sc_hd__dfstp_1
X_10433_ net823 net658 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__and2_1
XANTENNA__08786__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ net718 net553 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07882__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10295_ net861 net696 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__and2_1
Xfanout690 net694 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08917__S _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07821__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ clknet_leaf_66_clk _02351_ _01190_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08608__A3 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11749_ clknet_leaf_106_clk _00019_ _01139_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08652__S top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08777__C1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06252__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09991__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ top.WB.CPU_DAT_O\[8\] net1146 net320 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
X_07911_ top.findLeastValue.sum\[15\] _04454_ net391 vssd1 vssd1 vccd1 vccd1 _04455_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07792__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net1159 top.WB.CPU_DAT_O\[11\] net305 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__mux2_1
X_07842_ net470 _04398_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or2_1
X_07773_ net422 _04343_ _04344_ net262 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__o211a_1
X_09512_ net752 net587 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06724_ top.compVal\[35\] _02462_ _02463_ top.compVal\[34\] vssd1 vssd1 vccd1 vccd1
+ _03522_ sky130_fd_sc_hd__o22a_1
XANTENNA__06858__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net726 net561 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__and2_1
X_06655_ top.compVal\[14\] _02494_ _02495_ top.compVal\[13\] vssd1 vssd1 vccd1 vccd1
+ _03453_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout251_A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05606_ top.cb_syn.char_path\[52\] net530 net311 top.cb_syn.char_path\[116\] vssd1
+ vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
X_09374_ net1038 net222 _05262_ _05263_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout349_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06586_ top.cb_syn.zeroes\[1\] top.cb_syn.zeroes\[0\] vssd1 vssd1 vccd1 vccd1 _03386_
+ sky130_fd_sc_hd__or2_1
X_08325_ top.cb_syn.char_path_n\[42\] net379 net336 top.cb_syn.char_path_n\[40\] net182
+ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05537_ net1026 net169 net211 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a21o_1
X_08256_ net1741 net203 _04690_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_104_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05468_ net11 net416 net364 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 _02390_
+ sky130_fd_sc_hd__a22o_1
X_08187_ top.cb_syn.char_path_n\[111\] net383 net339 top.cb_syn.char_path_n\[109\]
+ net186 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10393__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07207_ top.findLeastValue.val2\[33\] top.findLeastValue.val1\[33\] vssd1 vssd1 vccd1
+ vccd1 _03883_ sky130_fd_sc_hd__nand2_1
XANTENNA__08232__A1 top.cb_syn.char_path_n\[88\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05399_ top.findLeastValue.least2\[5\] vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__inv_2
X_07138_ _02476_ _02497_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05597__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ top.findLeastValue.val2\[29\] top.findLeastValue.val1\[29\] vssd1 vssd1 vccd1
+ vccd1 _03745_ sky130_fd_sc_hd__or2_1
XANTENNA__07906__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ net757 net592 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10982_ clknet_leaf_42_clk _01547_ _00372_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07641__S _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ clknet_leaf_5_clk top.dut.bit_buf_next\[10\] _00993_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08472__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__A1 top.cb_syn.char_path_n\[88\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ clknet_leaf_68_clk _02099_ _00924_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07877__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ clknet_leaf_76_clk _02030_ _00855_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ net737 net572 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__and2_1
X_11396_ clknet_leaf_90_clk _01961_ _00786_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10347_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__and2_1
XANTENNA__05588__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__and2_1
XANTENNA__07816__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05860__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06440_ net1140 _03291_ net300 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06371_ _02512_ _02600_ _02603_ _02513_ _03236_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ _04590_ _04589_ top.cb_syn.num_lefts\[0\] vssd1 vssd1 vccd1 vccd1 _01755_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08462__A1 top.cb_syn.char_path_n\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09090_ top.sram_interface.CB_write_counter\[1\] top.sram_interface.CB_write_counter\[0\]
+ net460 _05107_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05322_ top.compVal\[7\] vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__inv_2
X_08041_ net550 _02894_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08214__A1 top.cb_syn.char_path_n\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05579__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ net832 net667 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__and2_1
X_08943_ top.WB.CPU_DAT_O\[25\] net1374 net322 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout299_A _03244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ net1156 top.WB.CPU_DAT_O\[28\] net303 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__mux2_1
XANTENNA__09190__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_A top.controller.state_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ top.hTree.tree_reg\[32\] top.findLeastValue.sum\[32\] net283 vssd1 vssd1
+ vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_1
X_07756_ top.hTree.tree_reg\[46\] top.findLeastValue.least2\[0\] net264 vssd1 vssd1
+ vccd1 vccd1 _04331_ sky130_fd_sc_hd__mux2_1
X_06707_ _03503_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ net257 _04273_ _04274_ net1195 net432 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a32o_1
X_09426_ net747 net582 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06638_ _02442_ top.findLeastValue.val1\[4\] vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__and2_1
X_09357_ net1015 net225 net217 _04347_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout800_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06569_ _03365_ _03369_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__nand2_1
X_08308_ net1747 net196 _04716_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__o21a_1
X_09288_ net504 _05228_ _05230_ _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07256__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08239_ top.cb_syn.char_path_n\[85\] net378 net334 top.cb_syn.char_path_n\[83\] net180
+ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a221o_1
XANTENNA__05929__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ clknet_leaf_75_clk net1547 _00640_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11181_ clknet_leaf_33_clk _01746_ _00571_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10201_ net754 net589 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__and2_1
XANTENNA_hold678_A top.hTree.node_reg\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold845_A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__and2_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08467__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10965_ clknet_leaf_56_clk _01530_ _00355_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ clknet_leaf_31_clk _01468_ _00286_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ clknet_leaf_118_clk _02082_ _00907_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold209 top.hTree.tree_reg\[62\] vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ clknet_leaf_89_clk _02013_ _00838_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ clknet_leaf_17_clk _01944_ _00769_ vssd1 vssd1 vccd1 vccd1 top.cw2\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07546__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05940_ top.compVal\[21\] net158 net145 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 _02238_ sky130_fd_sc_hd__a22o_1
X_05871_ net1774 top.WB.CPU_DAT_O\[27\] net350 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08590_ top.cb_syn.char_path_n\[105\] top.cb_syn.char_path_n\[106\] top.cb_syn.char_path_n\[109\]
+ top.cb_syn.char_path_n\[110\] net500 net494 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__mux4_1
X_07610_ _04205_ _04207_ _04209_ _04203_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__or4b_1
XFILLER_0_72_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07541_ _04137_ _04140_ _04110_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07472_ _04055_ _04077_ _04048_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ _02956_ _02964_ _02961_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a21o_1
X_06423_ top.hist_data_o\[24\] _03260_ top.hist_data_o\[25\] vssd1 vssd1 vccd1 vccd1
+ _03282_ sky130_fd_sc_hd__a21oi_1
X_06354_ net1261 net165 _03221_ net208 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a22o_1
X_09142_ _02840_ _03390_ _05148_ _02845_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a2bb2o_1
X_05305_ top.compVal\[30\] vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__inv_2
X_06285_ net445 top.TRN_char_index\[1\] top.TRN_char_index\[3\] vssd1 vssd1 vccd1
+ vccd1 _03156_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout214_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ net457 net1040 _05100_ net1237 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold710 top.cb_syn.num_lefts\[5\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 top.hTree.nullSumIndex\[0\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08024_ _02784_ _03395_ _04531_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_77_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold743 top.findLeastValue.histo_index\[5\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 top.findLeastValue.sum\[39\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 top.findLeastValue.sum\[31\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 top.cb_syn.char_path_n\[119\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold776 top.findLeastValue.sum\[43\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__and2_1
XANTENNA__09148__C1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ _04254_ _05060_ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or3b_1
X_08857_ top.translation.index\[4\] _05042_ _05040_ vssd1 vssd1 vccd1 vccd1 _01446_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout750_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ net418 _04371_ _04372_ net260 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o211a_1
X_08788_ top.path\[4\] top.path\[5\] top.path\[6\] top.path\[7\] net510 net507 vssd1
+ vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__mux4_1
XANTENNA__05724__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06596__A _02562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ _02518_ net389 _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__o21a_1
X_10750_ clknet_leaf_13_clk _00045_ _00140_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_43_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09409_ top.hTree.nulls\[63\] _02851_ net220 _05285_ vssd1 vssd1 vccd1 vccd1 _05286_
+ sky130_fd_sc_hd__a211o_1
X_10681_ clknet_leaf_3_clk _01312_ _00071_ vssd1 vssd1 vccd1 vccd1 top.path\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10565__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06988__B2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302_ clknet_leaf_2_clk _01867_ _00692_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11233_ clknet_leaf_82_clk _01798_ _00623_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11164_ clknet_leaf_59_clk _01729_ _00554_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08051__A top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07401__A2 _03611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ clknet_leaf_62_clk _01660_ _00485_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07412__A2_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10115_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__and2_1
X_11938__901 vssd1 vssd1 vccd1 vccd1 _11938__901/HI net901 sky130_fd_sc_hd__conb_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10046_ net811 net646 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__and2_1
Xhold81 net50 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 net51 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 top.hTree.node_reg\[15\] vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05715__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ clknet_leaf_39_clk _01513_ _00338_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05479__B2 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06140__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ clknet_leaf_24_clk top.header_synthesis.next_header\[1\] _00269_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06070_ top.cb_syn.cb_length\[6\] top.cb_syn.i\[6\] vssd1 vssd1 vccd1 vccd1 _02970_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_1 ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05651__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
Xfanout508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_4
X_09760_ net852 net687 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06972_ _02501_ _02502_ _02503_ _03669_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__nor4_1
X_09691_ net868 net703 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__and2_1
X_08711_ top.header_synthesis.count\[3\] _04899_ _04907_ vssd1 vssd1 vccd1 vccd1 _04908_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_72_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05923_ top.sram_interface.CB_write_counter\[1\] _02587_ vssd1 vssd1 vccd1 vccd1
+ _02905_ sky130_fd_sc_hd__nor2_1
X_08642_ _04792_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and2b_1
X_11878__881 vssd1 vssd1 vccd1 vccd1 _11878__881/HI net881 sky130_fd_sc_hd__conb_1
XANTENNA__05706__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05854_ _02870_ _02867_ top.sram_interface.counter_HTREE\[0\] vssd1 vssd1 vccd1 vccd1
+ _02287_ sky130_fd_sc_hd__mux2_1
X_08573_ top.cb_syn.char_path_n\[81\] top.cb_syn.char_path_n\[82\] top.cb_syn.char_path_n\[85\]
+ top.cb_syn.char_path_n\[86\] net501 net495 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05785_ _02809_ _02814_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout164_A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07524_ top.cb_syn.char_path_n\[114\] top.cb_syn.char_path_n\[113\] top.cb_syn.char_path_n\[116\]
+ top.cb_syn.char_path_n\[115\] net396 net294 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__mux4_1
XANTENNA__09520__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ top.dut.bit_buf\[11\] top.dut.bit_buf\[4\] net713 vssd1 vssd1 vccd1 vccd1
+ _04063_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout331_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ net1429 _03270_ net301 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07386_ net271 _04018_ _04022_ net278 top.findLeastValue.sum\[6\] vssd1 vssd1 vccd1
+ vccd1 _01893_ sky130_fd_sc_hd__a32o_1
X_06337_ _03088_ _03204_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__nor2_1
XANTENNA__05890__A1 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09125_ top.histogram.state\[7\] top.histogram.state\[3\] top.histogram.state\[5\]
+ top.histogram.state\[6\] vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09056_ net463 _05088_ net954 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a21o_1
X_06268_ net1233 net164 _03139_ net207 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07694__B _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ top.findLeastValue.least2\[2\] top.findLeastValue.least1\[2\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout798_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 top.cb_syn.char_path\[78\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05495__A top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07919__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06199_ top.cw1\[6\] _03072_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__and2_1
Xhold540 _01819_ vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 top.histogram.total\[18\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 top.hist_data_o\[28\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 top.hTree.tree_reg\[40\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 top.hTree.tree_reg\[26\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
X_09958_ net770 net605 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__and2_1
XANTENNA__07395__B2 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _02835_ _05050_ top.findLeastValue.least2\[8\] vssd1 vssd1 vccd1 vccd1 _05056_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__05945__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net875 net710 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__and2_1
X_11920_ net951 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__08895__A1 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ clknet_leaf_96_clk _02384_ _01223_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_10802_ clknet_leaf_20_clk _01405_ _00192_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ clknet_leaf_2_clk _02316_ _01154_ vssd1 vssd1 vccd1 vccd1 top.translation.write_fin
+ sky130_fd_sc_hd__dfrtp_1
X_10733_ clknet_leaf_17_clk _01364_ _00123_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10295__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ clknet_leaf_106_clk _01295_ _00054_ vssd1 vssd1 vccd1 vccd1 top.path\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05881__A1 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10595_ net797 net632 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06830__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216_ clknet_leaf_15_clk _01781_ _00606_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07386__A1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
X_11147_ clknet_leaf_34_clk _01712_ _00537_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[93\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__05936__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11078_ clknet_leaf_52_clk _01643_ _00468_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_10029_ net839 net674 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__and2_1
XANTENNA__08886__A1 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08638__A1 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05570_ top.cb_syn.char_path\[58\] net532 net309 top.cb_syn.char_path\[122\] vssd1
+ vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XANTENNA__07310__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07240_ top.findLeastValue.val2\[44\] top.findLeastValue.val1\[44\] vssd1 vssd1 vccd1
+ vccd1 _03916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05872__A1 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07171_ top.findLeastValue.val2\[6\] top.findLeastValue.val1\[6\] vssd1 vssd1 vccd1
+ vccd1 _03847_ sky130_fd_sc_hd__or2_1
XANTENNA__09994__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06122_ net1434 _02619_ net207 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a21o_1
XANTENNA__06903__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06053_ top.cb_syn.count\[7\] _02526_ _02527_ top.cb_syn.count\[6\] _02952_ vssd1
+ vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
Xfanout327 net331 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
Xfanout338 net341 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
X_09812_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__and2_1
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
Xfanout349 net352 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout379_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ top.findLeastValue.val1\[2\] net135 net112 net1651 vssd1 vssd1 vccd1 vccd1
+ _01963_ sky130_fd_sc_hd__o22a_1
X_05906_ top.cb_syn.end_check top.cb_syn.curr_state\[5\] vssd1 vssd1 vccd1 vccd1 _02888_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__05762__B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08877__A1 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06886_ top.findLeastValue.val2\[11\] net131 net120 _03648_ vssd1 vssd1 vccd1 vccd1
+ _02019_ sky130_fd_sc_hd__o22a_1
X_09674_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__and2_1
X_08625_ top.cb_syn.char_path_n\[57\] top.cb_syn.char_path_n\[58\] top.cb_syn.char_path_n\[61\]
+ top.cb_syn.char_path_n\[62\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__mux4_1
X_05837_ top.WorR _02553_ _02844_ _02847_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__or4_1
XANTENNA__06888__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ net1182 top.cb_syn.char_path_n\[3\] net237 vssd1 vssd1 vccd1 vccd1 _01486_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06352__A2 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _02972_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_85_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05560__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05768_ top.compVal\[40\] net163 _02806_ top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1
+ vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08487_ net1309 top.cb_syn.char_path_n\[72\] net239 vssd1 vssd1 vccd1 vccd1 _01555_
+ sky130_fd_sc_hd__mux2_1
X_05699_ top.histogram.sram_out\[5\] net357 net409 top.hTree.node_reg\[5\] vssd1 vssd1
+ vccd1 vccd1 _02756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07438_ _04043_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09054__A1 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07369_ _03810_ _04009_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nand2_1
X_09108_ net453 _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__nand2_1
X_10380_ net769 net604 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09039_ top.WB.CPU_DAT_O\[11\] net1259 net315 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
Xhold370 top.cb_syn.char_path\[10\] vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 top.path\[41\] vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09357__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ clknet_leaf_53_clk _01566_ _00391_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[83\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold392 top.path\[32\] vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout850 net854 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_2
Xfanout861 net865 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_2
Xfanout872 net875 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11903_ net934 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05551__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11834_ clknet_leaf_42_clk _02367_ _01206_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
X_11765_ clknet_leaf_72_clk _02304_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07828__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10716_ clknet_leaf_42_clk _01347_ _00106_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_11696_ clknet_leaf_98_clk _02246_ _01086_ vssd1 vssd1 vccd1 vccd1 top.compVal\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ clknet_leaf_103_clk _01278_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10578_ net727 net562 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__and2_1
XANTENNA__09348__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _02442_ top.findLeastValue.val2\[4\] vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06671_ top.compVal\[26\] _02491_ _03466_ _03467_ _03468_ vssd1 vssd1 vccd1 vccd1
+ _03469_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_108_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08410_ net488 net519 net424 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a21o_1
X_05622_ net1452 net169 _02691_ net210 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a22o_1
XANTENNA__09989__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05542__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09390_ top.hTree.nulls\[56\] net399 net228 vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__o21a_1
X_05553_ _02632_ _02633_ net465 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__o21a_1
X_08341_ top.cb_syn.char_path_n\[34\] net372 net329 top.cb_syn.char_path_n\[32\] net177
+ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ top.cb_syn.char_path_n\[68\] net196 _04698_ vssd1 vssd1 vccd1 vccd1 _01687_
+ sky130_fd_sc_hd__o21a_1
X_05484_ net24 net416 _02570_ top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 _02374_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07223_ top.findLeastValue.val2\[41\] top.findLeastValue.val1\[41\] vssd1 vssd1 vccd1
+ vccd1 _03899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_A _03611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07154_ top.findLeastValue.val2\[0\] top.findLeastValue.val1\[0\] _03828_ vssd1 vssd1
+ vccd1 vccd1 _03830_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06105_ top.cb_syn.count\[6\] _03003_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__nand2_1
X_07085_ _03751_ _03754_ _03755_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08795__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06036_ top.sram_interface.init_counter\[0\] _02924_ top.sram_interface.init_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09339__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
Xfanout124 _03612_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_1
Xfanout146 _02909_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net138 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
Xfanout179 net189 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
Xfanout168 net170 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
Xfanout157 _03017_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_4
X_07987_ net477 _04514_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__or2_1
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__and2_1
XANTENNA__07770__A1 top.findLeastValue.sum\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ top.findLeastValue.val1\[19\] net138 net115 top.compVal\[19\] vssd1 vssd1
+ vccd1 vccd1 _01980_ sky130_fd_sc_hd__o22a_1
X_09657_ net789 net624 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout830_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06869_ top.compVal\[19\] top.findLeastValue.val1\[19\] net152 vssd1 vssd1 vccd1
+ vccd1 _03640_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ top.cb_syn.char_path_n\[27\] top.cb_syn.char_path_n\[28\] top.cb_syn.char_path_n\[31\]
+ top.cb_syn.char_path_n\[32\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__mux4_1
X_09588_ net798 net633 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__and2_1
X_08539_ net1220 top.cb_syn.char_path_n\[20\] net235 vssd1 vssd1 vccd1 vccd1 _01503_
+ sky130_fd_sc_hd__mux2_1
X_11550_ clknet_leaf_45_clk _02115_ _00940_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07286__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ net734 net569 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__and2_1
X_11481_ clknet_leaf_95_clk _02046_ _00871_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[38\]
+ sky130_fd_sc_hd__dfstp_1
X_10432_ net822 net657 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__and2_1
XANTENNA__08250__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10363_ net718 net553 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__and2_1
X_10294_ net829 net664 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net693 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_2
Xfanout680 net712 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05772__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ clknet_leaf_66_clk _02350_ _01189_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07403__A _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07277__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ clknet_leaf_106_clk _00017_ _01138_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ clknet_leaf_86_clk _02229_ _01069_ vssd1 vssd1 vccd1 vccd1 top.compVal\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07549__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08624__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07910_ top.hTree.tree_reg\[15\] top.findLeastValue.sum\[15\] net286 vssd1 vssd1
+ vccd1 vccd1 _04454_ sky130_fd_sc_hd__mux2_1
X_08890_ net1224 top.WB.CPU_DAT_O\[12\] net306 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__mux2_1
X_07841_ top.findLeastValue.sum\[29\] _04398_ net390 vssd1 vssd1 vccd1 vccd1 _04399_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07772_ net479 _04342_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__or2_1
X_09511_ net732 net567 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__and2_1
X_06723_ top.compVal\[37\] _02460_ _02461_ top.compVal\[36\] vssd1 vssd1 vccd1 vccd1
+ _03521_ sky130_fd_sc_hd__o22a_1
XANTENNA__05763__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__and2_1
X_06654_ top.compVal\[13\] _02495_ _03450_ _03451_ _03429_ vssd1 vssd1 vccd1 vccd1
+ _03452_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06585_ top.cb_syn.zeroes\[5\] top.cb_syn.zeroes\[4\] top.cb_syn.zeroes\[3\] top.cb_syn.zeroes\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__or4_1
X_05605_ top.cb_syn.char_path\[20\] net548 net539 top.cb_syn.char_path\[84\] vssd1
+ vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ top.hTree.nulls\[50\] net398 net229 vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout244_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08324_ net1716 net202 _04724_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__o21a_1
XANTENNA__07268__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05536_ net207 _02619_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__and2b_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ top.cb_syn.char_path_n\[77\] net384 net339 top.cb_syn.char_path_n\[75\] net186
+ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a221o_1
X_05467_ net12 net415 net364 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 _02391_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout509_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08217__C1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ net1744 net205 _04655_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__o21a_1
X_05398_ top.findLeastValue.least2\[6\] vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__inv_2
X_07206_ _02464_ _02488_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07137_ top.findLeastValue.val2\[9\] top.findLeastValue.val1\[9\] vssd1 vssd1 vccd1
+ vccd1 _03813_ sky130_fd_sc_hd__nand2_1
XANTENNA__05487__B top.WB.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ top.findLeastValue.val2\[29\] top.findLeastValue.val1\[29\] vssd1 vssd1 vccd1
+ vccd1 _03744_ sky130_fd_sc_hd__nor2_1
XANTENNA__08615__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06019_ top.sram_interface.init_counter\[10\] top.sram_interface.init_counter\[9\]
+ _02931_ net1101 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a31o_1
XANTENNA__08940__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ clknet_leaf_39_clk _01546_ _00371_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_09709_ net839 net674 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10568__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ clknet_leaf_0_clk top.dut.bit_buf_next\[9\] _00992_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ clknet_leaf_70_clk _02098_ _00923_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ clknet_leaf_78_clk _02029_ _00854_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[21\]
+ sky130_fd_sc_hd__dfstp_1
X_10415_ net742 net577 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11395_ clknet_leaf_12_clk _01960_ _00785_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.wipe_the_char_2
+ sky130_fd_sc_hd__dfrtp_1
X_10346_ net776 net611 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__and2_1
X_10277_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__and2_1
XANTENNA__05993__A0 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__S _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05860__B top.WB.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__A2_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06370_ _02504_ net534 net407 _02578_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_64_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08998__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05321_ top.compVal\[8\] vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__inv_2
X_08040_ net488 net550 net412 net524 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or4b_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08214__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09991_ net860 net695 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__and2_1
XANTENNA__07422__B1 _03660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08942_ top.WB.CPU_DAT_O\[26\] net1265 net318 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__mux2_1
XANTENNA__05984__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ net1116 top.WB.CPU_DAT_O\[29\] net303 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__mux2_1
X_07824_ net435 net1585 net249 top.findLeastValue.sum\[33\] _04385_ vssd1 vssd1 vccd1
+ vccd1 _01822_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07755_ top.hTree.tree_reg\[46\] top.findLeastValue.least2\[0\] net281 vssd1 vssd1
+ vccd1 vccd1 _04330_ sky130_fd_sc_hd__mux2_1
X_07686_ net474 _04271_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__or2_1
X_06706_ _03490_ _03487_ _03485_ _03484_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__o2bb2a_1
X_11890__921 vssd1 vssd1 vccd1 vccd1 net921 _11890__921/LO sky130_fd_sc_hd__conb_1
X_06637_ _03433_ _03434_ _03432_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o21a_1
XANTENNA__07043__A _03394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ net754 net589 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout626_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ net1008 net225 net217 _04351_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__a22o_1
XANTENNA__08989__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06568_ _02417_ _02454_ _02561_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__or4b_1
X_08307_ top.cb_syn.char_path_n\[51\] net375 net332 top.cb_syn.char_path_n\[49\] net178
+ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05519_ _02600_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__or2_1
X_09287_ top.histogram.total\[16\] net402 net323 top.histogram.total\[17\] net429
+ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__o221a_1
X_06499_ top.histogram.total\[11\] top.histogram.total\[10\] top.histogram.total\[9\]
+ _03331_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__and4_1
X_08238_ top.cb_syn.char_path_n\[85\] net198 _04681_ vssd1 vssd1 vccd1 vccd1 _01704_
+ sky130_fd_sc_hd__o21a_1
X_08169_ top.cb_syn.char_path_n\[120\] net374 net330 top.cb_syn.char_path_n\[118\]
+ net177 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__a221o_1
XANTENNA__07413__A0 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ net819 net654 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08602__A _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ clknet_leaf_38_clk _01745_ _00570_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[126\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06821__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10131_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__and2_1
XANTENNA__05975__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__B2 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ net720 net555 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__and2_1
XANTENNA__05727__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ clknet_leaf_57_clk _01529_ _00354_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_10895_ clknet_leaf_31_clk _01467_ _00285_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07247__A3 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ clknet_leaf_118_clk _02081_ _00906_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05839__C net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11447_ clknet_leaf_89_clk _02012_ _00837_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ clknet_leaf_17_clk _01943_ _00768_ vssd1 vssd1 vccd1 vccd1 top.cw2\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07404__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10329_ net768 net603 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07707__A1 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05870_ net1524 top.WB.CPU_DAT_O\[28\] net353 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__mux2_1
XANTENNA__05718__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _04138_ _04139_ net289 vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__S0 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09997__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11915__946 vssd1 vssd1 vccd1 vccd1 net946 _11915__946/LO sky130_fd_sc_hd__conb_1
X_07471_ _04072_ _04076_ _04049_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
X_09210_ net491 top.header_synthesis.write_char_path _03382_ _02566_ _05186_ vssd1
+ vssd1 vccd1 vccd1 top.header_synthesis.next_write_char_path sky130_fd_sc_hd__o221a_1
X_06422_ net1180 _03281_ net301 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06353_ net458 _03211_ _03215_ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a211o_1
X_09141_ top.WorR _02856_ _02852_ net448 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ net447 _02562_ _03013_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__or3_1
X_05304_ top.compVal\[31\] vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06284_ net445 _03053_ top.TRN_char_index\[3\] vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a21oi_1
X_08023_ net287 _04534_ _04538_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__and3_1
Xhold711 top.cb_syn.count\[4\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold700 top.compVal\[2\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout207_A _02620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 top.cb_syn.count\[1\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold744 top.hTree.nullSumIndex\[4\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 top.findLeastValue.sum\[18\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 top.dut.bits_in_buf\[1\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 top.cb_syn.zeroes\[1\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 top.header_synthesis.count\[5\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 top.hTree.nullSumIndex\[6\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__and2_1
Xhold799 top.histogram.state\[1\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
X_08925_ top.cb_syn.max_index\[3\] top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\]
+ top.cb_syn.max_index\[4\] vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout576_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05709__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _05037_ net502 _02811_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__or3b_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05781__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ net476 _04370_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ _04971_ _04972_ _04974_ _04975_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a22o_1
XANTENNA__06921__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout743_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05999_ top.WB.CPU_DAT_O\[2\] net1138 net347 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
X_07738_ net389 _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nand2_1
XANTENNA__06134__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07669_ top.findLeastValue.least1\[7\] _04259_ net389 vssd1 vssd1 vccd1 vccd1 _04260_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09408_ _02851_ _04252_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nor2_1
X_10680_ clknet_leaf_116_clk _01311_ _00070_ vssd1 vssd1 vccd1 vccd1 top.path\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_09339_ net1516 net223 net214 _04419_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06988__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ clknet_leaf_2_clk _01866_ _00691_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05660__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ clknet_leaf_66_clk _01797_ _00622_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09387__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ clknet_leaf_60_clk _01728_ _00553_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_10114_ net802 net637 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__and2_1
XANTENNA__05948__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11094_ clknet_leaf_62_clk _01659_ _00484_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[40\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08478__S net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10045_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold82 net56 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 top.hTree.tree_reg\[47\] vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 top.hTree.node_reg\[52\] vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 top.path\[8\] vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06912__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07548__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__A2 _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10947_ clknet_leaf_38_clk net1427 _00337_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10878_ clknet_leaf_23_clk top.header_synthesis.next_header\[0\] _00268_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07557__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05651__A2 _02714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05866__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09057__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05939__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 net512 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_4
X_06971_ net482 top.findLeastValue.histo_index\[5\] _03670_ vssd1 vssd1 vccd1 vccd1
+ _03672_ sky130_fd_sc_hd__and3_1
X_09690_ net874 net709 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__and2_1
X_08710_ _03375_ _04906_ _04895_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_72_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05922_ top.sram_interface.CB_write_counter\[0\] _02587_ _02903_ vssd1 vssd1 vccd1
+ vccd1 _02904_ sky130_fd_sc_hd__o21ai_1
X_08641_ top.cb_syn.end_cnt\[6\] _04809_ _04826_ _04843_ _04860_ vssd1 vssd1 vccd1
+ vccd1 _04861_ sky130_fd_sc_hd__a32o_1
XANTENNA__08908__A2_N _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05853_ _02848_ _02855_ _02870_ _02867_ net1690 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a32o_1
XANTENNA__07539__S0 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ _04199_ _04630_ _04791_ top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1 vccd1 _04792_
+ sky130_fd_sc_hd__o22ai_2
X_05784_ top.translation.index\[6\] top.translation.index\[5\] _02812_ vssd1 vssd1
+ vccd1 vccd1 _02814_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07523_ top.cb_syn.char_path_n\[118\] top.cb_syn.char_path_n\[117\] top.cb_syn.char_path_n\[120\]
+ top.cb_syn.char_path_n\[119\] net394 net295 vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__mux4_1
XANTENNA__07864__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A _03017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09520__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ top.dut.bit_buf\[12\] top.dut.bit_buf\[5\] net713 vssd1 vssd1 vccd1 vccd1
+ _04062_ sky130_fd_sc_hd__mux2_1
X_06405_ top.hist_data_o\[31\] _03265_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout324_A _04917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07385_ _03845_ _03847_ _03842_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a21o_1
X_06336_ net487 top.findLeastValue.histo_index\[0\] top.findLeastValue.histo_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09081__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ top.histogram.state\[6\] _05124_ _05130_ net1479 vssd1 vssd1 vccd1 vccd1
+ _00035_ sky130_fd_sc_hd__a22o_1
X_09055_ top.CB_write_complete top.cb_syn.end_cond top.cb_syn.curr_state\[8\] _05087_
+ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a31o_1
X_06267_ _03124_ _03138_ _03128_ _03137_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__or4b_1
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05642__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 top.hist_data_o\[25\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
X_08006_ _04527_ net1655 _04522_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__mux2_1
X_06198_ top.cw1\[5\] top.cw1\[4\] _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__and3_1
Xhold563 top.histogram.state\[6\] vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 top.hTree.tree_reg\[35\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 top.histogram.total\[13\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05495__B top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 top.hist_data_o\[22\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _01815_ vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 net47 vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07395__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ net773 net608 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__and2_1
X_08908_ top.hTree.finish_check _04254_ _05053_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_
+ sky130_fd_sc_hd__o2bb2a_1
X_09888_ net875 net710 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__and2_1
XANTENNA__08344__A1 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _05026_ _05027_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__and2b_1
X_11850_ clknet_leaf_96_clk _02383_ _01222_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10801_ clknet_leaf_18_clk _01404_ _00191_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06370__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ clknet_leaf_3_clk _00016_ _01153_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.write_HT_fin_n
+ sky130_fd_sc_hd__dfrtp_1
X_10732_ clknet_leaf_25_clk _01363_ _00122_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10663_ clknet_leaf_106_clk _01294_ _00053_ vssd1 vssd1 vccd1 vccd1 top.path\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07607__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ net737 net572 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__and2_1
XANTENNA__08804__C1 top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05633__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
X_11215_ clknet_leaf_43_clk _01780_ _00605_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__clkbuf_4
X_11146_ clknet_leaf_34_clk _01711_ _00536_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[92\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput72 net441 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
X_11077_ clknet_leaf_52_clk _01642_ _00467_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_10028_ net855 net690 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07840__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07170_ top.findLeastValue.val2\[6\] top.findLeastValue.val1\[6\] _03844_ _03843_
+ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06121_ net453 top.histogram.eof_n _02561_ net1034 vssd1 vssd1 vccd1 vccd1 _02148_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__05624__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06052_ _02950_ _02951_ top.cb_syn.count\[6\] _02527_ vssd1 vssd1 vccd1 vccd1 _02952_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08810__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
Xfanout328 net331 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
X_09811_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 _02918_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_2
Xfanout317 _05083_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_2
X_09742_ net842 net677 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__and2_1
X_06954_ top.findLeastValue.val1\[3\] net135 net112 net1698 vssd1 vssd1 vccd1 vccd1
+ _01964_ sky130_fd_sc_hd__o22a_1
X_05905_ _02884_ _02885_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__nor2_1
X_06885_ top.compVal\[11\] top.findLeastValue.val1\[11\] net155 vssd1 vssd1 vccd1
+ vccd1 _03648_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout274_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ net734 net569 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ top.cb_syn.char_path_n\[59\] top.cb_syn.char_path_n\[60\] top.cb_syn.char_path_n\[63\]
+ top.cb_syn.char_path_n\[64\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__mux4_1
X_05836_ net448 _02845_ _02852_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_85_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ net1334 top.cb_syn.char_path_n\[4\] net237 vssd1 vssd1 vccd1 vccd1 _01487_
+ sky130_fd_sc_hd__mux2_1
X_05767_ top.compVal\[41\] net163 _02806_ top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1
+ vccd1 _02326_ sky130_fd_sc_hd__a22o_1
X_07506_ _02988_ _04105_ _02986_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout539_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05560__B2 top.hTree.node_reg\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09287__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ net1176 top.cb_syn.char_path_n\[73\] net240 vssd1 vssd1 vccd1 vccd1 _01556_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05698_ _02753_ _02754_ net468 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ _02405_ top.dut.bits_in_buf\[0\] top.dut.bits_in_buf\[1\] vssd1 vssd1 vccd1
+ vccd1 _04047_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_33_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07368_ _03810_ _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06319_ top.cw2\[3\] _03077_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__xnor2_1
X_09107_ _02594_ _05122_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__or2_1
XANTENNA__05615__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07299_ _03741_ _03745_ _03959_ top.findLeastValue.val1\[30\] top.findLeastValue.val2\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__a32o_1
XANTENNA__08660__B1_N _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ top.WB.CPU_DAT_O\[12\] net1095 net315 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
Xhold371 top.cb_syn.char_path\[44\] vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 top.path\[106\] vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ clknet_leaf_54_clk _01565_ _00390_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[82\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold382 top.cb_syn.char_path\[123\] vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 top.hTree.nulls\[57\] vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout851 net854 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout840 net844 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout873 net874 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout862 net865 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ net933 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_11833_ clknet_leaf_46_clk _02366_ _01205_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11764_ clknet_leaf_47_clk _02303_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10715_ clknet_leaf_75_clk _01346_ _00105_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_11695_ clknet_leaf_99_clk _02245_ _01085_ vssd1 vssd1 vccd1 vccd1 top.compVal\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_10646_ clknet_leaf_103_clk _01277_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10577_ net785 net620 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_102_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05606__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ clknet_leaf_60_clk _01694_ _00519_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[75\]
+ sky130_fd_sc_hd__dfrtp_2
X_06670_ _03459_ _03460_ _03462_ _03464_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_108_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05621_ top.hTree.node_reg\[50\] net355 _02689_ _02690_ vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__05542__B2 top.hTree.node_reg\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05552_ top.cb_syn.char_path\[29\] net546 net309 top.cb_syn.char_path\[125\] vssd1
+ vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__a22o_1
X_08340_ top.cb_syn.char_path_n\[34\] net200 _04732_ vssd1 vssd1 vccd1 vccd1 _01653_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_50_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07819__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08271_ top.cb_syn.char_path_n\[69\] net375 net333 top.cb_syn.char_path_n\[67\] net178
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a221o_1
X_05483_ net27 net416 _02570_ top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 _02375_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07222_ _03896_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__and2_1
X_07153_ top.findLeastValue.val2\[0\] top.findLeastValue.val1\[0\] vssd1 vssd1 vccd1
+ vccd1 _03829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06104_ _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06215__A top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ top.findLeastValue.val2\[31\] top.findLeastValue.val1\[31\] _03758_ _03759_
+ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a211oi_1
X_06035_ _02924_ _02926_ _02938_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09526__A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923__886 vssd1 vssd1 vccd1 vccd1 _11923__886/HI net886 sky130_fd_sc_hd__conb_1
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 _02806_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_4
Xfanout114 _03661_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_4
Xfanout136 net138 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_2
Xfanout169 net171 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_4
X_07986_ top.findLeastValue.sum\[0\] _04514_ net391 vssd1 vssd1 vccd1 vccd1 _04515_
+ sky130_fd_sc_hd__mux2_1
X_09725_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__and2_1
X_06937_ top.findLeastValue.val1\[20\] net138 net116 top.compVal\[20\] vssd1 vssd1
+ vccd1 vccd1 _01981_ sky130_fd_sc_hd__o22a_1
X_09656_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08607_ top.cb_syn.char_path_n\[25\] top.cb_syn.char_path_n\[26\] top.cb_syn.char_path_n\[29\]
+ top.cb_syn.char_path_n\[30\] net498 net492 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06868_ top.findLeastValue.val2\[20\] net132 net117 _03639_ vssd1 vssd1 vccd1 vccd1
+ _02028_ sky130_fd_sc_hd__o22a_1
X_09587_ net799 net634 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__and2_1
X_06799_ _03560_ _03596_ _03584_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__o21a_1
X_05819_ net442 top.sram_interface.counter_HTREE\[3\] top.sram_interface.counter_HTREE\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__nor3_1
X_08538_ net1171 top.cb_syn.char_path_n\[21\] net235 vssd1 vssd1 vccd1 vccd1 _01504_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08469_ net1132 top.cb_syn.char_path_n\[90\] net234 vssd1 vssd1 vccd1 vccd1 _01573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07286__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07286__B2 top.findLeastValue.sum\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ net734 net569 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__and2_1
X_11480_ clknet_leaf_95_clk _02045_ _00870_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[37\]
+ sky130_fd_sc_hd__dfstp_1
X_10431_ net822 net657 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08786__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ net727 net562 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__and2_1
X_10293_ net861 net696 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__and2_1
Xhold190 top.cb_syn.char_path\[36\] vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout681 net689 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_2
Xfanout692 net693 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_2
Xfanout670 net712 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05772__B2 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11816_ clknet_leaf_67_clk _02349_ _01188_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07277__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11747_ clknet_leaf_11_clk _02297_ _01137_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.zero_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11678_ clknet_leaf_86_clk _02228_ _01068_ vssd1 vssd1 vccd1 vccd1 top.compVal\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ clknet_leaf_66_clk _01260_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__S _04110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08624__S1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ top.hTree.tree_reg\[29\] top.findLeastValue.sum\[29\] net282 vssd1 vssd1
+ vccd1 vccd1 _04398_ sky130_fd_sc_hd__mux2_1
X_07771_ top.hTree.tree_reg\[43\] top.findLeastValue.sum\[43\] _04251_ vssd1 vssd1
+ vccd1 vccd1 _04343_ sky130_fd_sc_hd__mux2_1
X_09510_ net735 net570 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__and2_1
XANTENNA__06960__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06722_ top.compVal\[34\] _02463_ _02464_ top.compVal\[33\] _03519_ vssd1 vssd1 vccd1
+ vccd1 _03520_ sky130_fd_sc_hd__a221o_1
XANTENNA__05763__B2 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06653_ top.compVal\[12\] top.findLeastValue.val1\[12\] vssd1 vssd1 vccd1 vccd1 _03451_
+ sky130_fd_sc_hd__nand2b_1
X_09441_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_35_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06584_ top.header_synthesis.write_num_lefts _03377_ _03381_ _03383_ vssd1 vssd1
+ vccd1 vccd1 _03384_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_82_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05604_ net1484 net169 _02676_ net211 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a22o_1
X_09372_ net398 _04312_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__nand2_1
XANTENNA__10020__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ top.cb_syn.char_path_n\[43\] net381 net338 top.cb_syn.char_path_n\[41\] net184
+ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07268__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05535_ top.WB.curr_state\[0\] _02572_ _02617_ net213 vssd1 vssd1 vccd1 vccd1 _02620_
+ sky130_fd_sc_hd__a31o_1
X_08254_ top.cb_syn.char_path_n\[77\] net204 _04689_ vssd1 vssd1 vccd1 vccd1 _01696_
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05466_ net14 net413 net362 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 _02392_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08185_ top.cb_syn.char_path_n\[112\] net385 net340 top.cb_syn.char_path_n\[110\]
+ net188 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a221o_1
X_05397_ top.findLeastValue.least2\[8\] vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout404_A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07205_ _03877_ _03878_ _03879_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__or3_1
XANTENNA__06228__C1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ top.findLeastValue.val2\[9\] top.findLeastValue.val1\[9\] vssd1 vssd1 vccd1
+ vccd1 _03812_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07067_ top.findLeastValue.val2\[29\] top.findLeastValue.val1\[29\] vssd1 vssd1 vccd1
+ vccd1 _03743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06018_ top.sram_interface.init_counter\[8\] top.sram_interface.init_counter\[7\]
+ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__and3_1
XANTENNA__05784__A top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__S1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09708_ net784 net619 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__and2_1
XANTENNA__06951__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ net436 net1318 net249 top.findLeastValue.sum\[4\] _04501_ vssd1 vssd1 vccd1
+ vccd1 _01793_ sky130_fd_sc_hd__a221o_1
XANTENNA__08153__C1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ clknet_leaf_39_clk _01545_ _00370_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06819__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09639_ net760 net595 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ clknet_leaf_1_clk top.dut.bit_buf_next\[8\] _00991_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ clknet_leaf_81_clk _02097_ _00922_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11463_ clknet_leaf_78_clk _02028_ _00853_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[20\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05690__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ net737 net572 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_36_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11394_ clknet_leaf_13_clk _01959_ _00784_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.wipe_the_char_1
+ sky130_fd_sc_hd__dfrtp_1
X_10345_ net776 net611 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10276_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_45_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06942__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05320_ top.compVal\[9\] vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06464__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07422__B2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09990_ net831 net666 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__and2_1
X_08941_ top.WB.CPU_DAT_O\[27\] net1267 net319 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__mux2_1
X_08872_ net1062 top.WB.CPU_DAT_O\[30\] net303 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__mux2_1
XANTENNA__09175__A1 top.WB.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07823_ net418 _04383_ _04384_ net260 vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__o211a_1
XANTENNA__05736__A1 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06933__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ net257 _04328_ _04329_ net1011 net433 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a32o_1
X_07685_ net474 _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06705_ _03477_ _03502_ _03488_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout354_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
X_06636_ _02444_ top.findLeastValue.val1\[2\] top.findLeastValue.val1\[1\] _02445_
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__a22o_1
X_09424_ net747 net582 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__and2_1
XANTENNA__07043__B _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ net1014 net227 net217 _04355_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__a22o_1
X_06567_ top.dut.out\[2\] top.dut.out\[1\] _03367_ top.dut.out\[3\] vssd1 vssd1 vccd1
+ vccd1 _03368_ sky130_fd_sc_hd__and4b_1
X_08306_ net1756 net197 _04715_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_72_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05518_ _02563_ _02602_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__nor2_2
X_06498_ top.histogram.total\[8\] _03325_ _03328_ _03330_ vssd1 vssd1 vccd1 vccd1
+ _03331_ sky130_fd_sc_hd__and4_1
X_09286_ net425 _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__or2_1
X_08237_ top.cb_syn.char_path_n\[86\] net377 net334 top.cb_syn.char_path_n\[84\] net180
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a221o_1
X_05449_ top.header_synthesis.write_num_lefts vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__inv_2
X_11888__884 vssd1 vssd1 vccd1 vccd1 _11888__884/HI net884 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05672__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929__892 vssd1 vssd1 vccd1 vccd1 _11929__892/HI net892 sky130_fd_sc_hd__conb_1
X_08168_ top.cb_syn.char_path_n\[120\] net194 _04646_ vssd1 vssd1 vccd1 vccd1 _01739_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09402__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ _04590_ _04597_ _04599_ _04589_ net1682 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a32o_1
X_07119_ _03793_ _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__and2_1
X_10130_ net781 net616 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__and2_1
X_10061_ net720 net555 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__and2_1
XANTENNA__06924__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ clknet_leaf_61_clk _01528_ _00353_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10579__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_82_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
X_10894_ clknet_leaf_34_clk _01466_ _00284_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_26_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07652__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11515_ clknet_leaf_118_clk _02080_ _00905_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05663__B1 _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ clknet_leaf_89_clk _02011_ _00836_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11377_ clknet_leaf_40_clk _01942_ _00767_ vssd1 vssd1 vccd1 vccd1 top.cw2\[1\] sky130_fd_sc_hd__dfrtp_1
X_10328_ net767 net602 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__and2_1
XANTENNA__08365__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__and2_1
XANTENNA__06459__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07566__S1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_45_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07470_ top.dut.bit_buf\[5\] net43 net713 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__mux2_1
X_06421_ _03262_ _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06352_ top.cb_syn.char_index\[0\] _02607_ _03219_ vssd1 vssd1 vccd1 vccd1 _03220_
+ sky130_fd_sc_hd__a21o_1
X_09140_ net543 net466 _02901_ _05147_ _02802_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__a311o_1
X_06283_ net446 _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__nand2_1
X_09071_ _02715_ _05099_ _02915_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__or3b_1
X_05303_ top.hist_data_o\[0\] vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__inv_2
XANTENNA__05654__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08022_ net456 _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold701 top.header_synthesis.count\[6\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 top.hist_data_o\[17\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold723 top.header_synthesis.char_added vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold734 top.hist_addr\[6\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold745 top.findLeastValue.sum\[37\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 top.hist_data_o\[19\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ net782 net617 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__and2_1
Xhold756 top.findLeastValue.sum\[16\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 top.compVal\[12\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ _05068_ top.cb_syn.max_index\[5\] _05059_ vssd1 vssd1 vccd1 vccd1 _01405_
+ sky130_fd_sc_hd__mux2_1
Xhold789 top.hist_addr\[0\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05957__B2 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _02546_ _02812_ _05039_ _05041_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout471_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ top.path\[9\] net324 _04973_ net426 net429 vssd1 vssd1 vccd1 vccd1 _04975_
+ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05781__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ top.findLeastValue.sum\[36\] _04370_ net391 vssd1 vssd1 vccd1 vccd1 _04371_
+ sky130_fd_sc_hd__mux2_1
X_07737_ top.hTree.tree_reg\[49\] top.findLeastValue.least2\[3\] net280 vssd1 vssd1
+ vccd1 vccd1 _04315_ sky130_fd_sc_hd__mux2_1
X_05998_ top.WB.CPU_DAT_O\[3\] net1412 net347 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_64_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout736_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07668_ top.findLeastValue.least1\[7\] top.hTree.tree_reg\[62\] _04248_ vssd1 vssd1
+ vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07599_ top.cb_syn.cb_length\[6\] top.cb_syn.cb_length\[5\] _04198_ vssd1 vssd1 vccd1
+ vccd1 _04199_ sky130_fd_sc_hd__or3_1
X_09407_ net988 _05284_ net229 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_80_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06619_ top.findLeastValue.val1\[19\] top.compVal\[19\] vssd1 vssd1 vccd1 vccd1 _03417_
+ sky130_fd_sc_hd__and2b_1
X_09338_ net1006 net221 net214 _04423_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__a22o_1
XANTENNA__09084__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05302__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ _04046_ _04067_ _04090_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[2\]
+ sky130_fd_sc_hd__o21a_1
X_11300_ clknet_leaf_2_clk _01865_ _00690_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11231_ clknet_leaf_83_clk _01796_ _00621_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11162_ clknet_leaf_60_clk _01727_ _00552_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[108\]
+ sky130_fd_sc_hd__dfrtp_2
X_10113_ net806 net641 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__and2_1
XANTENNA__05948__B2 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897__928 vssd1 vssd1 vccd1 vccd1 net928 _11897__928/LO sky130_fd_sc_hd__conb_1
X_11093_ clknet_leaf_65_clk _01658_ _00483_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[39\]
+ sky130_fd_sc_hd__dfrtp_2
X_10044_ net783 net618 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__and2_1
Xhold50 top.hTree.node_reg\[33\] vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 net55 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 top.dut.out\[6\] vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 top.histogram.out_of_init vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 top.histogram.sram_out\[23\] vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_55_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
X_10946_ clknet_leaf_35_clk _01511_ _00336_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07548__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07322__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ clknet_leaf_26_clk top.header_synthesis.next_char_added _00267_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.char_added sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05636__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07625__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07625__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ clknet_leaf_96_clk _01994_ _00819_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[33\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_113_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07389__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05939__B2 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06970_ net483 _03670_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05921_ _02553_ net460 _02588_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__a31o_1
XANTENNA__08353__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ top.cb_syn.end_cnt\[5\] _04859_ top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1
+ vccd1 _04860_ sky130_fd_sc_hd__a21oi_1
X_05852_ net1640 _02872_ _02869_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__o21a_1
X_08571_ top.cb_syn.end_cnt\[5\] top.cb_syn.end_cnt\[4\] _04790_ vssd1 vssd1 vccd1
+ vccd1 _04791_ sky130_fd_sc_hd__or3_2
Xclkbuf_leaf_46_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
X_05783_ _02812_ _02546_ _02545_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__and3b_1
XANTENNA__07539__S1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07522_ _04120_ _04121_ net289 vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07864__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ net344 _04044_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__or2_1
X_06404_ top.hist_data_o\[20\] top.hist_data_o\[19\] _03268_ vssd1 vssd1 vccd1 vccd1
+ _03269_ sky130_fd_sc_hd__and3_1
X_09123_ _02417_ net1514 _05134_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07384_ net1789 net277 net272 _04021_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06335_ net487 _02787_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ top.cb_syn.char_path_n\[1\] _04202_ _04585_ _05085_ vssd1 vssd1 vccd1 vccd1
+ _05087_ sky130_fd_sc_hd__a22o_1
X_06266_ top.cb_syn.curr_index\[6\] _02584_ _03134_ net446 _03130_ vssd1 vssd1 vccd1
+ vccd1 _03138_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08005_ top.findLeastValue.least2\[3\] top.findLeastValue.least1\[3\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_1
Xhold520 top.path\[97\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 top.cb_syn.end_cond vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
X_06197_ top.cw1\[3\] _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__or2_1
Xhold553 _03355_ vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold542 top.hTree.tree_reg\[29\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 top.cb_syn.state8 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 top.hist_data_o\[31\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 top.hTree.tree_reg\[31\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 net46 vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09956_ net772 net607 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__and2_1
X_09887_ net873 net708 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__and2_1
X_08907_ net288 _04255_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ top.TRN_char_index\[2\] top.TRN_char_index\[1\] top.TRN_char_index\[4\] top.TRN_char_index\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_37_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_08769_ _04934_ _04935_ _04936_ net429 net502 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_28_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ clknet_leaf_17_clk _01403_ _00190_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_56_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07304__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06827__S net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ clknet_leaf_3_clk _00015_ _01152_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10731_ clknet_leaf_17_clk _01362_ _00121_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_10662_ clknet_leaf_68_clk _01293_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10593_ net745 net580 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__and2_1
XANTENNA__05618__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09158__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06830__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11214_ clknet_leaf_15_clk _01779_ _00604_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
X_11145_ clknet_leaf_35_clk _01710_ _00535_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[91\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_8_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
X_11076_ clknet_leaf_52_clk _01641_ _00466_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
X_10027_ net855 net690 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09902__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
X_10929_ clknet_leaf_60_clk _01494_ _00319_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09048__A0 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06120_ _02996_ _02997_ _02453_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XANTENNA__07568__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06051_ top.cb_syn.count\[5\] _02528_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout329 net331 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
X_09810_ net764 net599 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__and2_1
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
Xfanout318 net319 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
X_09741_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__and2_1
X_06953_ top.findLeastValue.val1\[4\] net135 net112 top.compVal\[4\] vssd1 vssd1 vccd1
+ vccd1 _01965_ sky130_fd_sc_hd__o22a_1
X_05904_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06884_ top.findLeastValue.val2\[12\] net130 net119 _03647_ vssd1 vssd1 vccd1 vccd1
+ _02020_ sky130_fd_sc_hd__o22a_1
X_09672_ net750 net585 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__and2_1
X_08623_ _02540_ _04838_ _04842_ _04834_ top.cb_syn.end_cnt\[5\] vssd1 vssd1 vccd1
+ vccd1 _04843_ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_19_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_05835_ top.WorR _02856_ net544 _02847_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__and4bb_1
XANTENNA__06888__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ net1420 top.cb_syn.char_path_n\[5\] net237 vssd1 vssd1 vccd1 vccd1 _01488_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout267_A _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05766_ top.compVal\[42\] net163 net147 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XANTENNA__09287__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _02979_ _02989_ _04103_ _02978_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__o31ai_2
XANTENNA__05560__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08485_ net1362 top.cb_syn.char_path_n\[74\] net241 vssd1 vssd1 vccd1 vccd1 _01557_
+ sky130_fd_sc_hd__mux2_1
X_05697_ top.cb_syn.char_path\[37\] net529 net310 top.cb_syn.char_path\[101\] vssd1
+ vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a22o_1
XANTENNA__09039__A0 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ top.dut.out_valid_next _04044_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout601_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ _03806_ _04008_ _03804_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06318_ top.findLeastValue.histo_index\[2\] net406 _03186_ net535 vssd1 vssd1 vccd1
+ vccd1 _03187_ sky130_fd_sc_hd__o211a_1
X_09106_ _02594_ _05122_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nor2_1
XANTENNA__08798__C1 _02547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ top.WB.CPU_DAT_O\[13\] net1181 net315 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
X_07298_ _03745_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__nand2_1
X_06249_ _02602_ _03073_ _03117_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold361 top.histogram.sram_out\[13\] vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 top.hTree.nulls\[63\] vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 top.cb_syn.char_path\[8\] vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 top.cb_syn.char_path\[4\] vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 top.path\[75\] vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_2
Xfanout841 net844 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_1
Xfanout830 net835 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_09939_ net791 net626 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__and2_1
Xfanout863 net865 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_1
XANTENNA__06130__B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07941__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11901_ net932 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_11832_ clknet_leaf_82_clk _02365_ _01204_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05551__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ clknet_leaf_72_clk _02302_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10714_ clknet_leaf_75_clk _01345_ _00104_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ clknet_leaf_103_clk _02244_ _01084_ vssd1 vssd1 vccd1 vccd1 top.compVal\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_10645_ clknet_leaf_104_clk _01276_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10576_ net784 net619 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08801__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ clknet_leaf_59_clk _01693_ _00518_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[74\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07764__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ clknet_leaf_71_clk _01624_ _00449_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07851__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05620_ top.histogram.sram_out\[18\] net358 net410 top.hTree.node_reg\[18\] vssd1
+ vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a22o_1
XANTENNA__06467__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05542__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05551_ top.cb_syn.char_path\[93\] net537 net528 top.cb_syn.char_path\[61\] vssd1
+ vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07819__B2 top.findLeastValue.sum\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08270_ net1773 net196 _04697_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05482_ net28 net414 net362 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 _02376_
+ sky130_fd_sc_hd__o22a_1
X_07221_ top.findLeastValue.val2\[40\] top.findLeastValue.val1\[40\] vssd1 vssd1 vccd1
+ vccd1 _03897_ sky130_fd_sc_hd__nand2_1
X_07152_ top.findLeastValue.val2\[1\] top.findLeastValue.val1\[1\] vssd1 vssd1 vccd1
+ vccd1 _03828_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_30_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06103_ _02448_ _03002_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08795__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ top.findLeastValue.val2\[31\] top.findLeastValue.val1\[31\] top.findLeastValue.val1\[30\]
+ top.findLeastValue.val2\[30\] vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06034_ net1614 _02925_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__nor2_1
XANTENNA__09526__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
Xfanout115 net116 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
Xfanout137 net138 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_4
Xfanout159 _02908_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_07985_ top.hTree.tree_reg\[0\] top.findLeastValue.sum\[0\] net284 vssd1 vssd1 vccd1
+ vccd1 _04514_ sky130_fd_sc_hd__mux2_1
X_09724_ net866 net701 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__and2_1
X_06936_ top.findLeastValue.val1\[21\] net138 net116 net1701 vssd1 vssd1 vccd1 vccd1
+ _01982_ sky130_fd_sc_hd__o22a_1
X_09655_ net774 net609 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__and2_1
XANTENNA__09542__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06867_ top.compVal\[20\] top.findLeastValue.val1\[20\] net156 vssd1 vssd1 vccd1
+ vccd1 _03639_ sky130_fd_sc_hd__mux2_1
X_08606_ _04817_ _04825_ top.cb_syn.end_cnt\[5\] vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05818_ net442 net431 _02838_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout649_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09586_ net743 net578 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__and2_1
X_06798_ top.compVal\[19\] _02469_ _02470_ top.compVal\[18\] _03594_ vssd1 vssd1 vccd1
+ vccd1 _03596_ sky130_fd_sc_hd__o221a_1
X_08537_ net1304 top.cb_syn.char_path_n\[22\] net235 vssd1 vssd1 vccd1 vccd1 _01505_
+ sky130_fd_sc_hd__mux2_1
X_05749_ top.findLeastValue.startup _02792_ net457 vssd1 vssd1 vccd1 vccd1 _02793_
+ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout816_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ net1439 top.cb_syn.char_path_n\[91\] net236 vssd1 vssd1 vccd1 vccd1 _01574_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ _02522_ net133 _03664_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_98_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08399_ top.cb_syn.char_path_n\[5\] net375 net332 top.cb_syn.char_path_n\[3\] net178
+ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ net822 net657 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__and2_1
XANTENNA__06125__B top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ net716 net551 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__and2_1
X_10292_ net857 net692 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__and2_1
XANTENNA__07936__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07994__B1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 top.hTree.tree_reg\[60\] vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold191 top.path\[38\] vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout660 net661 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_2
Xfanout682 net689 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_2
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout671 net680 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05772__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ clknet_leaf_67_clk _02348_ _01187_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ clknet_leaf_11_clk _02296_ _01136_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.zero_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06485__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11677_ clknet_leaf_91_clk _02227_ _01067_ vssd1 vssd1 vccd1 vccd1 top.compVal\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_10628_ clknet_leaf_67_clk _01259_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10559_ net860 net695 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07846__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05460__B2 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07410__A2_N net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ top.hTree.tree_reg\[43\] top.findLeastValue.sum\[43\] net285 vssd1 vssd1
+ vccd1 vccd1 _04342_ sky130_fd_sc_hd__mux2_1
X_06721_ top.findLeastValue.val2\[32\] _03518_ top.compVal\[32\] vssd1 vssd1 vccd1
+ vccd1 _03519_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_69_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09440_ net724 net559 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__and2_1
X_06652_ _03446_ _03447_ _03449_ _03445_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_35_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06583_ top.header_synthesis.write_num_lefts _03382_ vssd1 vssd1 vccd1 vccd1 _03383_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05603_ top.hTree.node_reg\[53\] net354 _02674_ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_
+ sky130_fd_sc_hd__a211o_1
X_09371_ net1275 net222 _05260_ _05261_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
XANTENNA__10020__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ top.cb_syn.char_path_n\[43\] net202 _04723_ vssd1 vssd1 vccd1 vccd1 _01662_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05534_ _02567_ _02572_ _02618_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__or3b_2
X_08253_ top.cb_syn.char_path_n\[78\] net384 net339 top.cb_syn.char_path_n\[76\] net187
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout132_A _03611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05465_ net15 net415 net364 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 _02393_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07204_ _03878_ _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nor2_1
XANTENNA__08217__A1 top.cb_syn.char_path_n\[96\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08184_ net1759 net199 _04654_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__o21a_1
X_05396_ top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07135_ _03806_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and2_1
XANTENNA__07756__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__A0 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ _03740_ _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06017_ top.sram_interface.init_counter\[6\] _02929_ vssd1 vssd1 vccd1 vccd1 _02930_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_30_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05784__B top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ net419 _04499_ _04500_ net261 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o211a_1
X_09707_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__and2_1
X_06919_ top.findLeastValue.val1\[38\] net137 net114 top.compVal\[38\] vssd1 vssd1
+ vccd1 vccd1 _01999_ sky130_fd_sc_hd__o22a_1
X_07899_ net438 net1570 net252 top.findLeastValue.sum\[18\] _04445_ vssd1 vssd1 vccd1
+ vccd1 _01807_ sky130_fd_sc_hd__a221o_1
X_09638_ net761 net596 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__and2_1
X_09569_ net787 net622 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__and2_1
X_11600_ clknet_leaf_0_clk top.dut.bit_buf_next\[7\] _00990_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[7\] sky130_fd_sc_hd__dfrtp_1
X_11531_ clknet_leaf_81_clk _02096_ _00921_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06835__S net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11462_ clknet_leaf_78_clk _02027_ _00852_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[19\]
+ sky130_fd_sc_hd__dfstp_2
X_11393_ clknet_leaf_12_clk _01958_ _00783_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_FLV
+ sky130_fd_sc_hd__dfrtp_1
X_10413_ net742 net577 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__and2_1
X_10344_ net775 net610 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ net721 net556 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__and2_1
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09182__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06155__C1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ clknet_leaf_42_clk _02279_ _01119_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05681__B2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ top.WB.CPU_DAT_O\[28\] net1468 net318 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08871_ net1057 top.WB.CPU_DAT_O\[31\] net303 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__mux2_1
X_07822_ net476 _04382_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__or2_1
X_07753_ net472 _04325_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or2_1
X_07684_ top.findLeastValue.least1\[4\] net264 _04270_ vssd1 vssd1 vccd1 vccd1 _04272_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_48_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06704_ top.compVal\[38\] _02485_ _03481_ _03501_ _03480_ vssd1 vssd1 vccd1 vccd1
+ _03502_ sky130_fd_sc_hd__o311a_1
X_06635_ _02445_ top.findLeastValue.val1\[1\] top.findLeastValue.val1\[0\] _02446_
+ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__o211a_1
X_09423_ net754 net589 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__and2_1
X_09354_ net1007 net227 net216 _04359_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout347_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ top.cb_syn.char_path_n\[52\] net376 net332 top.cb_syn.char_path_n\[50\] net179
+ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06566_ top.dut.out\[0\] _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__nor2_1
X_05517_ top.findLeastValue.wipe_the_char_1 _02576_ vssd1 vssd1 vccd1 vccd1 _02602_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06497_ top.histogram.total\[7\] top.histogram.total\[6\] vssd1 vssd1 vccd1 vccd1
+ _03330_ sky130_fd_sc_hd__and2_1
X_09285_ top.histogram.total\[18\] top.histogram.total\[19\] net508 vssd1 vssd1 vccd1
+ vccd1 _05229_ sky130_fd_sc_hd__mux2_1
X_08236_ top.cb_syn.char_path_n\[86\] net198 _04680_ vssd1 vssd1 vccd1 vccd1 _01705_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05448_ top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__inv_2
X_08167_ top.cb_syn.char_path_n\[121\] net373 net331 top.cb_syn.char_path_n\[119\]
+ net176 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07949__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05379_ top.findLeastValue.val1\[10\] vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__inv_2
X_07118_ top.findLeastValue.val2\[15\] top.findLeastValue.val1\[15\] vssd1 vssd1 vccd1
+ vccd1 _03794_ sky130_fd_sc_hd__or2_1
XANTENNA__08610__A1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ top.cb_syn.num_lefts\[6\] _04595_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__or2_1
X_07049_ _03721_ _03722_ _03723_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10060_ net720 net555 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__and2_1
XANTENNA__05727__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05734__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ clknet_leaf_61_clk _01527_ _00352_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ clknet_leaf_31_clk _01465_ _00283_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_66_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ clknet_leaf_118_clk _02079_ _00904_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05663__B2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ clknet_leaf_90_clk _02010_ _00835_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_34_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06860__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ clknet_leaf_17_clk _01941_ _00766_ vssd1 vssd1 vccd1 vccd1 top.cw2\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07404__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10327_ net730 net565 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__and2_1
X_10258_ net717 net552 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__and2_1
XANTENNA__08365__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10189_ net799 net634 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__and2_1
XANTENNA__05718__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06420_ top.hist_data_o\[26\] _03261_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06351_ top.cb_syn.curr_index\[2\] _02584_ _03216_ net446 _03218_ vssd1 vssd1 vccd1
+ vccd1 _03219_ sky130_fd_sc_hd__a221o_1
XANTENNA__09093__B2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06282_ top.cb_syn.max_index\[5\] _03102_ _03104_ top.hTree.nullSumIndex\[4\] vssd1
+ vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a22o_1
X_09070_ net462 net526 _02910_ _05097_ net546 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a32o_1
X_05302_ net448 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ top.findLeastValue.alternator_timer\[2\] top.findLeastValue.alternator_timer\[1\]
+ top.findLeastValue.alternator_timer\[0\] _02785_ _04536_ vssd1 vssd1 vccd1 vccd1
+ _04537_ sky130_fd_sc_hd__a32o_1
Xhold702 top.histogram.sram_out\[27\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold746 top.cb_syn.char_path_n\[52\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 top.cb_syn.setup vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold735 top.hist_data_o\[18\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 top.cw1\[5\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 top.cb_syn.char_path_n\[80\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 top.cb_syn.zero_count\[6\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 top.compVal\[43\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ net754 net589 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08923_ _04222_ _05067_ _04255_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05709__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ top.translation.index\[5\] _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__or2_1
X_08785_ top.path\[8\] net404 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__or2_1
X_05997_ top.WB.CPU_DAT_O\[4\] net1166 net348 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
X_07805_ top.hTree.tree_reg\[36\] top.findLeastValue.sum\[36\] net283 vssd1 vssd1
+ vccd1 vccd1 _04370_ sky130_fd_sc_hd__mux2_1
XANTENNA__08659__A1 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ net257 _04313_ _04314_ net994 net432 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a32o_1
XANTENNA__05590__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06134__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _04253_ net256 _04258_ net1371 net431 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout631_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ top.cb_syn.cb_length\[4\] top.cb_syn.cb_length\[3\] top.cb_syn.cb_length\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09406_ top.hTree.nulls\[62\] _04260_ net401 vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__mux2_1
X_06618_ top.compVal\[18\] top.findLeastValue.val1\[18\] vssd1 vssd1 vccd1 vccd1 _03416_
+ sky130_fd_sc_hd__and2b_1
X_09337_ net987 net222 net219 _04427_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__a22o_1
X_06549_ _03331_ _03358_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_23_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05893__A1 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09084__B2 top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _04046_ top.dut.bits_in_buf_next\[1\] _04094_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[1\]
+ sky130_fd_sc_hd__o21a_1
X_08219_ top.cb_syn.char_path_n\[95\] net369 net326 top.cb_syn.char_path_n\[93\] net173
+ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08831__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06842__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ net1778 top.controller.fin_reg\[2\] top.controller.fin_reg\[4\] top.controller.fin_reg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or4b_1
X_11230_ clknet_leaf_82_clk _01795_ _00620_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ clknet_leaf_61_clk _01726_ _00551_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[107\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05948__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ net809 net644 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__and2_1
XANTENNA__09139__A2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11092_ clknet_leaf_64_clk _01657_ _00482_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[38\]
+ sky130_fd_sc_hd__dfrtp_2
X_10043_ net838 net673 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__and2_1
XANTENNA__06358__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 _02310_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__A1 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold62 top.histogram.sram_out\[14\] vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 top.hTree.node_reg\[55\] vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 top.hTree.node_reg\[0\] vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 top.hTree.node_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 top.path\[22\] vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05581__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ clknet_leaf_37_clk _01510_ _00335_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07322__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ clknet_leaf_23_clk _01461_ _00266_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05884__A1 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09075__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09075__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__C1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945__908 vssd1 vssd1 vccd1 vccd1 _11945__908/HI net908 sky130_fd_sc_hd__conb_1
XANTENNA_output93_A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ clknet_leaf_98_clk _01993_ _00818_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[32\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_113_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07389__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__B2 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ clknet_leaf_94_clk _01924_ _00749_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[37\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05939__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ net542 net460 _02900_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__and3_1
XANTENNA__08889__A1 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05851_ _02855_ _02867_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nor2_1
X_08570_ top.cb_syn.end_cnt\[3\] net493 net496 net498 vssd1 vssd1 vccd1 vccd1 _04790_
+ sky130_fd_sc_hd__or4_1
X_07521_ top.cb_syn.char_path_n\[122\] top.cb_syn.char_path_n\[121\] top.cb_syn.char_path_n\[124\]
+ top.cb_syn.char_path_n\[123\] net394 net292 vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__mux4_1
X_05782_ top.translation.index\[4\] net502 net504 net402 vssd1 vssd1 vccd1 vccd1 _02812_
+ sky130_fd_sc_hd__or4_2
XFILLER_0_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07452_ net343 _04044_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__nor2_2
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06403_ top.hist_data_o\[18\] top.hist_data_o\[17\] _03267_ vssd1 vssd1 vccd1 vccd1
+ _03268_ sky130_fd_sc_hd__and3_1
XANTENNA__05875__A1 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09066__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07383_ _04019_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__xnor2_1
X_06334_ net1077 net165 _03202_ net208 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a22o_1
X_09122_ _02610_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09053_ net412 _05084_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout212_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06265_ _02585_ _03056_ _03131_ _03133_ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__o311a_1
XANTENNA__06824__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold510 top.histogram.sram_out\[29\] vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
X_06196_ top.cw1\[2\] top.cw1\[1\] top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__and3_1
X_08004_ _04526_ net1695 _04522_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__mux2_1
Xhold532 _01463_ vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 top.histogram.sram_out\[12\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 top.histogram.total\[28\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _01818_ vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 top.hTree.node_reg\[24\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 top.histogram.sram_out\[7\] vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 top.hTree.tree_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ net771 net606 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__and2_1
Xhold598 top.hist_data_o\[7\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ net872 net707 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _02418_ top.hTree.closing net470 _05051_ _05052_ vssd1 vssd1 vccd1 vccd1
+ _05053_ sky130_fd_sc_hd__a311o_1
XANTENNA__07001__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ top.TRN_char_index\[6\] top.TRN_char_index\[5\] top.TRN_char_index\[0\] top.TRN_sram_complete
+ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout846_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05563__B1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _02547_ _04929_ _04932_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_28_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ top.header_synthesis.count\[3\] top.header_synthesis.count\[2\] _04898_ vssd1
+ vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__and3_1
X_07719_ top.hTree.tree_reg\[52\] top.findLeastValue.least2\[6\] net280 vssd1 vssd1
+ vccd1 vccd1 _04300_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ clknet_leaf_17_clk _01361_ _00120_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ clknet_leaf_66_clk _01292_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06128__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08804__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10592_ net799 net634 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__and2_1
XANTENNA__06843__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06291__B2 _02607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08017__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08568__A0 _02538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ clknet_leaf_105_clk _01778_ _00603_ vssd1 vssd1 vccd1 vccd1 top.hTree.wait_cnt
+ sky130_fd_sc_hd__dfrtp_1
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
X_11905__936 vssd1 vssd1 vccd1 vccd1 net936 _11905__936/LO sky130_fd_sc_hd__conb_1
X_11144_ clknet_leaf_35_clk _01709_ _00534_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[90\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
X_11075_ clknet_leaf_52_clk _01640_ _00465_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07791__A1 top.findLeastValue.sum\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ net859 net694 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__and2_1
XANTENNA__09902__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05554__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10928_ clknet_leaf_61_clk _01493_ _00318_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ clknet_leaf_28_clk top.header_synthesis.next_zero_count\[0\] _00249_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06050_ _02448_ top.cb_syn.zeroes\[5\] top.cb_syn.zeroes\[4\] _02449_ _02949_ vssd1
+ vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09220__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__A3 top.cb_syn.char_path_n\[88\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 _02715_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
Xfanout319 net322 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_2
X_09740_ net779 net614 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__and2_1
XANTENNA__10304__A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06952_ top.findLeastValue.val1\[5\] net135 net112 net1650 vssd1 vssd1 vccd1 vccd1
+ _01966_ sky130_fd_sc_hd__o22a_1
.ends

