magic
tech sky130A
magscale 1 2
timestamp 1756832388
<< viali >>
rect 1685 37417 1719 37451
rect 3341 37417 3375 37451
rect 27813 37417 27847 37451
rect 29101 37417 29135 37451
rect 29745 37417 29779 37451
rect 34253 37417 34287 37451
rect 34897 37417 34931 37451
rect 35541 37417 35575 37451
rect 36185 37417 36219 37451
rect 36829 37417 36863 37451
rect 37933 37417 37967 37451
rect 38209 37417 38243 37451
rect 1409 37281 1443 37315
rect 5273 37213 5307 37247
rect 8217 37213 8251 37247
rect 24225 37213 24259 37247
rect 25513 37213 25547 37247
rect 25881 37213 25915 37247
rect 26801 37213 26835 37247
rect 27169 37213 27203 37247
rect 28457 37213 28491 37247
rect 30389 37213 30423 37247
rect 31033 37213 31067 37247
rect 31677 37213 31711 37247
rect 32321 37213 32355 37247
rect 32965 37213 32999 37247
rect 33609 37213 33643 37247
rect 20821 37145 20855 37179
rect 21005 37145 21039 37179
rect 7665 37077 7699 37111
rect 20637 37077 20671 37111
rect 24041 37077 24075 37111
rect 25697 37077 25731 37111
rect 26065 37077 26099 37111
rect 26617 37077 26651 37111
rect 38485 37077 38519 37111
rect 19809 36873 19843 36907
rect 21649 36873 21683 36907
rect 24225 36873 24259 36907
rect 26985 36873 27019 36907
rect 29377 36873 29411 36907
rect 19441 36805 19475 36839
rect 19657 36805 19691 36839
rect 20177 36805 20211 36839
rect 8677 36737 8711 36771
rect 8769 36737 8803 36771
rect 8953 36737 8987 36771
rect 24409 36737 24443 36771
rect 27169 36737 27203 36771
rect 38209 36737 38243 36771
rect 38485 36737 38519 36771
rect 4445 36669 4479 36703
rect 4721 36669 4755 36703
rect 6837 36669 6871 36703
rect 7113 36669 7147 36703
rect 19901 36669 19935 36703
rect 22385 36669 22419 36703
rect 22661 36669 22695 36703
rect 24869 36669 24903 36703
rect 25145 36669 25179 36703
rect 27629 36669 27663 36703
rect 27905 36669 27939 36703
rect 30941 36669 30975 36703
rect 31217 36669 31251 36703
rect 6193 36533 6227 36567
rect 8585 36533 8619 36567
rect 8953 36533 8987 36567
rect 19625 36533 19659 36567
rect 24133 36533 24167 36567
rect 26617 36533 26651 36567
rect 29469 36533 29503 36567
rect 4445 36329 4479 36363
rect 5181 36329 5215 36363
rect 7205 36329 7239 36363
rect 7481 36329 7515 36363
rect 8953 36329 8987 36363
rect 21189 36329 21223 36363
rect 21741 36329 21775 36363
rect 23489 36329 23523 36363
rect 24409 36329 24443 36363
rect 24777 36329 24811 36363
rect 27905 36329 27939 36363
rect 28365 36329 28399 36363
rect 28825 36329 28859 36363
rect 29193 36329 29227 36363
rect 29377 36329 29411 36363
rect 1409 36261 1443 36295
rect 4997 36261 5031 36295
rect 22201 36261 22235 36295
rect 5457 36193 5491 36227
rect 6929 36193 6963 36227
rect 8677 36193 8711 36227
rect 24041 36193 24075 36227
rect 25329 36193 25363 36227
rect 25973 36193 26007 36227
rect 30481 36193 30515 36227
rect 4445 36125 4479 36159
rect 4629 36125 4663 36159
rect 4721 36125 4755 36159
rect 5181 36125 5215 36159
rect 5365 36125 5399 36159
rect 5641 36125 5675 36159
rect 5825 36125 5859 36159
rect 6561 36125 6595 36159
rect 6837 36125 6871 36159
rect 7757 36125 7791 36159
rect 7941 36125 7975 36159
rect 8033 36125 8067 36159
rect 9505 36125 9539 36159
rect 19257 36125 19291 36159
rect 21097 36125 21131 36159
rect 21281 36125 21315 36159
rect 21373 36125 21407 36159
rect 21557 36125 21591 36159
rect 21649 36125 21683 36159
rect 22017 36125 22051 36159
rect 22293 36125 22327 36159
rect 22477 36125 22511 36159
rect 22845 36125 22879 36159
rect 23857 36125 23891 36159
rect 24409 36125 24443 36159
rect 24593 36125 24627 36159
rect 25145 36125 25179 36159
rect 26160 36125 26194 36159
rect 28089 36125 28123 36159
rect 28365 36125 28399 36159
rect 28549 36125 28583 36159
rect 28733 36125 28767 36159
rect 28917 36125 28951 36159
rect 30113 36125 30147 36159
rect 4997 36057 5031 36091
rect 7297 36057 7331 36091
rect 7497 36057 7531 36091
rect 19533 36057 19567 36091
rect 23949 36057 23983 36091
rect 26341 36057 26375 36091
rect 27629 36057 27663 36091
rect 27813 36057 27847 36091
rect 28273 36057 28307 36091
rect 29009 36057 29043 36091
rect 29561 36057 29595 36091
rect 30757 36057 30791 36091
rect 38485 36057 38519 36091
rect 4813 35989 4847 36023
rect 5917 35989 5951 36023
rect 7665 35989 7699 36023
rect 7849 35989 7883 36023
rect 21005 35989 21039 36023
rect 21465 35989 21499 36023
rect 22477 35989 22511 36023
rect 25237 35989 25271 36023
rect 27445 35989 27479 36023
rect 29209 35989 29243 36023
rect 32229 35989 32263 36023
rect 5549 35785 5583 35819
rect 8309 35785 8343 35819
rect 19441 35785 19475 35819
rect 23765 35785 23799 35819
rect 25329 35785 25363 35819
rect 29561 35785 29595 35819
rect 30573 35785 30607 35819
rect 20729 35717 20763 35751
rect 24041 35717 24075 35751
rect 24593 35717 24627 35751
rect 24961 35717 24995 35751
rect 25881 35717 25915 35751
rect 29745 35717 29779 35751
rect 30389 35717 30423 35751
rect 5273 35649 5307 35683
rect 6561 35649 6595 35683
rect 13093 35649 13127 35683
rect 19625 35649 19659 35683
rect 20177 35649 20211 35683
rect 23673 35649 23707 35683
rect 23857 35649 23891 35683
rect 23949 35649 23983 35683
rect 24133 35649 24167 35683
rect 24409 35649 24443 35683
rect 24501 35649 24535 35683
rect 24777 35649 24811 35683
rect 24869 35649 24903 35683
rect 25145 35649 25179 35683
rect 26249 35649 26283 35683
rect 26525 35649 26559 35683
rect 26985 35649 27019 35683
rect 29929 35649 29963 35683
rect 30941 35649 30975 35683
rect 31125 35649 31159 35683
rect 31493 35649 31527 35683
rect 1409 35581 1443 35615
rect 4537 35581 4571 35615
rect 6101 35581 6135 35615
rect 6837 35581 6871 35615
rect 9873 35581 9907 35615
rect 10149 35581 10183 35615
rect 13369 35581 13403 35615
rect 19901 35581 19935 35615
rect 20361 35581 20395 35615
rect 25421 35581 25455 35615
rect 28733 35581 28767 35615
rect 30849 35581 30883 35615
rect 31033 35581 31067 35615
rect 31309 35581 31343 35615
rect 13185 35513 13219 35547
rect 21097 35513 21131 35547
rect 25605 35513 25639 35547
rect 30021 35513 30055 35547
rect 3893 35445 3927 35479
rect 4629 35445 4663 35479
rect 8401 35445 8435 35479
rect 13093 35445 13127 35479
rect 19809 35445 19843 35479
rect 19993 35445 20027 35479
rect 20545 35445 20579 35479
rect 20729 35445 20763 35479
rect 24225 35445 24259 35479
rect 26341 35445 26375 35479
rect 27248 35445 27282 35479
rect 30389 35445 30423 35479
rect 30665 35445 30699 35479
rect 31677 35445 31711 35479
rect 38485 35445 38519 35479
rect 6101 35241 6135 35275
rect 7205 35241 7239 35275
rect 8033 35241 8067 35275
rect 12541 35241 12575 35275
rect 13737 35241 13771 35275
rect 17785 35241 17819 35275
rect 20710 35241 20744 35275
rect 22201 35241 22235 35275
rect 24225 35241 24259 35275
rect 25237 35241 25271 35275
rect 27261 35241 27295 35275
rect 27445 35241 27479 35275
rect 30941 35241 30975 35275
rect 31953 35241 31987 35275
rect 15301 35173 15335 35207
rect 15577 35173 15611 35207
rect 18245 35173 18279 35207
rect 24041 35173 24075 35207
rect 28273 35173 28307 35207
rect 30757 35173 30791 35207
rect 2881 35105 2915 35139
rect 3341 35105 3375 35139
rect 6745 35105 6779 35139
rect 7757 35105 7791 35139
rect 8677 35105 8711 35139
rect 10793 35105 10827 35139
rect 15945 35105 15979 35139
rect 20453 35105 20487 35139
rect 22937 35105 22971 35139
rect 24869 35105 24903 35139
rect 24961 35105 24995 35139
rect 29653 35105 29687 35139
rect 33701 35105 33735 35139
rect 1409 35037 1443 35071
rect 3249 35037 3283 35071
rect 4077 35037 4111 35071
rect 4261 35037 4295 35071
rect 4353 35037 4387 35071
rect 6837 35037 6871 35071
rect 7205 35037 7239 35071
rect 7665 35037 7699 35071
rect 8125 35037 8159 35071
rect 13277 35037 13311 35071
rect 13461 35037 13495 35071
rect 14657 35037 14691 35071
rect 15117 35037 15151 35071
rect 15669 35037 15703 35071
rect 18061 35037 18095 35071
rect 18337 35037 18371 35071
rect 22661 35037 22695 35071
rect 22753 35037 22787 35071
rect 23765 35037 23799 35071
rect 24777 35037 24811 35071
rect 25237 35037 25271 35071
rect 25329 35037 25363 35071
rect 27537 35037 27571 35071
rect 27721 35037 27755 35071
rect 28089 35037 28123 35071
rect 28273 35037 28307 35071
rect 29561 35037 29595 35071
rect 29745 35037 29779 35071
rect 30205 35037 30239 35071
rect 30389 35037 30423 35071
rect 31217 35037 31251 35071
rect 4169 34969 4203 35003
rect 4629 34969 4663 35003
rect 11069 34969 11103 35003
rect 13737 34969 13771 35003
rect 14105 34969 14139 35003
rect 15393 34969 15427 35003
rect 17969 34969 18003 35003
rect 27077 34969 27111 35003
rect 27293 34969 27327 35003
rect 30925 34969 30959 35003
rect 31125 34969 31159 35003
rect 33425 34969 33459 35003
rect 7389 34901 7423 34935
rect 12633 34901 12667 34935
rect 13553 34901 13587 34935
rect 15669 34901 15703 34935
rect 16589 34901 16623 34935
rect 17601 34901 17635 34935
rect 17769 34901 17803 34935
rect 18337 34901 18371 34935
rect 22937 34901 22971 34935
rect 24409 34901 24443 34935
rect 25605 34901 25639 34935
rect 27537 34901 27571 34935
rect 30389 34901 30423 34935
rect 31861 34901 31895 34935
rect 38485 34901 38519 34935
rect 10977 34697 11011 34731
rect 13921 34697 13955 34731
rect 15945 34697 15979 34731
rect 17417 34697 17451 34731
rect 20170 34697 20204 34731
rect 21833 34697 21867 34731
rect 22477 34697 22511 34731
rect 25421 34697 25455 34731
rect 25513 34697 25547 34731
rect 28273 34697 28307 34731
rect 30849 34697 30883 34731
rect 31677 34697 31711 34731
rect 2881 34629 2915 34663
rect 4629 34629 4663 34663
rect 12449 34629 12483 34663
rect 15485 34629 15519 34663
rect 18889 34629 18923 34663
rect 20269 34629 20303 34663
rect 20361 34629 20395 34663
rect 22753 34629 22787 34663
rect 24593 34629 24627 34663
rect 25881 34629 25915 34663
rect 30757 34629 30791 34663
rect 31861 34629 31895 34663
rect 32137 34629 32171 34663
rect 5365 34561 5399 34595
rect 5917 34561 5951 34595
rect 9781 34561 9815 34595
rect 10149 34561 10183 34595
rect 10793 34561 10827 34595
rect 10885 34561 10919 34595
rect 11069 34561 11103 34595
rect 11161 34561 11195 34595
rect 11345 34561 11379 34595
rect 11897 34561 11931 34595
rect 15853 34561 15887 34595
rect 16037 34561 16071 34595
rect 16313 34561 16347 34595
rect 16497 34561 16531 34595
rect 17049 34561 17083 34595
rect 19993 34561 20027 34595
rect 20085 34561 20119 34595
rect 20637 34561 20671 34595
rect 22293 34561 22327 34595
rect 22661 34561 22695 34595
rect 22845 34561 22879 34595
rect 24869 34561 24903 34595
rect 25237 34561 25271 34595
rect 25605 34561 25639 34595
rect 26065 34561 26099 34595
rect 26157 34561 26191 34595
rect 28549 34561 28583 34595
rect 28733 34561 28767 34595
rect 28917 34561 28951 34595
rect 29101 34561 29135 34595
rect 29653 34561 29687 34595
rect 29837 34561 29871 34595
rect 30113 34561 30147 34595
rect 30297 34561 30331 34595
rect 30389 34561 30423 34595
rect 30481 34561 30515 34595
rect 31033 34561 31067 34595
rect 31493 34561 31527 34595
rect 31585 34561 31619 34595
rect 32321 34561 32355 34595
rect 32413 34561 32447 34595
rect 34069 34561 34103 34595
rect 2605 34493 2639 34527
rect 6193 34493 6227 34527
rect 9597 34493 9631 34527
rect 9965 34493 9999 34527
rect 10425 34493 10459 34527
rect 11805 34493 11839 34527
rect 12173 34493 12207 34527
rect 14013 34493 14047 34527
rect 15761 34493 15795 34527
rect 17141 34493 17175 34527
rect 19165 34493 19199 34527
rect 20361 34493 20395 34527
rect 20729 34493 20763 34527
rect 21281 34493 21315 34527
rect 22009 34493 22043 34527
rect 22109 34493 22143 34527
rect 22201 34493 22235 34527
rect 23121 34493 23155 34527
rect 25145 34493 25179 34527
rect 28457 34493 28491 34527
rect 28641 34493 28675 34527
rect 29561 34493 29595 34527
rect 29745 34493 29779 34527
rect 30021 34493 30055 34527
rect 31125 34493 31159 34527
rect 32137 34493 32171 34527
rect 32965 34493 32999 34527
rect 33241 34493 33275 34527
rect 10609 34425 10643 34459
rect 11529 34425 11563 34459
rect 16681 34425 16715 34459
rect 23029 34425 23063 34459
rect 31861 34425 31895 34459
rect 4353 34357 4387 34391
rect 10241 34357 10275 34391
rect 10333 34357 10367 34391
rect 11345 34357 11379 34391
rect 16497 34357 16531 34391
rect 20545 34357 20579 34391
rect 29009 34357 29043 34391
rect 31217 34357 31251 34391
rect 38485 34357 38519 34391
rect 5181 34153 5215 34187
rect 5641 34153 5675 34187
rect 6837 34153 6871 34187
rect 13093 34153 13127 34187
rect 13369 34153 13403 34187
rect 13553 34153 13587 34187
rect 15301 34153 15335 34187
rect 18521 34153 18555 34187
rect 29193 34153 29227 34187
rect 30849 34153 30883 34187
rect 5365 34085 5399 34119
rect 30481 34085 30515 34119
rect 3525 34017 3559 34051
rect 5089 34017 5123 34051
rect 10701 34017 10735 34051
rect 10977 34017 11011 34051
rect 11345 34017 11379 34051
rect 15945 34017 15979 34051
rect 16221 34017 16255 34051
rect 17785 34017 17819 34051
rect 19257 34017 19291 34051
rect 21741 34017 21775 34051
rect 21925 34017 21959 34051
rect 25421 34017 25455 34051
rect 27445 34017 27479 34051
rect 29837 34017 29871 34051
rect 32321 34017 32355 34051
rect 32597 34017 32631 34051
rect 3157 33949 3191 33983
rect 3341 33949 3375 33983
rect 3433 33949 3467 33983
rect 3617 33949 3651 33983
rect 3985 33949 4019 33983
rect 4537 33949 4571 33983
rect 4721 33949 4755 33983
rect 5181 33949 5215 33983
rect 6745 33949 6779 33983
rect 6929 33949 6963 33983
rect 15025 33949 15059 33983
rect 15117 33949 15151 33983
rect 18797 33949 18831 33983
rect 30481 33949 30515 33983
rect 30757 33949 30791 33983
rect 33241 33949 33275 33983
rect 5825 33881 5859 33915
rect 11621 33881 11655 33915
rect 13185 33881 13219 33915
rect 13401 33881 13435 33915
rect 18429 33881 18463 33915
rect 18521 33881 18555 33915
rect 19533 33881 19567 33915
rect 22201 33881 22235 33915
rect 27721 33881 27755 33915
rect 3249 33813 3283 33847
rect 5457 33813 5491 33847
rect 5625 33813 5659 33847
rect 7113 33813 7147 33847
rect 9229 33813 9263 33847
rect 17693 33813 17727 33847
rect 18705 33813 18739 33847
rect 21005 33813 21039 33847
rect 21189 33813 21223 33847
rect 23673 33813 23707 33847
rect 24777 33813 24811 33847
rect 30389 33813 30423 33847
rect 30665 33813 30699 33847
rect 6637 33609 6671 33643
rect 11253 33609 11287 33643
rect 21649 33609 21683 33643
rect 22201 33609 22235 33643
rect 27537 33609 27571 33643
rect 28365 33609 28399 33643
rect 29285 33609 29319 33643
rect 2513 33541 2547 33575
rect 6837 33541 6871 33575
rect 9229 33541 9263 33575
rect 10853 33541 10887 33575
rect 11069 33541 11103 33575
rect 20177 33541 20211 33575
rect 23213 33541 23247 33575
rect 30757 33541 30791 33575
rect 4353 33473 4387 33507
rect 4629 33473 4663 33507
rect 4721 33473 4755 33507
rect 4905 33473 4939 33507
rect 5181 33473 5215 33507
rect 7113 33473 7147 33507
rect 7297 33473 7331 33507
rect 11161 33473 11195 33507
rect 11345 33473 11379 33507
rect 15577 33473 15611 33507
rect 18889 33473 18923 33507
rect 22017 33473 22051 33507
rect 22293 33473 22327 33507
rect 22385 33473 22419 33507
rect 23397 33473 23431 33507
rect 23489 33473 23523 33507
rect 23673 33473 23707 33507
rect 24869 33473 24903 33507
rect 27261 33473 27295 33507
rect 27445 33473 27479 33507
rect 27813 33473 27847 33507
rect 27905 33473 27939 33507
rect 27997 33473 28031 33507
rect 28181 33473 28215 33507
rect 28273 33473 28307 33507
rect 28457 33473 28491 33507
rect 29193 33473 29227 33507
rect 33241 33473 33275 33507
rect 2237 33405 2271 33439
rect 3985 33405 4019 33439
rect 4537 33405 4571 33439
rect 5733 33405 5767 33439
rect 7757 33405 7791 33439
rect 9505 33405 9539 33439
rect 10057 33405 10091 33439
rect 10609 33405 10643 33439
rect 15761 33405 15795 33439
rect 19625 33405 19659 33439
rect 19901 33405 19935 33439
rect 23765 33405 23799 33439
rect 25145 33405 25179 33439
rect 28549 33405 28583 33439
rect 31033 33405 31067 33439
rect 31677 33405 31711 33439
rect 33517 33405 33551 33439
rect 34989 33405 35023 33439
rect 35633 33405 35667 33439
rect 35081 33337 35115 33371
rect 38485 33337 38519 33371
rect 4169 33269 4203 33303
rect 4905 33269 4939 33303
rect 6469 33269 6503 33303
rect 6653 33269 6687 33303
rect 6929 33269 6963 33303
rect 10701 33269 10735 33303
rect 10885 33269 10919 33303
rect 15393 33269 15427 33303
rect 18705 33269 18739 33303
rect 21833 33269 21867 33303
rect 23581 33269 23615 33303
rect 26617 33269 26651 33303
rect 27077 33269 27111 33303
rect 31125 33269 31159 33303
rect 9689 33065 9723 33099
rect 10609 33065 10643 33099
rect 10977 33065 11011 33099
rect 11161 33065 11195 33099
rect 17049 33065 17083 33099
rect 18153 33065 18187 33099
rect 19901 33065 19935 33099
rect 22017 33065 22051 33099
rect 22201 33065 22235 33099
rect 24409 33065 24443 33099
rect 26249 33065 26283 33099
rect 27997 33065 28031 33099
rect 30665 33065 30699 33099
rect 33609 33065 33643 33099
rect 15209 32997 15243 33031
rect 16681 32997 16715 33031
rect 17969 32997 18003 33031
rect 20085 32997 20119 33031
rect 34529 32997 34563 33031
rect 3893 32929 3927 32963
rect 5733 32929 5767 32963
rect 6009 32929 6043 32963
rect 8953 32929 8987 32963
rect 9597 32929 9631 32963
rect 10149 32929 10183 32963
rect 20361 32929 20395 32963
rect 26157 32929 26191 32963
rect 26893 32929 26927 32963
rect 30849 32929 30883 32963
rect 31769 32929 31803 32963
rect 33977 32929 34011 32963
rect 34161 32929 34195 32963
rect 34897 32929 34931 32963
rect 35173 32929 35207 32963
rect 3433 32861 3467 32895
rect 3617 32861 3651 32895
rect 7757 32861 7791 32895
rect 7849 32861 7883 32895
rect 8401 32861 8435 32895
rect 8585 32861 8619 32895
rect 9873 32861 9907 32895
rect 10057 32861 10091 32895
rect 10701 32861 10735 32895
rect 10885 32861 10919 32895
rect 11437 32861 11471 32895
rect 11621 32861 11655 32895
rect 15025 32861 15059 32895
rect 15301 32861 15335 32895
rect 15761 32861 15795 32895
rect 16313 32861 16347 32895
rect 17509 32861 17543 32895
rect 17601 32861 17635 32895
rect 17693 32861 17727 32895
rect 17785 32861 17819 32895
rect 19349 32861 19383 32895
rect 22385 32861 22419 32895
rect 27077 32861 27111 32895
rect 27261 32861 27295 32895
rect 27445 32861 27479 32895
rect 27721 32861 27755 32895
rect 28733 32861 28767 32895
rect 29009 32861 29043 32895
rect 29561 32861 29595 32895
rect 30757 32861 30791 32895
rect 33885 32861 33919 32895
rect 34253 32861 34287 32895
rect 34345 32861 34379 32895
rect 34529 32861 34563 32895
rect 3525 32793 3559 32827
rect 4169 32793 4203 32827
rect 8493 32793 8527 32827
rect 10241 32793 10275 32827
rect 10425 32793 10459 32827
rect 10793 32793 10827 32827
rect 11345 32793 11379 32827
rect 12449 32793 12483 32827
rect 17049 32793 17083 32827
rect 18337 32793 18371 32827
rect 21833 32793 21867 32827
rect 25881 32793 25915 32827
rect 26617 32793 26651 32827
rect 27629 32793 27663 32827
rect 30297 32793 30331 32827
rect 32045 32793 32079 32827
rect 33609 32793 33643 32827
rect 33977 32793 34011 32827
rect 5641 32725 5675 32759
rect 7481 32725 7515 32759
rect 7573 32725 7607 32759
rect 11145 32725 11179 32759
rect 14841 32725 14875 32759
rect 17233 32725 17267 32759
rect 17325 32725 17359 32759
rect 18137 32725 18171 32759
rect 22033 32725 22067 32759
rect 26709 32725 26743 32759
rect 27169 32725 27203 32759
rect 27813 32725 27847 32759
rect 28181 32725 28215 32759
rect 33517 32725 33551 32759
rect 33793 32725 33827 32759
rect 36645 32725 36679 32759
rect 4011 32521 4045 32555
rect 4905 32521 4939 32555
rect 6929 32521 6963 32555
rect 7113 32521 7147 32555
rect 11805 32521 11839 32555
rect 14197 32521 14231 32555
rect 16129 32521 16163 32555
rect 24159 32521 24193 32555
rect 25605 32521 25639 32555
rect 25789 32521 25823 32555
rect 28273 32521 28307 32555
rect 32137 32521 32171 32555
rect 32305 32521 32339 32555
rect 33517 32521 33551 32555
rect 33885 32521 33919 32555
rect 34621 32521 34655 32555
rect 3801 32453 3835 32487
rect 14657 32453 14691 32487
rect 16957 32453 16991 32487
rect 18521 32453 18555 32487
rect 18737 32453 18771 32487
rect 23949 32453 23983 32487
rect 32505 32453 32539 32487
rect 33793 32453 33827 32487
rect 6561 32385 6595 32419
rect 6653 32385 6687 32419
rect 6745 32385 6779 32419
rect 7205 32385 7239 32419
rect 9597 32385 9631 32419
rect 13553 32385 13587 32419
rect 14105 32385 14139 32419
rect 14289 32385 14323 32419
rect 14381 32385 14415 32419
rect 16681 32385 16715 32419
rect 18981 32385 19015 32419
rect 19165 32385 19199 32419
rect 22109 32385 22143 32419
rect 24593 32385 24627 32419
rect 24685 32385 24719 32419
rect 24961 32385 24995 32419
rect 25054 32385 25088 32419
rect 25237 32385 25271 32419
rect 25329 32385 25363 32419
rect 25467 32385 25501 32419
rect 25697 32385 25731 32419
rect 25881 32385 25915 32419
rect 27169 32385 27203 32419
rect 27537 32385 27571 32419
rect 27721 32385 27755 32419
rect 27813 32385 27847 32419
rect 27905 32385 27939 32419
rect 30021 32385 30055 32419
rect 31401 32385 31435 32419
rect 31493 32385 31527 32419
rect 31769 32385 31803 32419
rect 33057 32385 33091 32419
rect 33333 32385 33367 32419
rect 33517 32385 33551 32419
rect 33609 32385 33643 32419
rect 34069 32385 34103 32419
rect 34253 32385 34287 32419
rect 34345 32385 34379 32419
rect 4353 32317 4387 32351
rect 4997 32317 5031 32351
rect 9873 32317 9907 32351
rect 13277 32317 13311 32351
rect 16497 32317 16531 32351
rect 22385 32317 22419 32351
rect 23857 32317 23891 32351
rect 29745 32317 29779 32351
rect 31033 32317 31067 32351
rect 31585 32317 31619 32351
rect 33149 32317 33183 32351
rect 33241 32317 33275 32351
rect 34621 32317 34655 32351
rect 4169 32249 4203 32283
rect 5273 32249 5307 32283
rect 19349 32249 19383 32283
rect 24317 32249 24351 32283
rect 28181 32249 28215 32283
rect 34437 32249 34471 32283
rect 3985 32181 4019 32215
rect 5457 32181 5491 32215
rect 11345 32181 11379 32215
rect 18429 32181 18463 32215
rect 18705 32181 18739 32215
rect 18889 32181 18923 32215
rect 24133 32181 24167 32215
rect 24685 32181 24719 32215
rect 27353 32181 27387 32215
rect 31217 32181 31251 32215
rect 32321 32181 32355 32215
rect 32873 32181 32907 32215
rect 4721 31977 4755 32011
rect 6193 31977 6227 32011
rect 10241 31977 10275 32011
rect 12541 31977 12575 32011
rect 14841 31977 14875 32011
rect 15945 31977 15979 32011
rect 18613 31977 18647 32011
rect 18981 31977 19015 32011
rect 25973 31977 26007 32011
rect 27077 31977 27111 32011
rect 28549 31977 28583 32011
rect 33149 31977 33183 32011
rect 3617 31909 3651 31943
rect 6285 31909 6319 31943
rect 10333 31909 10367 31943
rect 10609 31909 10643 31943
rect 17141 31909 17175 31943
rect 18245 31909 18279 31943
rect 18797 31909 18831 31943
rect 22569 31909 22603 31943
rect 27169 31909 27203 31943
rect 1869 31841 1903 31875
rect 2145 31841 2179 31875
rect 3985 31841 4019 31875
rect 4997 31841 5031 31875
rect 5549 31841 5583 31875
rect 6034 31841 6068 31875
rect 6561 31841 6595 31875
rect 6653 31841 6687 31875
rect 10149 31841 10183 31875
rect 11529 31841 11563 31875
rect 17877 31841 17911 31875
rect 19257 31841 19291 31875
rect 20729 31841 20763 31875
rect 23305 31841 23339 31875
rect 27905 31841 27939 31875
rect 30389 31841 30423 31875
rect 30665 31841 30699 31875
rect 32137 31841 32171 31875
rect 4629 31773 4663 31807
rect 5089 31773 5123 31807
rect 6469 31773 6503 31807
rect 6745 31773 6779 31807
rect 7113 31773 7147 31807
rect 8125 31773 8159 31807
rect 10425 31773 10459 31807
rect 10885 31773 10919 31807
rect 12265 31773 12299 31807
rect 12449 31773 12483 31807
rect 12633 31773 12667 31807
rect 14657 31773 14691 31807
rect 14933 31773 14967 31807
rect 15025 31773 15059 31807
rect 15577 31773 15611 31807
rect 17601 31773 17635 31807
rect 18889 31773 18923 31807
rect 19073 31773 19107 31807
rect 21005 31773 21039 31807
rect 21189 31773 21223 31807
rect 23949 31773 23983 31807
rect 24961 31773 24995 31807
rect 25329 31773 25363 31807
rect 26525 31773 26559 31807
rect 26709 31773 26743 31807
rect 26801 31773 26835 31807
rect 27445 31773 27479 31807
rect 27537 31773 27571 31807
rect 27650 31773 27684 31807
rect 27813 31773 27847 31807
rect 28089 31773 28123 31807
rect 28365 31773 28399 31807
rect 28641 31773 28675 31807
rect 32413 31773 32447 31807
rect 32965 31773 32999 31807
rect 33057 31773 33091 31807
rect 35541 31773 35575 31807
rect 36185 31773 36219 31807
rect 38485 31773 38519 31807
rect 7297 31705 7331 31739
rect 7481 31705 7515 31739
rect 10609 31705 10643 31739
rect 10977 31705 11011 31739
rect 15761 31705 15795 31739
rect 15961 31705 15995 31739
rect 17141 31705 17175 31739
rect 17693 31705 17727 31739
rect 21456 31705 21490 31739
rect 26617 31705 26651 31739
rect 27077 31705 27111 31739
rect 5825 31637 5859 31671
rect 5917 31637 5951 31671
rect 7573 31637 7607 31671
rect 10793 31637 10827 31671
rect 11713 31637 11747 31671
rect 14473 31637 14507 31671
rect 16129 31637 16163 31671
rect 18613 31637 18647 31671
rect 22661 31637 22695 31671
rect 23397 31637 23431 31671
rect 24409 31637 24443 31671
rect 26893 31637 26927 31671
rect 28273 31637 28307 31671
rect 6745 31433 6779 31467
rect 7757 31433 7791 31467
rect 12081 31433 12115 31467
rect 14841 31433 14875 31467
rect 15301 31433 15335 31467
rect 17049 31433 17083 31467
rect 18153 31433 18187 31467
rect 18613 31433 18647 31467
rect 22477 31433 22511 31467
rect 24317 31433 24351 31467
rect 25053 31433 25087 31467
rect 29101 31433 29135 31467
rect 36645 31433 36679 31467
rect 6561 31365 6595 31399
rect 17385 31365 17419 31399
rect 17601 31365 17635 31399
rect 20177 31365 20211 31399
rect 22845 31365 22879 31399
rect 27629 31365 27663 31399
rect 35173 31365 35207 31399
rect 3341 31297 3375 31331
rect 5825 31297 5859 31331
rect 6653 31297 6687 31331
rect 7297 31297 7331 31331
rect 10977 31297 11011 31331
rect 11713 31297 11747 31331
rect 13093 31297 13127 31331
rect 15209 31297 15243 31331
rect 15393 31297 15427 31331
rect 16037 31297 16071 31331
rect 16221 31297 16255 31331
rect 16313 31297 16347 31331
rect 16957 31297 16991 31331
rect 17141 31297 17175 31331
rect 17969 31297 18003 31331
rect 18245 31297 18279 31331
rect 18429 31297 18463 31331
rect 20453 31297 20487 31331
rect 21833 31297 21867 31331
rect 22017 31297 22051 31331
rect 22109 31297 22143 31331
rect 22201 31297 22235 31331
rect 22569 31297 22603 31331
rect 24501 31297 24535 31331
rect 24593 31297 24627 31331
rect 27353 31297 27387 31331
rect 32781 31297 32815 31331
rect 32965 31297 32999 31331
rect 3617 31229 3651 31263
rect 5089 31229 5123 31263
rect 7389 31229 7423 31263
rect 9229 31229 9263 31263
rect 9505 31229 9539 31263
rect 10701 31229 10735 31263
rect 11805 31229 11839 31263
rect 13369 31229 13403 31263
rect 17785 31229 17819 31263
rect 18705 31229 18739 31263
rect 26525 31229 26559 31263
rect 26801 31229 26835 31263
rect 33977 31229 34011 31263
rect 34253 31229 34287 31263
rect 34897 31229 34931 31263
rect 5181 31161 5215 31195
rect 6929 31161 6963 31195
rect 7665 31161 7699 31195
rect 6377 31093 6411 31127
rect 10793 31093 10827 31127
rect 10885 31093 10919 31127
rect 16037 31093 16071 31127
rect 17233 31093 17267 31127
rect 17417 31093 17451 31127
rect 24777 31093 24811 31127
rect 29929 31093 29963 31127
rect 30481 31093 30515 31127
rect 32597 31093 32631 31127
rect 32965 31093 32999 31127
rect 3893 30889 3927 30923
rect 6745 30889 6779 30923
rect 7297 30889 7331 30923
rect 12449 30889 12483 30923
rect 15945 30889 15979 30923
rect 16129 30889 16163 30923
rect 23581 30889 23615 30923
rect 26985 30889 27019 30923
rect 32229 30889 32263 30923
rect 33425 30889 33459 30923
rect 33793 30889 33827 30923
rect 33977 30889 34011 30923
rect 35081 30889 35115 30923
rect 13921 30821 13955 30855
rect 15485 30821 15519 30855
rect 22477 30821 22511 30855
rect 26157 30821 26191 30855
rect 34713 30821 34747 30855
rect 5273 30753 5307 30787
rect 7481 30753 7515 30787
rect 9873 30753 9907 30787
rect 11621 30753 11655 30787
rect 12265 30753 12299 30787
rect 12817 30753 12851 30787
rect 14657 30753 14691 30787
rect 15209 30753 15243 30787
rect 17325 30753 17359 30787
rect 21097 30753 21131 30787
rect 24225 30753 24259 30787
rect 26341 30753 26375 30787
rect 29653 30753 29687 30787
rect 31401 30753 31435 30787
rect 32505 30753 32539 30787
rect 33517 30753 33551 30787
rect 34345 30753 34379 30787
rect 34529 30753 34563 30787
rect 3893 30685 3927 30719
rect 4077 30685 4111 30719
rect 4445 30685 4479 30719
rect 4629 30685 4663 30719
rect 4997 30685 5031 30719
rect 7205 30685 7239 30719
rect 7389 30685 7423 30719
rect 7665 30685 7699 30719
rect 12633 30685 12667 30719
rect 13369 30685 13403 30719
rect 13553 30685 13587 30719
rect 13645 30685 13679 30719
rect 13737 30685 13771 30719
rect 14381 30685 14415 30719
rect 14565 30685 14599 30719
rect 14841 30685 14875 30719
rect 15761 30685 15795 30719
rect 16037 30685 16071 30719
rect 16681 30685 16715 30719
rect 17969 30685 18003 30719
rect 18153 30685 18187 30719
rect 23765 30685 23799 30719
rect 23857 30685 23891 30719
rect 23949 30685 23983 30719
rect 24067 30685 24101 30719
rect 25421 30685 25455 30719
rect 25605 30685 25639 30719
rect 25789 30685 25823 30719
rect 25973 30685 26007 30719
rect 32321 30685 32355 30719
rect 32413 30685 32447 30719
rect 32781 30685 32815 30719
rect 32873 30685 32907 30719
rect 32965 30685 32999 30719
rect 33149 30685 33183 30719
rect 33425 30685 33459 30719
rect 33701 30685 33735 30719
rect 34253 30685 34287 30719
rect 35357 30685 35391 30719
rect 38485 30685 38519 30719
rect 4537 30617 4571 30651
rect 10149 30617 10183 30651
rect 13461 30617 13495 30651
rect 13921 30617 13955 30651
rect 14197 30617 14231 30651
rect 15326 30617 15360 30651
rect 16313 30617 16347 30651
rect 16497 30617 16531 30651
rect 17509 30617 17543 30651
rect 17877 30617 17911 30651
rect 18337 30617 18371 30651
rect 21364 30617 21398 30651
rect 22753 30617 22787 30651
rect 24409 30617 24443 30651
rect 24593 30617 24627 30651
rect 24777 30617 24811 30651
rect 25881 30617 25915 30651
rect 29929 30617 29963 30651
rect 32137 30617 32171 30651
rect 34161 30617 34195 30651
rect 35633 30617 35667 30651
rect 7849 30549 7883 30583
rect 11713 30549 11747 30583
rect 15117 30549 15151 30583
rect 15577 30549 15611 30583
rect 18429 30549 18463 30583
rect 22845 30549 22879 30583
rect 24869 30549 24903 30583
rect 33241 30549 33275 30583
rect 33956 30549 33990 30583
rect 34529 30549 34563 30583
rect 35081 30549 35115 30583
rect 35265 30549 35299 30583
rect 37105 30549 37139 30583
rect 7573 30345 7607 30379
rect 14841 30345 14875 30379
rect 16129 30345 16163 30379
rect 17325 30345 17359 30379
rect 20729 30345 20763 30379
rect 21281 30345 21315 30379
rect 35449 30345 35483 30379
rect 5181 30277 5215 30311
rect 9045 30277 9079 30311
rect 10241 30277 10275 30311
rect 15577 30277 15611 30311
rect 16497 30277 16531 30311
rect 17049 30277 17083 30311
rect 22109 30277 22143 30311
rect 23305 30277 23339 30311
rect 24409 30277 24443 30311
rect 30389 30277 30423 30311
rect 34529 30277 34563 30311
rect 4077 30209 4111 30243
rect 5365 30209 5399 30243
rect 5549 30209 5583 30243
rect 6837 30209 6871 30243
rect 9321 30209 9355 30243
rect 9597 30209 9631 30243
rect 9781 30209 9815 30243
rect 11069 30209 11103 30243
rect 11253 30209 11287 30243
rect 12357 30209 12391 30243
rect 14381 30209 14415 30243
rect 15761 30209 15795 30243
rect 16037 30209 16071 30243
rect 16313 30209 16347 30243
rect 19073 30209 19107 30243
rect 19441 30209 19475 30243
rect 19625 30209 19659 30243
rect 20269 30209 20303 30243
rect 20361 30209 20395 30243
rect 20913 30209 20947 30243
rect 21465 30209 21499 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 22201 30209 22235 30243
rect 23489 30209 23523 30243
rect 23857 30209 23891 30243
rect 24041 30209 24075 30243
rect 24133 30209 24167 30243
rect 29653 30209 29687 30243
rect 30113 30209 30147 30243
rect 32505 30209 32539 30243
rect 32689 30209 32723 30243
rect 32781 30209 32815 30243
rect 32965 30209 32999 30243
rect 34253 30209 34287 30243
rect 34345 30209 34379 30243
rect 35265 30209 35299 30243
rect 35725 30209 35759 30243
rect 35817 30209 35851 30243
rect 10885 30141 10919 30175
rect 12633 30141 12667 30175
rect 14197 30141 14231 30175
rect 14565 30141 14599 30175
rect 14657 30141 14691 30175
rect 15393 30141 15427 30175
rect 15945 30141 15979 30175
rect 16681 30141 16715 30175
rect 18797 30141 18831 30175
rect 21649 30141 21683 30175
rect 23673 30141 23707 30175
rect 23765 30141 23799 30175
rect 26525 30141 26559 30175
rect 26985 30141 27019 30175
rect 35633 30141 35667 30175
rect 35909 30141 35943 30175
rect 1409 30073 1443 30107
rect 3893 30073 3927 30107
rect 11069 30073 11103 30107
rect 14105 30073 14139 30107
rect 17233 30073 17267 30107
rect 22385 30073 22419 30107
rect 31861 30073 31895 30107
rect 32597 30073 32631 30107
rect 34529 30073 34563 30107
rect 9689 30005 9723 30039
rect 17049 30005 17083 30039
rect 19257 30005 19291 30039
rect 20545 30005 20579 30039
rect 25881 30005 25915 30039
rect 25973 30005 26007 30039
rect 27629 30005 27663 30039
rect 29929 30005 29963 30039
rect 32229 30005 32263 30039
rect 12725 29801 12759 29835
rect 14381 29801 14415 29835
rect 17233 29801 17267 29835
rect 17325 29801 17359 29835
rect 17509 29801 17543 29835
rect 19349 29801 19383 29835
rect 24133 29801 24167 29835
rect 25973 29801 26007 29835
rect 30481 29801 30515 29835
rect 31125 29801 31159 29835
rect 32781 29801 32815 29835
rect 34345 29801 34379 29835
rect 11253 29733 11287 29767
rect 11529 29733 11563 29767
rect 18889 29733 18923 29767
rect 26065 29733 26099 29767
rect 28549 29733 28583 29767
rect 36737 29733 36771 29767
rect 4537 29665 4571 29699
rect 4997 29665 5031 29699
rect 7941 29665 7975 29699
rect 9229 29665 9263 29699
rect 11345 29665 11379 29699
rect 15025 29665 15059 29699
rect 15761 29665 15795 29699
rect 25513 29665 25547 29699
rect 27537 29665 27571 29699
rect 27813 29665 27847 29699
rect 28917 29665 28951 29699
rect 29101 29665 29135 29699
rect 34713 29665 34747 29699
rect 1409 29597 1443 29631
rect 3801 29597 3835 29631
rect 4905 29597 4939 29631
rect 5365 29597 5399 29631
rect 6009 29597 6043 29631
rect 7573 29597 7607 29631
rect 7849 29597 7883 29631
rect 8677 29597 8711 29631
rect 8953 29597 8987 29631
rect 10977 29597 11011 29631
rect 11621 29597 11655 29631
rect 15485 29597 15519 29631
rect 18797 29597 18831 29631
rect 19533 29597 19567 29631
rect 19625 29597 19659 29631
rect 19901 29597 19935 29631
rect 21106 29597 21140 29631
rect 21373 29597 21407 29631
rect 21741 29597 21775 29631
rect 23489 29597 23523 29631
rect 23949 29597 23983 29631
rect 24409 29597 24443 29631
rect 25237 29597 25271 29631
rect 25421 29597 25455 29631
rect 25605 29597 25639 29631
rect 25789 29597 25823 29631
rect 28825 29597 28859 29631
rect 29193 29597 29227 29631
rect 30113 29597 30147 29631
rect 30849 29597 30883 29631
rect 32965 29597 32999 29631
rect 33057 29597 33091 29631
rect 33241 29597 33275 29631
rect 33333 29597 33367 29631
rect 33977 29597 34011 29631
rect 36737 29597 36771 29631
rect 37013 29597 37047 29631
rect 3525 29529 3559 29563
rect 6377 29529 6411 29563
rect 7205 29529 7239 29563
rect 11253 29529 11287 29563
rect 12449 29529 12483 29563
rect 17493 29529 17527 29563
rect 17693 29529 17727 29563
rect 19717 29529 19751 29563
rect 22008 29529 22042 29563
rect 23305 29529 23339 29563
rect 23765 29529 23799 29563
rect 28549 29529 28583 29563
rect 28733 29529 28767 29563
rect 29561 29529 29595 29563
rect 31309 29529 31343 29563
rect 34989 29529 35023 29563
rect 3433 29461 3467 29495
rect 4445 29461 4479 29495
rect 7389 29461 7423 29495
rect 7757 29461 7791 29495
rect 8125 29461 8159 29495
rect 10701 29461 10735 29495
rect 11069 29461 11103 29495
rect 11345 29461 11379 29495
rect 13001 29461 13035 29495
rect 19993 29461 20027 29495
rect 23121 29461 23155 29495
rect 23673 29461 23707 29495
rect 25053 29461 25087 29495
rect 28917 29461 28951 29495
rect 30297 29461 30331 29495
rect 30481 29461 30515 29495
rect 30941 29461 30975 29495
rect 31109 29461 31143 29495
rect 34345 29461 34379 29495
rect 34529 29461 34563 29495
rect 36461 29461 36495 29495
rect 36921 29461 36955 29495
rect 8953 29257 8987 29291
rect 11529 29257 11563 29291
rect 12633 29257 12667 29291
rect 14841 29257 14875 29291
rect 20269 29257 20303 29291
rect 20361 29257 20395 29291
rect 21097 29257 21131 29291
rect 26525 29257 26559 29291
rect 29745 29257 29779 29291
rect 32689 29257 32723 29291
rect 33057 29257 33091 29291
rect 33885 29257 33919 29291
rect 34529 29257 34563 29291
rect 7113 29189 7147 29223
rect 12265 29189 12299 29223
rect 12465 29189 12499 29223
rect 18337 29189 18371 29223
rect 20637 29189 20671 29223
rect 22017 29189 22051 29223
rect 22109 29189 22143 29223
rect 23397 29189 23431 29223
rect 25329 29189 25363 29223
rect 25697 29189 25731 29223
rect 28273 29189 28307 29223
rect 30481 29189 30515 29223
rect 33517 29189 33551 29223
rect 33717 29189 33751 29223
rect 36461 29189 36495 29223
rect 3985 29121 4019 29155
rect 4077 29121 4111 29155
rect 4261 29121 4295 29155
rect 4445 29121 4479 29155
rect 6837 29121 6871 29155
rect 9045 29121 9079 29155
rect 9413 29121 9447 29155
rect 10609 29121 10643 29155
rect 12173 29121 12207 29155
rect 15209 29121 15243 29155
rect 18889 29121 18923 29155
rect 19156 29121 19190 29155
rect 20545 29121 20579 29155
rect 20729 29121 20763 29155
rect 20913 29121 20947 29155
rect 21189 29121 21223 29155
rect 21833 29121 21867 29155
rect 22201 29121 22235 29155
rect 22661 29121 22695 29155
rect 23581 29121 23615 29155
rect 30205 29121 30239 29155
rect 32781 29121 32815 29155
rect 34345 29121 34379 29155
rect 34621 29121 34655 29155
rect 36645 29121 36679 29155
rect 36921 29121 36955 29155
rect 37105 29121 37139 29155
rect 37473 29121 37507 29155
rect 1409 29053 1443 29087
rect 2237 29053 2271 29087
rect 3709 29053 3743 29087
rect 4721 29053 4755 29087
rect 9505 29053 9539 29087
rect 9873 29053 9907 29087
rect 11253 29053 11287 29087
rect 13093 29053 13127 29087
rect 13369 29053 13403 29087
rect 22845 29053 22879 29087
rect 23765 29053 23799 29087
rect 25605 29053 25639 29087
rect 26341 29053 26375 29087
rect 27537 29053 27571 29087
rect 27997 29053 28031 29087
rect 32413 29053 32447 29087
rect 32505 29053 32539 29087
rect 32873 29053 32907 29087
rect 34069 29053 34103 29087
rect 34161 29053 34195 29087
rect 34253 29053 34287 29087
rect 35449 29053 35483 29087
rect 37381 29053 37415 29087
rect 8585 28985 8619 29019
rect 9781 28985 9815 29019
rect 18153 28985 18187 29019
rect 21465 28985 21499 29019
rect 22385 28985 22419 29019
rect 22477 28985 22511 29019
rect 23857 28985 23891 29019
rect 4077 28917 4111 28951
rect 6193 28917 6227 28951
rect 10517 28917 10551 28951
rect 12409 28917 12443 28951
rect 26985 28917 27019 28951
rect 31953 28917 31987 28951
rect 33701 28917 33735 28951
rect 36829 28917 36863 28951
rect 37013 28917 37047 28951
rect 37749 28917 37783 28951
rect 3157 28713 3191 28747
rect 3985 28713 4019 28747
rect 7389 28713 7423 28747
rect 7573 28713 7607 28747
rect 11069 28713 11103 28747
rect 12909 28713 12943 28747
rect 21833 28713 21867 28747
rect 26065 28713 26099 28747
rect 30389 28713 30423 28747
rect 31309 28713 31343 28747
rect 34529 28713 34563 28747
rect 34805 28713 34839 28747
rect 34989 28713 35023 28747
rect 36001 28713 36035 28747
rect 24685 28645 24719 28679
rect 33701 28645 33735 28679
rect 4813 28577 4847 28611
rect 5089 28577 5123 28611
rect 6561 28577 6595 28611
rect 7205 28577 7239 28611
rect 8401 28577 8435 28611
rect 9321 28577 9355 28611
rect 11437 28577 11471 28611
rect 13645 28577 13679 28611
rect 15209 28577 15243 28611
rect 16037 28577 16071 28611
rect 23949 28577 23983 28611
rect 27537 28577 27571 28611
rect 27905 28577 27939 28611
rect 29653 28577 29687 28611
rect 30113 28577 30147 28611
rect 30849 28577 30883 28611
rect 32781 28577 32815 28611
rect 33517 28577 33551 28611
rect 34253 28577 34287 28611
rect 35449 28577 35483 28611
rect 35909 28577 35943 28611
rect 36461 28577 36495 28611
rect 36829 28577 36863 28611
rect 2973 28509 3007 28543
rect 3157 28509 3191 28543
rect 3341 28509 3375 28543
rect 3433 28509 3467 28543
rect 3801 28509 3835 28543
rect 3985 28509 4019 28543
rect 4077 28509 4111 28543
rect 4721 28509 4755 28543
rect 7941 28509 7975 28543
rect 11161 28509 11195 28543
rect 17049 28509 17083 28543
rect 21741 28509 21775 28543
rect 22385 28509 22419 28543
rect 22569 28509 22603 28543
rect 22661 28509 22695 28543
rect 22753 28509 22787 28543
rect 23397 28509 23431 28543
rect 24501 28509 24535 28543
rect 24961 28509 24995 28543
rect 27813 28509 27847 28543
rect 28457 28509 28491 28543
rect 28917 28509 28951 28543
rect 29009 28509 29043 28543
rect 29101 28509 29135 28543
rect 29285 28509 29319 28543
rect 29745 28509 29779 28543
rect 29929 28509 29963 28543
rect 30021 28509 30055 28543
rect 30205 28509 30239 28543
rect 30665 28509 30699 28543
rect 30941 28509 30975 28543
rect 33241 28509 33275 28543
rect 33793 28509 33827 28543
rect 34069 28509 34103 28543
rect 35541 28509 35575 28543
rect 36185 28509 36219 28543
rect 36277 28509 36311 28543
rect 36369 28509 36403 28543
rect 37013 28509 37047 28543
rect 37473 28509 37507 28543
rect 37749 28509 37783 28543
rect 37933 28509 37967 28543
rect 7573 28441 7607 28475
rect 8033 28441 8067 28475
rect 8217 28441 8251 28475
rect 9597 28441 9631 28475
rect 13461 28441 13495 28475
rect 14381 28441 14415 28475
rect 17325 28441 17359 28475
rect 19073 28441 19107 28475
rect 25697 28441 25731 28475
rect 31125 28441 31159 28475
rect 33885 28441 33919 28475
rect 34973 28441 35007 28475
rect 35173 28441 35207 28475
rect 37197 28441 37231 28475
rect 3617 28373 3651 28407
rect 6653 28373 6687 28407
rect 13001 28373 13035 28407
rect 13369 28373 13403 28407
rect 14197 28373 14231 28407
rect 15393 28373 15427 28407
rect 15761 28373 15795 28407
rect 15853 28373 15887 28407
rect 23029 28373 23063 28407
rect 28641 28373 28675 28407
rect 30481 28373 30515 28407
rect 33057 28373 33091 28407
rect 33149 28373 33183 28407
rect 33517 28373 33551 28407
rect 35265 28373 35299 28407
rect 37289 28373 37323 28407
rect 4905 28169 4939 28203
rect 10425 28169 10459 28203
rect 16037 28169 16071 28203
rect 17601 28169 17635 28203
rect 17969 28169 18003 28203
rect 20269 28169 20303 28203
rect 21373 28169 21407 28203
rect 23949 28169 23983 28203
rect 25973 28169 26007 28203
rect 29745 28169 29779 28203
rect 37933 28169 37967 28203
rect 2145 28101 2179 28135
rect 5365 28101 5399 28135
rect 5609 28101 5643 28135
rect 5825 28101 5859 28135
rect 7021 28101 7055 28135
rect 19717 28101 19751 28135
rect 22017 28101 22051 28135
rect 28273 28101 28307 28135
rect 30205 28101 30239 28135
rect 37565 28101 37599 28135
rect 37657 28101 37691 28135
rect 4261 28033 4295 28067
rect 4445 28033 4479 28067
rect 4537 28033 4571 28067
rect 4721 28033 4755 28067
rect 4813 28033 4847 28067
rect 4997 28033 5031 28067
rect 5089 28033 5123 28067
rect 5181 28033 5215 28067
rect 6745 28033 6779 28067
rect 7297 28033 7331 28067
rect 7573 28033 7607 28067
rect 10425 28033 10459 28067
rect 10609 28033 10643 28067
rect 12081 28033 12115 28067
rect 15761 28033 15795 28067
rect 15853 28033 15887 28067
rect 17049 28033 17083 28067
rect 17141 28033 17175 28067
rect 19533 28033 19567 28067
rect 19993 28033 20027 28067
rect 21005 28033 21039 28067
rect 22201 28033 22235 28067
rect 22569 28033 22603 28067
rect 22836 28033 22870 28067
rect 24409 28033 24443 28067
rect 24593 28033 24627 28067
rect 24685 28033 24719 28067
rect 24961 28033 24995 28067
rect 25237 28033 25271 28067
rect 25421 28033 25455 28067
rect 25513 28033 25547 28067
rect 25789 28033 25823 28067
rect 26065 28033 26099 28067
rect 27997 28033 28031 28067
rect 30665 28033 30699 28067
rect 31585 28033 31619 28067
rect 31769 28033 31803 28067
rect 34345 28033 34379 28067
rect 34529 28033 34563 28067
rect 37289 28033 37323 28067
rect 37437 28033 37471 28067
rect 37754 28033 37788 28067
rect 38025 28033 38059 28067
rect 1869 27965 1903 27999
rect 3617 27965 3651 27999
rect 6929 27965 6963 27999
rect 7113 27965 7147 27999
rect 7481 27965 7515 27999
rect 7849 27965 7883 27999
rect 9321 27965 9355 27999
rect 12357 27965 12391 27999
rect 14013 27965 14047 27999
rect 15485 27965 15519 27999
rect 17233 27965 17267 27999
rect 18061 27965 18095 27999
rect 18153 27965 18187 27999
rect 20269 27965 20303 27999
rect 20913 27965 20947 27999
rect 21097 27965 21131 27999
rect 21189 27965 21223 27999
rect 24777 27965 24811 27999
rect 25605 27965 25639 27999
rect 26617 27965 26651 27999
rect 26985 27965 27019 27999
rect 29929 27965 29963 27999
rect 30941 27965 30975 27999
rect 31493 27965 31527 27999
rect 32229 27965 32263 27999
rect 33977 27965 34011 27999
rect 34253 27965 34287 27999
rect 4721 27897 4755 27931
rect 25145 27897 25179 27931
rect 30757 27897 30791 27931
rect 3709 27829 3743 27863
rect 5365 27829 5399 27863
rect 5457 27829 5491 27863
rect 5641 27829 5675 27863
rect 6561 27829 6595 27863
rect 7021 27829 7055 27863
rect 13829 27829 13863 27863
rect 16681 27829 16715 27863
rect 19901 27829 19935 27863
rect 20085 27829 20119 27863
rect 21833 27829 21867 27863
rect 27629 27829 27663 27863
rect 30849 27829 30883 27863
rect 31953 27829 31987 27863
rect 34529 27829 34563 27863
rect 38209 27829 38243 27863
rect 3433 27625 3467 27659
rect 3617 27625 3651 27659
rect 3985 27625 4019 27659
rect 7389 27625 7423 27659
rect 11332 27625 11366 27659
rect 14381 27625 14415 27659
rect 16969 27625 17003 27659
rect 20085 27625 20119 27659
rect 27371 27625 27405 27659
rect 28181 27625 28215 27659
rect 28825 27625 28859 27659
rect 31309 27625 31343 27659
rect 31769 27625 31803 27659
rect 33241 27625 33275 27659
rect 38393 27625 38427 27659
rect 4261 27557 4295 27591
rect 13001 27557 13035 27591
rect 15117 27557 15151 27591
rect 20453 27557 20487 27591
rect 25881 27557 25915 27591
rect 28549 27557 28583 27591
rect 28641 27557 28675 27591
rect 32137 27557 32171 27591
rect 32873 27557 32907 27591
rect 37105 27557 37139 27591
rect 3893 27489 3927 27523
rect 13553 27489 13587 27523
rect 17233 27489 17267 27523
rect 19717 27489 19751 27523
rect 21557 27489 21591 27523
rect 24225 27489 24259 27523
rect 25329 27489 25363 27523
rect 25789 27489 25823 27523
rect 27629 27489 27663 27523
rect 30849 27489 30883 27523
rect 31125 27489 31159 27523
rect 31861 27489 31895 27523
rect 32781 27489 32815 27523
rect 1409 27421 1443 27455
rect 3801 27421 3835 27455
rect 4077 27421 4111 27455
rect 7297 27421 7331 27455
rect 7481 27421 7515 27455
rect 11069 27421 11103 27455
rect 14289 27421 14323 27455
rect 14657 27421 14691 27455
rect 15209 27421 15243 27455
rect 17498 27421 17532 27455
rect 17602 27421 17636 27455
rect 18061 27421 18095 27455
rect 18245 27431 18279 27465
rect 18429 27421 18463 27455
rect 19349 27421 19383 27455
rect 19533 27421 19567 27455
rect 19625 27421 19659 27455
rect 19809 27421 19843 27455
rect 20085 27421 20119 27455
rect 20269 27421 20303 27455
rect 21281 27421 21315 27455
rect 21465 27421 21499 27455
rect 21649 27421 21683 27455
rect 21833 27421 21867 27455
rect 22109 27421 22143 27455
rect 23949 27421 23983 27455
rect 24133 27421 24167 27455
rect 24777 27421 24811 27455
rect 25053 27421 25087 27455
rect 25237 27421 25271 27455
rect 25421 27421 25455 27455
rect 25605 27421 25639 27455
rect 30757 27421 30791 27455
rect 31217 27421 31251 27455
rect 31493 27421 31527 27455
rect 31769 27421 31803 27455
rect 33057 27421 33091 27455
rect 35173 27421 35207 27455
rect 35357 27421 35391 27455
rect 37013 27421 37047 27455
rect 37532 27421 37566 27455
rect 37749 27421 37783 27455
rect 37933 27421 37967 27455
rect 38025 27421 38059 27455
rect 38117 27421 38151 27455
rect 1685 27353 1719 27387
rect 3249 27353 3283 27387
rect 3449 27353 3483 27387
rect 4353 27353 4387 27387
rect 5181 27353 5215 27387
rect 18705 27353 18739 27387
rect 18889 27353 18923 27387
rect 20821 27353 20855 27387
rect 20913 27353 20947 27387
rect 21189 27353 21223 27387
rect 22017 27353 22051 27387
rect 22354 27353 22388 27387
rect 24409 27353 24443 27387
rect 24593 27353 24627 27387
rect 29009 27353 29043 27387
rect 31677 27353 31711 27387
rect 3157 27285 3191 27319
rect 5457 27285 5491 27319
rect 12817 27285 12851 27319
rect 13369 27285 13403 27319
rect 13461 27285 13495 27319
rect 14841 27285 14875 27319
rect 17877 27285 17911 27319
rect 18153 27285 18187 27319
rect 18521 27285 18555 27319
rect 19073 27285 19107 27319
rect 19993 27285 20027 27319
rect 20637 27285 20671 27319
rect 21005 27285 21039 27319
rect 23489 27285 23523 27319
rect 27997 27285 28031 27319
rect 28181 27285 28215 27319
rect 28809 27285 28843 27319
rect 35265 27285 35299 27319
rect 37473 27285 37507 27319
rect 37657 27285 37691 27319
rect 3525 27081 3559 27115
rect 13001 27081 13035 27115
rect 21373 27081 21407 27115
rect 22661 27081 22695 27115
rect 25973 27081 26007 27115
rect 33701 27081 33735 27115
rect 37013 27081 37047 27115
rect 38393 27081 38427 27115
rect 12909 27013 12943 27047
rect 15209 27013 15243 27047
rect 15577 27013 15611 27047
rect 16221 27013 16255 27047
rect 18889 27013 18923 27047
rect 19257 27013 19291 27047
rect 21925 27013 21959 27047
rect 27721 27013 27755 27047
rect 28917 27013 28951 27047
rect 30849 27013 30883 27047
rect 38025 27013 38059 27047
rect 2329 26945 2363 26979
rect 2789 26945 2823 26979
rect 3341 26945 3375 26979
rect 5365 26945 5399 26979
rect 6009 26945 6043 26979
rect 6193 26945 6227 26979
rect 13829 26945 13863 26979
rect 14013 26945 14047 26979
rect 14105 26945 14139 26979
rect 14289 26945 14323 26979
rect 15117 26945 15151 26979
rect 15301 26945 15335 26979
rect 15485 26945 15519 26979
rect 15669 26945 15703 26979
rect 15945 26945 15979 26979
rect 19073 26945 19107 26979
rect 19625 26945 19659 26979
rect 19809 26945 19843 26979
rect 20085 26945 20119 26979
rect 21465 26945 21499 26979
rect 21833 26945 21867 26979
rect 22017 26945 22051 26979
rect 23305 26945 23339 26979
rect 24225 26945 24259 26979
rect 26065 26945 26099 26979
rect 26249 26945 26283 26979
rect 26433 26945 26467 26979
rect 26617 26945 26651 26979
rect 27537 26945 27571 26979
rect 28641 26945 28675 26979
rect 31033 26945 31067 26979
rect 32229 26945 32263 26979
rect 32413 26945 32447 26979
rect 32689 26945 32723 26979
rect 35449 26945 35483 26979
rect 35725 26945 35759 26979
rect 36461 26945 36495 26979
rect 36553 26945 36587 26979
rect 36737 26945 36771 26979
rect 36829 26945 36863 26979
rect 37657 26945 37691 26979
rect 37933 26945 37967 26979
rect 38117 26945 38151 26979
rect 38209 26945 38243 26979
rect 1961 26877 1995 26911
rect 2421 26877 2455 26911
rect 4997 26877 5031 26911
rect 5273 26877 5307 26911
rect 7573 26877 7607 26911
rect 7849 26877 7883 26911
rect 9413 26877 9447 26911
rect 9689 26877 9723 26911
rect 11161 26877 11195 26911
rect 12081 26877 12115 26911
rect 15761 26877 15795 26911
rect 16313 26877 16347 26911
rect 23581 26877 23615 26911
rect 24133 26877 24167 26911
rect 24501 26877 24535 26911
rect 26341 26877 26375 26911
rect 28273 26877 28307 26911
rect 35173 26877 35207 26911
rect 35633 26877 35667 26911
rect 36093 26877 36127 26911
rect 37381 26877 37415 26911
rect 37841 26877 37875 26911
rect 26801 26809 26835 26843
rect 6009 26741 6043 26775
rect 9321 26741 9355 26775
rect 11529 26741 11563 26775
rect 13921 26741 13955 26775
rect 14289 26741 14323 26775
rect 19441 26741 19475 26775
rect 19993 26741 20027 26775
rect 26985 26741 27019 26775
rect 30389 26741 30423 26775
rect 31125 26741 31159 26775
rect 32873 26741 32907 26775
rect 37473 26741 37507 26775
rect 3065 26537 3099 26571
rect 3985 26537 4019 26571
rect 8309 26537 8343 26571
rect 9873 26537 9907 26571
rect 13185 26537 13219 26571
rect 19441 26537 19475 26571
rect 20361 26537 20395 26571
rect 24409 26537 24443 26571
rect 25513 26537 25547 26571
rect 28089 26537 28123 26571
rect 30205 26537 30239 26571
rect 35265 26537 35299 26571
rect 35449 26537 35483 26571
rect 36553 26537 36587 26571
rect 37473 26537 37507 26571
rect 17877 26469 17911 26503
rect 20729 26469 20763 26503
rect 2881 26401 2915 26435
rect 6469 26401 6503 26435
rect 8217 26401 8251 26435
rect 10241 26401 10275 26435
rect 14105 26401 14139 26435
rect 14565 26401 14599 26435
rect 15853 26401 15887 26435
rect 16221 26401 16255 26435
rect 16338 26401 16372 26435
rect 17693 26401 17727 26435
rect 19533 26401 19567 26435
rect 20269 26401 20303 26435
rect 20453 26401 20487 26435
rect 27261 26401 27295 26435
rect 27905 26401 27939 26435
rect 29929 26401 29963 26435
rect 30573 26401 30607 26435
rect 37657 26401 37691 26435
rect 2789 26333 2823 26367
rect 2973 26333 3007 26367
rect 3249 26333 3283 26367
rect 3433 26333 3467 26367
rect 3801 26333 3835 26367
rect 3985 26333 4019 26367
rect 4629 26333 4663 26367
rect 8493 26333 8527 26367
rect 8677 26333 8711 26367
rect 8769 26333 8803 26367
rect 9137 26333 9171 26367
rect 9689 26333 9723 26367
rect 9873 26333 9907 26367
rect 10057 26333 10091 26367
rect 13093 26333 13127 26367
rect 13277 26333 13311 26367
rect 13553 26333 13587 26367
rect 13646 26333 13680 26367
rect 14473 26333 14507 26367
rect 15301 26333 15335 26367
rect 15485 26333 15519 26367
rect 17325 26333 17359 26367
rect 17479 26333 17513 26367
rect 17785 26333 17819 26367
rect 17969 26333 18003 26367
rect 18153 26333 18187 26367
rect 18337 26333 18371 26367
rect 18613 26333 18647 26367
rect 18797 26333 18831 26367
rect 19441 26333 19475 26367
rect 19901 26333 19935 26367
rect 20361 26333 20395 26367
rect 20821 26333 20855 26367
rect 24593 26333 24627 26367
rect 24777 26333 24811 26367
rect 24869 26333 24903 26367
rect 24961 26333 24995 26367
rect 25145 26333 25179 26367
rect 28273 26333 28307 26367
rect 28457 26333 28491 26367
rect 29101 26333 29135 26367
rect 29285 26333 29319 26367
rect 29561 26333 29595 26367
rect 29745 26333 29779 26367
rect 31033 26333 31067 26367
rect 31217 26333 31251 26367
rect 35081 26333 35115 26367
rect 35357 26333 35391 26367
rect 35541 26333 35575 26367
rect 35909 26333 35943 26367
rect 36093 26333 36127 26367
rect 36185 26333 36219 26367
rect 36277 26333 36311 26367
rect 37749 26333 37783 26367
rect 4905 26265 4939 26299
rect 6745 26265 6779 26299
rect 10517 26265 10551 26299
rect 14197 26265 14231 26299
rect 20085 26265 20119 26299
rect 23857 26265 23891 26299
rect 24041 26265 24075 26299
rect 24225 26265 24259 26299
rect 26985 26265 27019 26299
rect 27353 26265 27387 26299
rect 28549 26265 28583 26299
rect 30113 26265 30147 26299
rect 30481 26265 30515 26299
rect 34897 26265 34931 26299
rect 38117 26265 38151 26299
rect 6377 26197 6411 26231
rect 11989 26197 12023 26231
rect 13921 26197 13955 26231
rect 14749 26197 14783 26231
rect 15301 26197 15335 26231
rect 16129 26197 16163 26231
rect 16497 26197 16531 26231
rect 18521 26197 18555 26231
rect 18705 26197 18739 26231
rect 19809 26197 19843 26231
rect 20913 26197 20947 26231
rect 29193 26197 29227 26231
rect 31033 26197 31067 26231
rect 8769 25993 8803 26027
rect 9597 25993 9631 26027
rect 13277 25993 13311 26027
rect 13645 25993 13679 26027
rect 15945 25993 15979 26027
rect 24225 25993 24259 26027
rect 25421 25993 25455 26027
rect 29837 25993 29871 26027
rect 31493 25993 31527 26027
rect 31861 25993 31895 26027
rect 33517 25993 33551 26027
rect 35725 25993 35759 26027
rect 36277 25993 36311 26027
rect 5641 25925 5675 25959
rect 6009 25925 6043 25959
rect 6377 25925 6411 25959
rect 9105 25925 9139 25959
rect 9321 25925 9355 25959
rect 9781 25925 9815 25959
rect 10669 25925 10703 25959
rect 10885 25925 10919 25959
rect 15209 25925 15243 25959
rect 20177 25925 20211 25959
rect 20913 25925 20947 25959
rect 21281 25925 21315 25959
rect 21833 25925 21867 25959
rect 25053 25925 25087 25959
rect 28365 25925 28399 25959
rect 32413 25925 32447 25959
rect 37657 25925 37691 25959
rect 3249 25857 3283 25891
rect 3433 25857 3467 25891
rect 5825 25857 5859 25891
rect 6101 25857 6135 25891
rect 7205 25857 7239 25891
rect 7389 25857 7423 25891
rect 7665 25857 7699 25891
rect 8677 25857 8711 25891
rect 8861 25857 8895 25891
rect 9505 25857 9539 25891
rect 10057 25857 10091 25891
rect 11529 25857 11563 25891
rect 12081 25857 12115 25891
rect 12541 25857 12575 25891
rect 12725 25857 12759 25891
rect 12817 25857 12851 25891
rect 13961 25857 13995 25891
rect 14105 25857 14139 25891
rect 14197 25857 14231 25891
rect 14381 25857 14415 25891
rect 14933 25857 14967 25891
rect 15301 25857 15335 25891
rect 15485 25857 15519 25891
rect 15761 25857 15795 25891
rect 16221 25857 16255 25891
rect 17601 25857 17635 25891
rect 17785 25857 17819 25891
rect 18245 25857 18279 25891
rect 18429 25857 18463 25891
rect 18521 25857 18555 25891
rect 18705 25857 18739 25891
rect 18889 25857 18923 25891
rect 19073 25857 19107 25891
rect 19349 25857 19383 25891
rect 19533 25857 19567 25891
rect 19625 25857 19659 25891
rect 19717 25857 19751 25891
rect 20545 25857 20579 25891
rect 20637 25857 20671 25891
rect 21097 25857 21131 25891
rect 21373 25857 21407 25891
rect 21557 25857 21591 25891
rect 22293 25857 22327 25891
rect 22845 25857 22879 25891
rect 23112 25857 23146 25891
rect 24869 25857 24903 25891
rect 25237 25857 25271 25891
rect 27813 25857 27847 25891
rect 27905 25857 27939 25891
rect 30021 25857 30055 25891
rect 32137 25857 32171 25891
rect 32321 25857 32355 25891
rect 32505 25857 32539 25891
rect 32781 25857 32815 25891
rect 32965 25857 32999 25891
rect 33333 25857 33367 25891
rect 33609 25857 33643 25891
rect 33793 25857 33827 25891
rect 34161 25857 34195 25891
rect 34345 25857 34379 25891
rect 35081 25857 35115 25891
rect 35173 25857 35207 25891
rect 35357 25857 35391 25891
rect 35449 25857 35483 25891
rect 35541 25857 35575 25891
rect 35817 25857 35851 25891
rect 35909 25857 35943 25891
rect 36093 25857 36127 25891
rect 37841 25857 37875 25891
rect 5733 25789 5767 25823
rect 6929 25789 6963 25823
rect 7481 25789 7515 25823
rect 7849 25789 7883 25823
rect 8493 25789 8527 25823
rect 10149 25789 10183 25823
rect 10425 25789 10459 25823
rect 13093 25789 13127 25823
rect 13185 25789 13219 25823
rect 15025 25789 15059 25823
rect 15209 25789 15243 25823
rect 16129 25789 16163 25823
rect 18797 25789 18831 25823
rect 20269 25789 20303 25823
rect 22201 25789 22235 25823
rect 27629 25789 27663 25823
rect 28089 25789 28123 25823
rect 33057 25789 33091 25823
rect 33149 25789 33183 25823
rect 34253 25789 34287 25823
rect 37473 25789 37507 25823
rect 7941 25721 7975 25755
rect 9781 25721 9815 25755
rect 20821 25721 20855 25755
rect 32689 25721 32723 25755
rect 33701 25721 33735 25755
rect 3433 25653 3467 25687
rect 7205 25653 7239 25687
rect 8953 25653 8987 25687
rect 9137 25653 9171 25687
rect 10517 25653 10551 25687
rect 10701 25653 10735 25687
rect 12357 25653 12391 25687
rect 13829 25653 13863 25687
rect 17601 25653 17635 25687
rect 17969 25653 18003 25687
rect 18429 25653 18463 25687
rect 19257 25653 19291 25687
rect 19993 25653 20027 25687
rect 21373 25653 21407 25687
rect 22109 25653 22143 25687
rect 22477 25653 22511 25687
rect 24317 25653 24351 25687
rect 27721 25653 27755 25687
rect 3249 25449 3283 25483
rect 3433 25449 3467 25483
rect 6101 25449 6135 25483
rect 7113 25449 7147 25483
rect 8309 25449 8343 25483
rect 12817 25449 12851 25483
rect 13645 25449 13679 25483
rect 15209 25449 15243 25483
rect 15577 25449 15611 25483
rect 15669 25449 15703 25483
rect 18245 25449 18279 25483
rect 20085 25449 20119 25483
rect 20545 25449 20579 25483
rect 21925 25449 21959 25483
rect 23305 25449 23339 25483
rect 24961 25449 24995 25483
rect 25881 25449 25915 25483
rect 31125 25449 31159 25483
rect 32505 25449 32539 25483
rect 33241 25449 33275 25483
rect 35081 25449 35115 25483
rect 36737 25449 36771 25483
rect 37013 25449 37047 25483
rect 37749 25449 37783 25483
rect 37841 25449 37875 25483
rect 9873 25381 9907 25415
rect 16037 25381 16071 25415
rect 28641 25381 28675 25415
rect 1409 25313 1443 25347
rect 3801 25313 3835 25347
rect 4077 25313 4111 25347
rect 13461 25313 13495 25347
rect 18337 25313 18371 25347
rect 20269 25313 20303 25347
rect 21005 25313 21039 25347
rect 26157 25313 26191 25347
rect 30481 25313 30515 25347
rect 31493 25313 31527 25347
rect 31585 25313 31619 25347
rect 37289 25313 37323 25347
rect 5641 25245 5675 25279
rect 5825 25245 5859 25279
rect 6929 25245 6963 25279
rect 7113 25245 7147 25279
rect 7849 25245 7883 25279
rect 7941 25245 7975 25279
rect 8309 25245 8343 25279
rect 10241 25245 10275 25279
rect 10425 25245 10459 25279
rect 12357 25245 12391 25279
rect 12541 25245 12575 25279
rect 13001 25245 13035 25279
rect 13303 25245 13337 25279
rect 13737 25245 13771 25279
rect 15117 25245 15151 25279
rect 15393 25245 15427 25279
rect 15669 25245 15703 25279
rect 15853 25245 15887 25279
rect 15945 25245 15979 25279
rect 16313 25245 16347 25279
rect 18061 25245 18095 25279
rect 18153 25245 18187 25279
rect 18429 25245 18463 25279
rect 18613 25245 18647 25279
rect 19901 25245 19935 25279
rect 20361 25245 20395 25279
rect 20913 25245 20947 25279
rect 21097 25245 21131 25279
rect 21189 25245 21223 25279
rect 21281 25245 21315 25279
rect 22017 25245 22051 25279
rect 22201 25245 22235 25279
rect 22661 25245 22695 25279
rect 22845 25245 22879 25279
rect 22937 25245 22971 25279
rect 23029 25245 23063 25279
rect 25513 25245 25547 25279
rect 27997 25245 28031 25279
rect 28181 25245 28215 25279
rect 28273 25245 28307 25279
rect 28365 25245 28399 25279
rect 30941 25245 30975 25279
rect 31217 25245 31251 25279
rect 31401 25245 31435 25279
rect 31769 25245 31803 25279
rect 32229 25245 32263 25279
rect 32321 25245 32355 25279
rect 32689 25245 32723 25279
rect 32781 25245 32815 25279
rect 33425 25245 33459 25279
rect 33609 25245 33643 25279
rect 36553 25245 36587 25279
rect 36737 25245 36771 25279
rect 37381 25245 37415 25279
rect 37565 25245 37599 25279
rect 37841 25245 37875 25279
rect 37933 25245 37967 25279
rect 1685 25177 1719 25211
rect 3401 25177 3435 25211
rect 3617 25177 3651 25211
rect 6085 25177 6119 25211
rect 6285 25177 6319 25211
rect 10057 25177 10091 25211
rect 13093 25177 13127 25211
rect 13185 25177 13219 25211
rect 16037 25177 16071 25211
rect 16221 25177 16255 25211
rect 21557 25177 21591 25211
rect 22109 25177 22143 25211
rect 25145 25177 25179 25211
rect 26433 25177 26467 25211
rect 30619 25177 30653 25211
rect 30757 25177 30791 25211
rect 30849 25177 30883 25211
rect 32045 25177 32079 25211
rect 34713 25177 34747 25211
rect 34897 25177 34931 25211
rect 37197 25177 37231 25211
rect 38117 25177 38151 25211
rect 3157 25109 3191 25143
rect 5549 25109 5583 25143
rect 5733 25109 5767 25143
rect 5917 25109 5951 25143
rect 8493 25109 8527 25143
rect 10333 25109 10367 25143
rect 11069 25109 11103 25143
rect 12633 25109 12667 25143
rect 18613 25109 18647 25143
rect 21465 25109 21499 25143
rect 21643 25109 21677 25143
rect 24777 25109 24811 25143
rect 24945 25109 24979 25143
rect 25881 25109 25915 25143
rect 26065 25109 26099 25143
rect 27905 25109 27939 25143
rect 29837 25109 29871 25143
rect 31953 25109 31987 25143
rect 36829 25109 36863 25143
rect 36997 25109 37031 25143
rect 6193 24905 6227 24939
rect 13737 24905 13771 24939
rect 15301 24905 15335 24939
rect 16221 24905 16255 24939
rect 18521 24905 18555 24939
rect 19165 24905 19199 24939
rect 21557 24905 21591 24939
rect 22845 24905 22879 24939
rect 30941 24905 30975 24939
rect 31309 24905 31343 24939
rect 32597 24905 32631 24939
rect 32689 24905 32723 24939
rect 33793 24905 33827 24939
rect 34529 24905 34563 24939
rect 35633 24905 35667 24939
rect 36001 24905 36035 24939
rect 9045 24837 9079 24871
rect 14565 24837 14599 24871
rect 18797 24837 18831 24871
rect 24777 24837 24811 24871
rect 31585 24837 31619 24871
rect 33609 24837 33643 24871
rect 34161 24837 34195 24871
rect 34361 24837 34395 24871
rect 1685 24769 1719 24803
rect 2145 24769 2179 24803
rect 2605 24769 2639 24803
rect 4169 24769 4203 24803
rect 6561 24769 6595 24803
rect 6929 24769 6963 24803
rect 7205 24769 7239 24803
rect 7481 24769 7515 24803
rect 8217 24769 8251 24803
rect 8493 24769 8527 24803
rect 8769 24769 8803 24803
rect 8861 24769 8895 24803
rect 9137 24769 9171 24803
rect 9597 24769 9631 24803
rect 10241 24769 10275 24803
rect 10517 24769 10551 24803
rect 10609 24769 10643 24803
rect 10793 24769 10827 24803
rect 11069 24769 11103 24803
rect 11529 24769 11563 24803
rect 12081 24769 12115 24803
rect 13001 24769 13035 24803
rect 13185 24769 13219 24803
rect 13369 24769 13403 24803
rect 13921 24769 13955 24803
rect 14013 24769 14047 24803
rect 14197 24769 14231 24803
rect 14289 24769 14323 24803
rect 14381 24769 14415 24803
rect 15209 24769 15243 24803
rect 15485 24769 15519 24803
rect 15577 24769 15611 24803
rect 15761 24769 15795 24803
rect 15853 24769 15887 24803
rect 16129 24769 16163 24803
rect 16313 24769 16347 24803
rect 18153 24769 18187 24803
rect 18337 24769 18371 24803
rect 18613 24769 18647 24803
rect 18889 24769 18923 24803
rect 18981 24769 19015 24803
rect 21189 24769 21223 24803
rect 21373 24769 21407 24803
rect 21833 24769 21867 24803
rect 22109 24769 22143 24803
rect 22385 24769 22419 24803
rect 22661 24769 22695 24803
rect 23296 24769 23330 24803
rect 24501 24769 24535 24803
rect 27169 24769 27203 24803
rect 27445 24769 27479 24803
rect 30573 24769 30607 24803
rect 30757 24769 30791 24803
rect 30849 24769 30883 24803
rect 31125 24769 31159 24803
rect 31401 24769 31435 24803
rect 31769 24769 31803 24803
rect 32137 24769 32171 24803
rect 32229 24769 32263 24803
rect 32413 24769 32447 24803
rect 32689 24769 32723 24803
rect 32781 24769 32815 24803
rect 32965 24769 32999 24803
rect 33149 24769 33183 24803
rect 33241 24769 33275 24803
rect 33425 24769 33459 24803
rect 33701 24769 33735 24803
rect 33885 24769 33919 24803
rect 33977 24769 34011 24803
rect 34621 24769 34655 24803
rect 34713 24769 34747 24803
rect 34897 24769 34931 24803
rect 35265 24769 35299 24803
rect 35725 24769 35759 24803
rect 36737 24769 36771 24803
rect 36829 24769 36863 24803
rect 37013 24769 37047 24803
rect 1777 24701 1811 24735
rect 2053 24701 2087 24735
rect 2697 24701 2731 24735
rect 3249 24701 3283 24735
rect 4445 24701 4479 24735
rect 4721 24701 4755 24735
rect 6469 24701 6503 24735
rect 7297 24701 7331 24735
rect 9505 24701 9539 24735
rect 10977 24701 11011 24735
rect 15117 24701 15151 24735
rect 22017 24701 22051 24735
rect 22477 24701 22511 24735
rect 23029 24701 23063 24735
rect 26985 24701 27019 24735
rect 27261 24701 27295 24735
rect 27353 24701 27387 24735
rect 29101 24701 29135 24735
rect 29561 24701 29595 24735
rect 35357 24701 35391 24735
rect 36001 24701 36035 24735
rect 1501 24633 1535 24667
rect 2421 24633 2455 24667
rect 7113 24633 7147 24667
rect 29193 24633 29227 24667
rect 30665 24633 30699 24667
rect 34897 24633 34931 24667
rect 35817 24633 35851 24667
rect 37013 24633 37047 24667
rect 3525 24565 3559 24599
rect 6837 24565 6871 24599
rect 7205 24565 7239 24599
rect 7665 24565 7699 24599
rect 9229 24565 9263 24599
rect 9781 24565 9815 24599
rect 10793 24565 10827 24599
rect 14749 24565 14783 24599
rect 21281 24565 21315 24599
rect 21833 24565 21867 24599
rect 22293 24565 22327 24599
rect 22385 24565 22419 24599
rect 24409 24565 24443 24599
rect 26249 24565 26283 24599
rect 34345 24565 34379 24599
rect 35449 24565 35483 24599
rect 3249 24361 3283 24395
rect 4537 24361 4571 24395
rect 5641 24361 5675 24395
rect 7389 24361 7423 24395
rect 7849 24361 7883 24395
rect 8217 24361 8251 24395
rect 9597 24361 9631 24395
rect 11989 24361 12023 24395
rect 13277 24361 13311 24395
rect 14105 24361 14139 24395
rect 14933 24361 14967 24395
rect 18061 24361 18095 24395
rect 19441 24361 19475 24395
rect 19901 24361 19935 24395
rect 21373 24361 21407 24395
rect 21833 24361 21867 24395
rect 23489 24361 23523 24395
rect 25145 24361 25179 24395
rect 25697 24361 25731 24395
rect 26433 24361 26467 24395
rect 27721 24361 27755 24395
rect 28641 24361 28675 24395
rect 29561 24361 29595 24395
rect 31861 24361 31895 24395
rect 32689 24361 32723 24395
rect 33885 24361 33919 24395
rect 35541 24361 35575 24395
rect 37657 24361 37691 24395
rect 4997 24293 5031 24327
rect 9413 24293 9447 24327
rect 13185 24293 13219 24327
rect 15669 24293 15703 24327
rect 16957 24293 16991 24327
rect 18337 24293 18371 24327
rect 19717 24293 19751 24327
rect 27169 24293 27203 24327
rect 30205 24293 30239 24327
rect 36461 24293 36495 24327
rect 4721 24225 4755 24259
rect 6561 24225 6595 24259
rect 7297 24225 7331 24259
rect 7481 24225 7515 24259
rect 8217 24225 8251 24259
rect 9781 24225 9815 24259
rect 10241 24225 10275 24259
rect 10517 24225 10551 24259
rect 12909 24225 12943 24259
rect 13737 24225 13771 24259
rect 14657 24225 14691 24259
rect 15117 24225 15151 24259
rect 15577 24225 15611 24259
rect 18521 24225 18555 24259
rect 19809 24225 19843 24259
rect 21741 24225 21775 24259
rect 21925 24225 21959 24259
rect 25053 24225 25087 24259
rect 27077 24225 27111 24259
rect 28825 24225 28859 24259
rect 29285 24225 29319 24259
rect 31401 24225 31435 24259
rect 35909 24225 35943 24259
rect 2973 24157 3007 24191
rect 3249 24157 3283 24191
rect 3341 24157 3375 24191
rect 3525 24157 3559 24191
rect 3801 24157 3835 24191
rect 4353 24157 4387 24191
rect 4813 24157 4847 24191
rect 5917 24157 5951 24191
rect 6837 24157 6871 24191
rect 6929 24157 6963 24191
rect 7389 24157 7423 24191
rect 7665 24157 7699 24191
rect 8125 24157 8159 24191
rect 9597 24157 9631 24191
rect 12817 24157 12851 24191
rect 13645 24157 13679 24191
rect 15209 24157 15243 24191
rect 15945 24157 15979 24191
rect 16129 24157 16163 24191
rect 16221 24157 16255 24191
rect 16405 24157 16439 24191
rect 16681 24157 16715 24191
rect 16773 24157 16807 24191
rect 17877 24157 17911 24191
rect 18061 24157 18095 24191
rect 18245 24157 18279 24191
rect 18613 24157 18647 24191
rect 18791 24157 18825 24191
rect 18889 24159 18923 24193
rect 19073 24157 19107 24191
rect 19993 24157 20027 24191
rect 20177 24157 20211 24191
rect 21373 24157 21407 24191
rect 21557 24157 21591 24191
rect 21649 24157 21683 24191
rect 22845 24157 22879 24191
rect 23029 24157 23063 24191
rect 23121 24157 23155 24191
rect 23213 24157 23247 24191
rect 24409 24157 24443 24191
rect 25329 24157 25363 24191
rect 25605 24157 25639 24191
rect 25697 24157 25731 24191
rect 25789 24157 25823 24191
rect 26801 24157 26835 24191
rect 27540 24157 27574 24191
rect 28365 24157 28399 24191
rect 28641 24157 28675 24191
rect 28917 24157 28951 24191
rect 29745 24157 29779 24191
rect 30205 24157 30239 24191
rect 30389 24157 30423 24191
rect 31033 24157 31067 24191
rect 31493 24157 31527 24191
rect 31677 24157 31711 24191
rect 31769 24157 31803 24191
rect 31953 24157 31987 24191
rect 32597 24157 32631 24191
rect 32781 24157 32815 24191
rect 33793 24157 33827 24191
rect 33977 24157 34011 24191
rect 35817 24157 35851 24191
rect 36082 24157 36116 24191
rect 36247 24157 36281 24191
rect 3065 24089 3099 24123
rect 4537 24089 4571 24123
rect 5641 24089 5675 24123
rect 6009 24089 6043 24123
rect 7021 24089 7055 24123
rect 7113 24089 7147 24123
rect 10057 24089 10091 24123
rect 14565 24089 14599 24123
rect 15669 24089 15703 24123
rect 16957 24089 16991 24123
rect 18521 24089 18555 24123
rect 25513 24089 25547 24123
rect 25973 24089 26007 24123
rect 26985 24089 27019 24123
rect 28457 24089 28491 24123
rect 30113 24089 30147 24123
rect 31217 24089 31251 24123
rect 37289 24089 37323 24123
rect 37473 24089 37507 24123
rect 3433 24021 3467 24055
rect 5825 24021 5859 24055
rect 8493 24021 8527 24055
rect 14473 24021 14507 24055
rect 15853 24021 15887 24055
rect 16589 24021 16623 24055
rect 18705 24021 18739 24055
rect 18981 24021 19015 24055
rect 26617 24021 26651 24055
rect 26709 24021 26743 24055
rect 27537 24021 27571 24055
rect 29837 24021 29871 24055
rect 29929 24021 29963 24055
rect 31677 24021 31711 24055
rect 3249 23817 3283 23851
rect 3969 23817 4003 23851
rect 8033 23817 8067 23851
rect 8493 23817 8527 23851
rect 8585 23817 8619 23851
rect 9229 23817 9263 23851
rect 14473 23817 14507 23851
rect 14841 23817 14875 23851
rect 18521 23817 18555 23851
rect 22201 23817 22235 23851
rect 29009 23817 29043 23851
rect 30573 23817 30607 23851
rect 31677 23817 31711 23851
rect 32873 23817 32907 23851
rect 33149 23817 33183 23851
rect 33977 23817 34011 23851
rect 34529 23817 34563 23851
rect 35265 23817 35299 23851
rect 36369 23817 36403 23851
rect 37933 23817 37967 23851
rect 4169 23749 4203 23783
rect 9873 23749 9907 23783
rect 10609 23749 10643 23783
rect 11253 23749 11287 23783
rect 13461 23749 13495 23783
rect 14657 23749 14691 23783
rect 15025 23749 15059 23783
rect 16773 23749 16807 23783
rect 17601 23749 17635 23783
rect 17969 23749 18003 23783
rect 18153 23749 18187 23783
rect 19441 23749 19475 23783
rect 26985 23749 27019 23783
rect 28273 23749 28307 23783
rect 30389 23749 30423 23783
rect 32689 23749 32723 23783
rect 34161 23749 34195 23783
rect 36645 23749 36679 23783
rect 37013 23749 37047 23783
rect 3433 23681 3467 23715
rect 7941 23681 7975 23715
rect 8376 23681 8410 23715
rect 8953 23681 8987 23715
rect 9137 23681 9171 23715
rect 9229 23681 9263 23715
rect 9597 23681 9631 23715
rect 9781 23681 9815 23715
rect 10885 23681 10919 23715
rect 11069 23681 11103 23715
rect 14381 23681 14415 23715
rect 14749 23681 14783 23715
rect 16687 23681 16721 23715
rect 16865 23681 16899 23715
rect 17325 23681 17359 23715
rect 17509 23681 17543 23715
rect 17785 23681 17819 23715
rect 18061 23681 18095 23715
rect 18239 23681 18273 23715
rect 19067 23671 19101 23705
rect 19257 23681 19291 23715
rect 19533 23681 19567 23715
rect 19625 23681 19659 23715
rect 19993 23681 20027 23715
rect 20269 23681 20303 23715
rect 20361 23681 20395 23715
rect 21189 23681 21223 23715
rect 21373 23681 21407 23715
rect 21833 23681 21867 23715
rect 22017 23681 22051 23715
rect 24409 23681 24443 23715
rect 25053 23681 25087 23715
rect 25421 23681 25455 23715
rect 25513 23681 25547 23715
rect 26709 23681 26743 23715
rect 27997 23681 28031 23715
rect 28181 23681 28215 23715
rect 29193 23681 29227 23715
rect 29285 23681 29319 23715
rect 29377 23681 29411 23715
rect 29469 23681 29503 23715
rect 30205 23681 30239 23715
rect 30481 23681 30515 23715
rect 30665 23681 30699 23715
rect 31585 23681 31619 23715
rect 31769 23681 31803 23715
rect 32505 23681 32539 23715
rect 32965 23681 32999 23715
rect 33149 23681 33183 23715
rect 34345 23681 34379 23715
rect 34437 23681 34471 23715
rect 34621 23681 34655 23715
rect 34897 23681 34931 23715
rect 35081 23681 35115 23715
rect 36277 23681 36311 23715
rect 36461 23681 36495 23715
rect 37105 23681 37139 23715
rect 37289 23681 37323 23715
rect 37473 23681 37507 23715
rect 37565 23681 37599 23715
rect 37657 23681 37691 23715
rect 1409 23613 1443 23647
rect 1685 23613 1719 23647
rect 3157 23613 3191 23647
rect 3617 23613 3651 23647
rect 8861 23613 8895 23647
rect 9689 23613 9723 23647
rect 11621 23613 11655 23647
rect 13921 23613 13955 23647
rect 18797 23613 18831 23647
rect 19901 23613 19935 23647
rect 24133 23613 24167 23647
rect 27721 23613 27755 23647
rect 30021 23613 30055 23647
rect 36737 23613 36771 23647
rect 3801 23545 3835 23579
rect 8217 23545 8251 23579
rect 13737 23545 13771 23579
rect 14657 23545 14691 23579
rect 15025 23545 15059 23579
rect 19809 23545 19843 23579
rect 21189 23545 21223 23579
rect 24317 23545 24351 23579
rect 3985 23477 4019 23511
rect 17417 23477 17451 23511
rect 18705 23477 18739 23511
rect 20545 23477 20579 23511
rect 21833 23477 21867 23511
rect 24225 23477 24259 23511
rect 24501 23477 24535 23511
rect 25237 23477 25271 23511
rect 28089 23477 28123 23511
rect 36829 23477 36863 23511
rect 2145 23273 2179 23307
rect 5181 23273 5215 23307
rect 5365 23273 5399 23307
rect 10701 23273 10735 23307
rect 18705 23273 18739 23307
rect 20545 23273 20579 23307
rect 28089 23273 28123 23307
rect 28273 23273 28307 23307
rect 31493 23273 31527 23307
rect 32137 23273 32171 23307
rect 32965 23273 32999 23307
rect 36369 23273 36403 23307
rect 36921 23273 36955 23307
rect 37657 23273 37691 23307
rect 4813 23205 4847 23239
rect 23949 23205 23983 23239
rect 30113 23205 30147 23239
rect 37841 23205 37875 23239
rect 5917 23137 5951 23171
rect 8953 23137 8987 23171
rect 16405 23137 16439 23171
rect 18613 23137 18647 23171
rect 19809 23137 19843 23171
rect 21281 23137 21315 23171
rect 22845 23137 22879 23171
rect 24409 23137 24443 23171
rect 27353 23137 27387 23171
rect 28181 23137 28215 23171
rect 29837 23137 29871 23171
rect 36829 23137 36863 23171
rect 2145 23069 2179 23103
rect 2329 23069 2363 23103
rect 2973 23069 3007 23103
rect 3157 23069 3191 23103
rect 4077 23069 4111 23103
rect 5089 23069 5123 23103
rect 5825 23069 5859 23103
rect 6009 23069 6043 23103
rect 6101 23069 6135 23103
rect 6469 23069 6503 23103
rect 6653 23069 6687 23103
rect 6745 23069 6779 23103
rect 6837 23069 6871 23103
rect 8309 23069 8343 23103
rect 8585 23069 8619 23103
rect 18889 23069 18923 23103
rect 19349 23069 19383 23103
rect 19625 23069 19659 23103
rect 19901 23069 19935 23103
rect 19993 23069 20027 23103
rect 20177 23069 20211 23103
rect 20361 23069 20395 23103
rect 21097 23069 21131 23103
rect 22109 23069 22143 23103
rect 22201 23069 22235 23103
rect 23949 23069 23983 23103
rect 24225 23069 24259 23103
rect 26433 23069 26467 23103
rect 26709 23069 26743 23103
rect 26893 23069 26927 23103
rect 26985 23069 27019 23103
rect 27077 23069 27111 23103
rect 27445 23069 27479 23103
rect 27537 23069 27571 23103
rect 27813 23069 27847 23103
rect 27905 23069 27939 23103
rect 28365 23069 28399 23103
rect 28457 23069 28491 23103
rect 28549 23069 28583 23103
rect 29745 23069 29779 23103
rect 31677 23069 31711 23103
rect 31769 23069 31803 23103
rect 31953 23069 31987 23103
rect 32137 23069 32171 23103
rect 33149 23069 33183 23103
rect 33241 23069 33275 23103
rect 36553 23069 36587 23103
rect 36737 23069 36771 23103
rect 36921 23069 36955 23103
rect 37105 23069 37139 23103
rect 37197 23069 37231 23103
rect 37473 23069 37507 23103
rect 37933 23069 37967 23103
rect 4721 23001 4755 23035
rect 4813 23001 4847 23035
rect 5349 23001 5383 23035
rect 5549 23001 5583 23035
rect 9229 23001 9263 23035
rect 16221 23001 16255 23035
rect 19073 23001 19107 23035
rect 20269 23001 20303 23035
rect 21005 23001 21039 23035
rect 24685 23001 24719 23035
rect 27721 23001 27755 23035
rect 28641 23001 28675 23035
rect 3065 22933 3099 22967
rect 4997 22933 5031 22967
rect 5641 22933 5675 22967
rect 7113 22933 7147 22967
rect 8401 22933 8435 22967
rect 8769 22933 8803 22967
rect 12081 22933 12115 22967
rect 15761 22933 15795 22967
rect 16129 22933 16163 22967
rect 19441 22933 19475 22967
rect 24133 22933 24167 22967
rect 37289 22933 37323 22967
rect 8493 22729 8527 22763
rect 8877 22729 8911 22763
rect 9045 22729 9079 22763
rect 11713 22729 11747 22763
rect 12357 22729 12391 22763
rect 12633 22729 12667 22763
rect 12817 22729 12851 22763
rect 19349 22729 19383 22763
rect 20269 22729 20303 22763
rect 21005 22729 21039 22763
rect 21925 22729 21959 22763
rect 25329 22729 25363 22763
rect 26801 22729 26835 22763
rect 27629 22729 27663 22763
rect 28917 22729 28951 22763
rect 30205 22729 30239 22763
rect 30297 22729 30331 22763
rect 30849 22729 30883 22763
rect 32137 22729 32171 22763
rect 32597 22729 32631 22763
rect 33885 22729 33919 22763
rect 34529 22729 34563 22763
rect 34805 22729 34839 22763
rect 36093 22729 36127 22763
rect 36921 22729 36955 22763
rect 37841 22729 37875 22763
rect 37933 22729 37967 22763
rect 2329 22661 2363 22695
rect 6469 22661 6503 22695
rect 7021 22661 7055 22695
rect 8677 22661 8711 22695
rect 11989 22661 12023 22695
rect 23213 22661 23247 22695
rect 24961 22661 24995 22695
rect 28733 22661 28767 22695
rect 29193 22661 29227 22695
rect 29285 22661 29319 22695
rect 34957 22661 34991 22695
rect 35173 22661 35207 22695
rect 38085 22661 38119 22695
rect 38301 22661 38335 22695
rect 5825 22593 5859 22627
rect 6009 22593 6043 22627
rect 6377 22593 6411 22627
rect 6745 22593 6779 22627
rect 12173 22593 12207 22627
rect 19263 22593 19297 22627
rect 19441 22593 19475 22627
rect 19717 22593 19751 22627
rect 20177 22593 20211 22627
rect 20361 22593 20395 22627
rect 20637 22593 20671 22627
rect 21833 22593 21867 22627
rect 22109 22593 22143 22627
rect 25421 22593 25455 22627
rect 26249 22593 26283 22627
rect 26525 22593 26559 22627
rect 26617 22593 26651 22627
rect 27169 22593 27203 22627
rect 27997 22593 28031 22627
rect 28641 22593 28675 22627
rect 28825 22593 28859 22627
rect 29101 22593 29135 22627
rect 29423 22593 29457 22627
rect 30021 22593 30055 22627
rect 30511 22593 30545 22627
rect 30665 22593 30699 22627
rect 30757 22593 30791 22627
rect 31033 22593 31067 22627
rect 32137 22593 32171 22627
rect 32321 22593 32355 22627
rect 32505 22593 32539 22627
rect 32689 22593 32723 22627
rect 33149 22593 33183 22627
rect 33701 22593 33735 22627
rect 34437 22593 34471 22627
rect 34621 22593 34655 22627
rect 35265 22593 35299 22627
rect 35357 22593 35391 22627
rect 35541 22593 35575 22627
rect 36001 22593 36035 22627
rect 36185 22593 36219 22627
rect 36277 22593 36311 22627
rect 36461 22593 36495 22627
rect 36737 22593 36771 22627
rect 37657 22593 37691 22627
rect 2053 22525 2087 22559
rect 3893 22525 3927 22559
rect 4169 22525 4203 22559
rect 5733 22525 5767 22559
rect 13553 22525 13587 22559
rect 19533 22525 19567 22559
rect 22293 22525 22327 22559
rect 22937 22525 22971 22559
rect 27353 22525 27387 22559
rect 27537 22525 27571 22559
rect 28089 22525 28123 22559
rect 29561 22525 29595 22559
rect 29745 22525 29779 22559
rect 29837 22525 29871 22559
rect 33057 22525 33091 22559
rect 33425 22525 33459 22559
rect 36369 22525 36403 22559
rect 36553 22525 36587 22559
rect 37381 22525 37415 22559
rect 27261 22457 27295 22491
rect 31033 22457 31067 22491
rect 33517 22457 33551 22491
rect 35541 22457 35575 22491
rect 3801 22389 3835 22423
rect 5641 22389 5675 22423
rect 6193 22389 6227 22423
rect 8861 22389 8895 22423
rect 12909 22389 12943 22423
rect 19901 22389 19935 22423
rect 21005 22389 21039 22423
rect 21189 22389 21223 22423
rect 22201 22389 22235 22423
rect 22569 22389 22603 22423
rect 26341 22389 26375 22423
rect 27353 22389 27387 22423
rect 32781 22389 32815 22423
rect 34989 22389 35023 22423
rect 37473 22389 37507 22423
rect 38117 22389 38151 22423
rect 5365 22185 5399 22219
rect 5904 22185 5938 22219
rect 7389 22185 7423 22219
rect 14933 22185 14967 22219
rect 15380 22185 15414 22219
rect 22550 22185 22584 22219
rect 28273 22185 28307 22219
rect 28641 22185 28675 22219
rect 30113 22185 30147 22219
rect 32045 22185 32079 22219
rect 32597 22185 32631 22219
rect 33241 22185 33275 22219
rect 34437 22185 34471 22219
rect 34713 22185 34747 22219
rect 36553 22185 36587 22219
rect 37841 22185 37875 22219
rect 4353 22049 4387 22083
rect 8401 22049 8435 22083
rect 8677 22049 8711 22083
rect 12081 22049 12115 22083
rect 12173 22049 12207 22083
rect 13921 22049 13955 22083
rect 17141 22049 17175 22083
rect 18981 22049 19015 22083
rect 22293 22049 22327 22083
rect 27077 22049 27111 22083
rect 30481 22049 30515 22083
rect 35541 22049 35575 22083
rect 37289 22049 37323 22083
rect 3065 21981 3099 22015
rect 5181 21981 5215 22015
rect 5641 21981 5675 22015
rect 8309 21981 8343 22015
rect 8953 21981 8987 22015
rect 9505 21981 9539 22015
rect 15117 21981 15151 22015
rect 20080 21981 20114 22015
rect 20452 21981 20486 22015
rect 20545 21981 20579 22015
rect 21189 21981 21223 22015
rect 21347 21981 21381 22015
rect 21649 21981 21683 22015
rect 21833 21981 21867 22015
rect 26985 21981 27019 22015
rect 28089 21981 28123 22015
rect 28273 21981 28307 22015
rect 28457 21981 28491 22015
rect 28641 21981 28675 22015
rect 30297 21981 30331 22015
rect 32505 21981 32539 22015
rect 32689 21981 32723 22015
rect 32873 21981 32907 22015
rect 34345 21981 34379 22015
rect 34529 21981 34563 22015
rect 35081 21981 35115 22015
rect 35173 21981 35207 22015
rect 35357 21981 35391 22015
rect 36921 21981 36955 22015
rect 37197 21981 37231 22015
rect 37381 21981 37415 22015
rect 37657 21981 37691 22015
rect 11805 21913 11839 21947
rect 12449 21913 12483 21947
rect 18705 21913 18739 21947
rect 20177 21913 20211 21947
rect 20269 21913 20303 21947
rect 21465 21913 21499 21947
rect 21557 21913 21591 21947
rect 32229 21913 32263 21947
rect 32413 21913 32447 21947
rect 33057 21913 33091 21947
rect 34897 21913 34931 21947
rect 36737 21913 36771 21947
rect 37473 21913 37507 21947
rect 2881 21845 2915 21879
rect 10333 21845 10367 21879
rect 17233 21845 17267 21879
rect 19901 21845 19935 21879
rect 24041 21845 24075 21879
rect 4353 21641 4387 21675
rect 6009 21641 6043 21675
rect 8769 21641 8803 21675
rect 11069 21641 11103 21675
rect 11805 21641 11839 21675
rect 13185 21641 13219 21675
rect 17601 21641 17635 21675
rect 21833 21641 21867 21675
rect 26433 21641 26467 21675
rect 29101 21641 29135 21675
rect 33977 21641 34011 21675
rect 35081 21641 35115 21675
rect 35357 21641 35391 21675
rect 3985 21573 4019 21607
rect 5089 21573 5123 21607
rect 10241 21573 10275 21607
rect 12173 21573 12207 21607
rect 12265 21573 12299 21607
rect 13553 21573 13587 21607
rect 34713 21573 34747 21607
rect 3801 21505 3835 21539
rect 4077 21505 4111 21539
rect 4537 21505 4571 21539
rect 4813 21505 4847 21539
rect 4997 21505 5031 21539
rect 5733 21505 5767 21539
rect 5825 21505 5859 21539
rect 6377 21505 6411 21539
rect 6561 21505 6595 21539
rect 10977 21505 11011 21539
rect 12633 21505 12667 21539
rect 12817 21505 12851 21539
rect 12909 21505 12943 21539
rect 13645 21505 13679 21539
rect 14197 21505 14231 21539
rect 17233 21505 17267 21539
rect 17693 21505 17727 21539
rect 20637 21505 20671 21539
rect 22201 21505 22235 21539
rect 22293 21505 22327 21539
rect 22477 21505 22511 21539
rect 25053 21505 25087 21539
rect 25789 21505 25823 21539
rect 25881 21505 25915 21539
rect 26341 21505 26375 21539
rect 26985 21505 27019 21539
rect 27169 21505 27203 21539
rect 28917 21505 28951 21539
rect 29285 21505 29319 21539
rect 29469 21505 29503 21539
rect 30021 21505 30055 21539
rect 30205 21505 30239 21539
rect 32321 21505 32355 21539
rect 33885 21505 33919 21539
rect 34069 21505 34103 21539
rect 34897 21505 34931 21539
rect 35173 21505 35207 21539
rect 35357 21505 35391 21539
rect 8585 21437 8619 21471
rect 10517 21437 10551 21471
rect 11161 21437 11195 21471
rect 12449 21437 12483 21471
rect 13737 21437 13771 21471
rect 14473 21437 14507 21471
rect 17049 21437 17083 21471
rect 17141 21437 17175 21471
rect 18245 21437 18279 21471
rect 22017 21437 22051 21471
rect 22109 21437 22143 21471
rect 25145 21437 25179 21471
rect 25329 21437 25363 21471
rect 28733 21437 28767 21471
rect 32229 21437 32263 21471
rect 32689 21437 32723 21471
rect 6377 21369 6411 21403
rect 26065 21369 26099 21403
rect 8033 21301 8067 21335
rect 10609 21301 10643 21335
rect 12817 21301 12851 21335
rect 13093 21301 13127 21335
rect 15945 21301 15979 21335
rect 20361 21301 20395 21335
rect 20913 21301 20947 21335
rect 22569 21301 22603 21335
rect 24685 21301 24719 21335
rect 25605 21301 25639 21335
rect 27077 21301 27111 21335
rect 29469 21301 29503 21335
rect 30389 21301 30423 21335
rect 7573 21097 7607 21131
rect 13461 21097 13495 21131
rect 13645 21097 13679 21131
rect 14749 21097 14783 21131
rect 17969 21097 18003 21131
rect 21005 21097 21039 21131
rect 21741 21097 21775 21131
rect 22385 21097 22419 21131
rect 26341 21097 26375 21131
rect 28273 21097 28307 21131
rect 29653 21097 29687 21131
rect 31769 21097 31803 21131
rect 32597 21097 32631 21131
rect 33793 21097 33827 21131
rect 34345 21097 34379 21131
rect 35909 21097 35943 21131
rect 36737 21097 36771 21131
rect 37565 21097 37599 21131
rect 7941 21029 7975 21063
rect 14289 21029 14323 21063
rect 16221 21029 16255 21063
rect 18521 21029 18555 21063
rect 21557 21029 21591 21063
rect 36369 21029 36403 21063
rect 38117 21029 38151 21063
rect 5641 20961 5675 20995
rect 8585 20961 8619 20995
rect 10701 20961 10735 20995
rect 13737 20961 13771 20995
rect 14381 20961 14415 20995
rect 15209 20961 15243 20995
rect 15301 20961 15335 20995
rect 16957 20961 16991 20995
rect 17877 20961 17911 20995
rect 18705 20961 18739 20995
rect 19257 20961 19291 20995
rect 24409 20961 24443 20995
rect 24777 20961 24811 20995
rect 26893 20961 26927 20995
rect 29101 20961 29135 20995
rect 38301 20961 38335 20995
rect 2881 20893 2915 20927
rect 3065 20893 3099 20927
rect 7389 20893 7423 20927
rect 7573 20893 7607 20927
rect 7665 20893 7699 20927
rect 7941 20893 7975 20927
rect 10425 20893 10459 20927
rect 12725 20893 12759 20927
rect 12909 20893 12943 20927
rect 13185 20893 13219 20927
rect 14197 20893 14231 20927
rect 14473 20893 14507 20927
rect 15577 20893 15611 20927
rect 15761 20893 15795 20927
rect 16037 20893 16071 20927
rect 17969 20893 18003 20927
rect 18061 20893 18095 20927
rect 18429 20893 18463 20927
rect 21833 20893 21867 20927
rect 22109 20893 22143 20927
rect 22385 20893 22419 20927
rect 22753 20893 22787 20927
rect 22845 20893 22879 20927
rect 23029 20893 23063 20927
rect 23305 20893 23339 20927
rect 26801 20893 26835 20927
rect 27169 20893 27203 20927
rect 27353 20893 27387 20927
rect 28089 20893 28123 20927
rect 28181 20893 28215 20927
rect 28365 20893 28399 20927
rect 28641 20893 28675 20927
rect 28825 20893 28859 20927
rect 28917 20893 28951 20927
rect 29009 20893 29043 20927
rect 29193 20893 29227 20927
rect 29561 20893 29595 20927
rect 30021 20893 30055 20927
rect 31401 20893 31435 20927
rect 31585 20893 31619 20927
rect 31677 20893 31711 20927
rect 31861 20893 31895 20927
rect 32321 20893 32355 20927
rect 32413 20893 32447 20927
rect 32689 20893 32723 20927
rect 33701 20893 33735 20927
rect 33885 20893 33919 20927
rect 33977 20893 34011 20927
rect 34161 20893 34195 20927
rect 35817 20893 35851 20927
rect 36001 20893 36035 20927
rect 36093 20893 36127 20927
rect 36369 20893 36403 20927
rect 36507 20893 36541 20927
rect 36645 20893 36679 20927
rect 36829 20893 36863 20927
rect 37841 20893 37875 20927
rect 37933 20893 37967 20927
rect 38117 20893 38151 20927
rect 38209 20893 38243 20927
rect 38393 20893 38427 20927
rect 3525 20825 3559 20859
rect 5365 20825 5399 20859
rect 8033 20825 8067 20859
rect 13461 20825 13495 20859
rect 13829 20825 13863 20859
rect 14657 20825 14691 20859
rect 16773 20825 16807 20859
rect 17233 20825 17267 20859
rect 19533 20825 19567 20859
rect 23213 20825 23247 20859
rect 26249 20825 26283 20859
rect 27537 20825 27571 20859
rect 27721 20825 27755 20859
rect 27905 20825 27939 20859
rect 29837 20825 29871 20859
rect 31493 20825 31527 20859
rect 31953 20825 31987 20859
rect 32873 20825 32907 20859
rect 33057 20825 33091 20859
rect 37549 20825 37583 20859
rect 37749 20825 37783 20859
rect 2973 20757 3007 20791
rect 3433 20757 3467 20791
rect 3893 20757 3927 20791
rect 7757 20757 7791 20791
rect 12173 20757 12207 20791
rect 13369 20757 13403 20791
rect 15117 20757 15151 20791
rect 16405 20757 16439 20791
rect 16865 20757 16899 20791
rect 18337 20757 18371 20791
rect 18705 20757 18739 20791
rect 19073 20757 19107 20791
rect 22201 20757 22235 20791
rect 26709 20757 26743 20791
rect 28457 20757 28491 20791
rect 30205 20757 30239 20791
rect 37381 20757 37415 20791
rect 5365 20553 5399 20587
rect 7941 20553 7975 20587
rect 11621 20553 11655 20587
rect 15945 20553 15979 20587
rect 17325 20553 17359 20587
rect 18337 20553 18371 20587
rect 25329 20553 25363 20587
rect 25973 20553 26007 20587
rect 27261 20553 27295 20587
rect 34437 20553 34471 20587
rect 35541 20553 35575 20587
rect 37105 20553 37139 20587
rect 37841 20553 37875 20587
rect 2513 20485 2547 20519
rect 4905 20485 4939 20519
rect 9413 20485 9447 20519
rect 12817 20485 12851 20519
rect 16405 20485 16439 20519
rect 17693 20485 17727 20519
rect 18153 20485 18187 20519
rect 21189 20485 21223 20519
rect 23857 20485 23891 20519
rect 25513 20485 25547 20519
rect 25697 20485 25731 20519
rect 27077 20485 27111 20519
rect 29653 20485 29687 20519
rect 37473 20485 37507 20519
rect 37657 20485 37691 20519
rect 2237 20417 2271 20451
rect 5549 20417 5583 20451
rect 5825 20417 5859 20451
rect 6009 20417 6043 20451
rect 6929 20417 6963 20451
rect 7205 20417 7239 20451
rect 7757 20417 7791 20451
rect 9689 20417 9723 20451
rect 12265 20417 12299 20451
rect 13645 20417 13679 20451
rect 15853 20417 15887 20451
rect 16497 20417 16531 20451
rect 16681 20417 16715 20451
rect 17601 20417 17635 20451
rect 18521 20417 18555 20451
rect 18613 20417 18647 20451
rect 18705 20417 18739 20451
rect 18843 20417 18877 20451
rect 19073 20417 19107 20451
rect 21465 20417 21499 20451
rect 21833 20417 21867 20451
rect 22109 20417 22143 20451
rect 22385 20417 22419 20451
rect 23121 20417 23155 20451
rect 23213 20417 23247 20451
rect 23305 20417 23339 20451
rect 23489 20417 23523 20451
rect 26157 20417 26191 20451
rect 26341 20417 26375 20451
rect 26433 20417 26467 20451
rect 26525 20417 26559 20451
rect 27169 20417 27203 20451
rect 27261 20417 27295 20451
rect 27445 20417 27479 20451
rect 27905 20417 27939 20451
rect 28089 20417 28123 20451
rect 30021 20417 30055 20451
rect 30205 20417 30239 20451
rect 31585 20417 31619 20451
rect 31769 20417 31803 20451
rect 33517 20417 33551 20451
rect 33977 20417 34011 20451
rect 34069 20417 34103 20451
rect 34253 20417 34287 20451
rect 35909 20417 35943 20451
rect 36369 20417 36403 20451
rect 36645 20417 36679 20451
rect 36921 20417 36955 20451
rect 4629 20349 4663 20383
rect 5733 20349 5767 20383
rect 5917 20349 5951 20383
rect 7021 20349 7055 20383
rect 13001 20349 13035 20383
rect 13921 20349 13955 20383
rect 16037 20349 16071 20383
rect 18981 20349 19015 20383
rect 19349 20349 19383 20383
rect 21281 20349 21315 20383
rect 21925 20349 21959 20383
rect 22477 20349 22511 20383
rect 22937 20349 22971 20383
rect 23397 20349 23431 20383
rect 23581 20349 23615 20383
rect 27997 20349 28031 20383
rect 33609 20349 33643 20383
rect 33885 20349 33919 20383
rect 35817 20349 35851 20383
rect 36461 20349 36495 20383
rect 18153 20281 18187 20315
rect 21649 20281 21683 20315
rect 3985 20213 4019 20247
rect 4077 20213 4111 20247
rect 4997 20213 5031 20247
rect 6561 20213 6595 20247
rect 13553 20213 13587 20247
rect 15393 20213 15427 20247
rect 15485 20213 15519 20247
rect 17417 20213 17451 20247
rect 20821 20213 20855 20247
rect 21189 20213 21223 20247
rect 22293 20213 22327 20247
rect 22569 20213 22603 20247
rect 22753 20213 22787 20247
rect 23029 20213 23063 20247
rect 26801 20213 26835 20247
rect 29561 20213 29595 20247
rect 30205 20213 30239 20247
rect 31585 20213 31619 20247
rect 35909 20213 35943 20247
rect 36001 20213 36035 20247
rect 36737 20213 36771 20247
rect 3433 20009 3467 20043
rect 3801 20009 3835 20043
rect 4445 20009 4479 20043
rect 8125 20009 8159 20043
rect 8401 20009 8435 20043
rect 8585 20009 8619 20043
rect 13921 20009 13955 20043
rect 14289 20009 14323 20043
rect 17509 20009 17543 20043
rect 19809 20009 19843 20043
rect 21741 20009 21775 20043
rect 22845 20009 22879 20043
rect 23489 20009 23523 20043
rect 28089 20009 28123 20043
rect 29193 20009 29227 20043
rect 36461 20009 36495 20043
rect 36921 20009 36955 20043
rect 3249 19941 3283 19975
rect 22937 19941 22971 19975
rect 31815 19941 31849 19975
rect 33609 19941 33643 19975
rect 1409 19873 1443 19907
rect 6285 19873 6319 19907
rect 6377 19873 6411 19907
rect 6653 19873 6687 19907
rect 10609 19873 10643 19907
rect 12541 19873 12575 19907
rect 13369 19873 13403 19907
rect 13461 19873 13495 19907
rect 16037 19873 16071 19907
rect 17693 19873 17727 19907
rect 22201 19873 22235 19907
rect 22661 19873 22695 19907
rect 29377 19873 29411 19907
rect 29561 19873 29595 19907
rect 30021 19873 30055 19907
rect 34437 19873 34471 19907
rect 36001 19873 36035 19907
rect 36645 19873 36679 19907
rect 3985 19805 4019 19839
rect 4261 19805 4295 19839
rect 14381 19805 14415 19839
rect 14749 19805 14783 19839
rect 15761 19805 15795 19839
rect 17601 19805 17635 19839
rect 17785 19805 17819 19839
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 19533 19805 19567 19839
rect 19625 19805 19659 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 22569 19805 22603 19839
rect 23062 19805 23096 19839
rect 23581 19805 23615 19839
rect 25973 19805 26007 19839
rect 26065 19805 26099 19839
rect 26249 19805 26283 19839
rect 26341 19805 26375 19839
rect 27537 19805 27571 19839
rect 27813 19805 27847 19839
rect 27905 19805 27939 19839
rect 28825 19805 28859 19839
rect 29101 19805 29135 19839
rect 29745 19805 29779 19839
rect 30389 19805 30423 19839
rect 32413 19805 32447 19839
rect 32591 19805 32625 19839
rect 33823 19805 33857 19839
rect 33977 19805 34011 19839
rect 36185 19805 36219 19839
rect 36277 19805 36311 19839
rect 36369 19805 36403 19839
rect 1685 19737 1719 19771
rect 3617 19737 3651 19771
rect 4077 19737 4111 19771
rect 6009 19737 6043 19771
rect 8217 19737 8251 19771
rect 12265 19737 12299 19771
rect 15485 19737 15519 19771
rect 27721 19737 27755 19771
rect 28733 19737 28767 19771
rect 34069 19737 34103 19771
rect 34253 19737 34287 19771
rect 36001 19737 36035 19771
rect 3157 19669 3191 19703
rect 3417 19669 3451 19703
rect 4537 19669 4571 19703
rect 8401 19669 8435 19703
rect 9965 19669 9999 19703
rect 10333 19669 10367 19703
rect 10425 19669 10459 19703
rect 10793 19669 10827 19703
rect 13553 19669 13587 19703
rect 22109 19669 22143 19703
rect 23121 19669 23155 19703
rect 23673 19669 23707 19703
rect 26525 19669 26559 19703
rect 29377 19669 29411 19703
rect 29929 19669 29963 19703
rect 32505 19669 32539 19703
rect 21557 19465 21591 19499
rect 25881 19465 25915 19499
rect 28457 19465 28491 19499
rect 33425 19465 33459 19499
rect 33977 19465 34011 19499
rect 35633 19465 35667 19499
rect 36369 19465 36403 19499
rect 36829 19465 36863 19499
rect 3709 19397 3743 19431
rect 11805 19397 11839 19431
rect 12725 19397 12759 19431
rect 13461 19397 13495 19431
rect 14197 19397 14231 19431
rect 18797 19397 18831 19431
rect 21833 19397 21867 19431
rect 24317 19397 24351 19431
rect 25237 19397 25271 19431
rect 28089 19397 28123 19431
rect 28181 19397 28215 19431
rect 29285 19397 29319 19431
rect 29377 19397 29411 19431
rect 29929 19397 29963 19431
rect 30113 19397 30147 19431
rect 31677 19397 31711 19431
rect 31861 19397 31895 19431
rect 32229 19397 32263 19431
rect 32505 19397 32539 19431
rect 32689 19397 32723 19431
rect 35817 19397 35851 19431
rect 36185 19397 36219 19431
rect 36921 19397 36955 19431
rect 2145 19329 2179 19363
rect 2697 19329 2731 19363
rect 3433 19329 3467 19363
rect 3525 19329 3559 19363
rect 4261 19329 4295 19363
rect 4721 19329 4755 19363
rect 7481 19329 7515 19363
rect 7665 19329 7699 19363
rect 11897 19329 11931 19363
rect 12909 19329 12943 19363
rect 13185 19329 13219 19363
rect 13369 19329 13403 19363
rect 14105 19329 14139 19363
rect 14473 19329 14507 19363
rect 14749 19329 14783 19363
rect 16681 19329 16715 19363
rect 18521 19329 18555 19363
rect 18705 19329 18739 19363
rect 18889 19329 18923 19363
rect 19533 19329 19567 19363
rect 23673 19329 23707 19363
rect 23857 19329 23891 19363
rect 23949 19329 23983 19363
rect 24041 19329 24075 19363
rect 24685 19329 24719 19363
rect 25145 19329 25179 19363
rect 25329 19329 25363 19363
rect 25789 19329 25823 19363
rect 25973 19329 26007 19363
rect 26985 19329 27019 19363
rect 27169 19329 27203 19363
rect 27537 19329 27571 19363
rect 27813 19329 27847 19363
rect 27906 19329 27940 19363
rect 28319 19329 28353 19363
rect 29101 19329 29135 19363
rect 29469 19329 29503 19363
rect 32137 19329 32171 19363
rect 32321 19329 32355 19363
rect 33241 19329 33275 19363
rect 33517 19329 33551 19363
rect 33793 19329 33827 19363
rect 34621 19329 34655 19363
rect 35541 19329 35575 19363
rect 35725 19329 35759 19363
rect 36001 19329 36035 19363
rect 36277 19329 36311 19363
rect 36553 19329 36587 19363
rect 36829 19329 36863 19363
rect 37105 19329 37139 19363
rect 1777 19261 1811 19295
rect 2237 19261 2271 19295
rect 3341 19261 3375 19295
rect 4353 19261 4387 19295
rect 5273 19261 5307 19295
rect 9505 19261 9539 19295
rect 9781 19261 9815 19295
rect 11253 19261 11287 19295
rect 11621 19261 11655 19295
rect 14289 19261 14323 19295
rect 15025 19261 15059 19295
rect 16497 19261 16531 19295
rect 19809 19261 19843 19295
rect 24777 19261 24811 19295
rect 27261 19261 27295 19295
rect 27353 19261 27387 19295
rect 27721 19261 27755 19295
rect 33609 19261 33643 19295
rect 36737 19261 36771 19295
rect 3709 19193 3743 19227
rect 4629 19193 4663 19227
rect 12265 19193 12299 19227
rect 25053 19193 25087 19227
rect 29653 19193 29687 19227
rect 7665 19125 7699 19159
rect 14197 19125 14231 19159
rect 14657 19125 14691 19159
rect 16865 19125 16899 19159
rect 19073 19125 19107 19159
rect 21281 19125 21315 19159
rect 23121 19125 23155 19159
rect 30297 19125 30331 19159
rect 31493 19125 31527 19159
rect 32781 19125 32815 19159
rect 33057 19125 33091 19159
rect 34805 19125 34839 19159
rect 3433 18921 3467 18955
rect 3893 18921 3927 18955
rect 4169 18921 4203 18955
rect 4629 18921 4663 18955
rect 8493 18921 8527 18955
rect 13093 18921 13127 18955
rect 14657 18921 14691 18955
rect 16129 18921 16163 18955
rect 17049 18921 17083 18955
rect 23581 18921 23615 18955
rect 25145 18921 25179 18955
rect 27445 18921 27479 18955
rect 28733 18921 28767 18955
rect 34897 18921 34931 18955
rect 36001 18921 36035 18955
rect 3617 18853 3651 18887
rect 4261 18853 4295 18887
rect 17233 18853 17267 18887
rect 25605 18853 25639 18887
rect 31769 18853 31803 18887
rect 33701 18853 33735 18887
rect 34713 18853 34747 18887
rect 36185 18853 36219 18887
rect 36829 18853 36863 18887
rect 37289 18853 37323 18887
rect 6929 18785 6963 18819
rect 13185 18785 13219 18819
rect 15945 18785 15979 18819
rect 16773 18785 16807 18819
rect 19717 18785 19751 18819
rect 22385 18785 22419 18819
rect 23305 18785 23339 18819
rect 25513 18785 25547 18819
rect 25697 18785 25731 18819
rect 28365 18785 28399 18819
rect 31861 18785 31895 18819
rect 33149 18785 33183 18819
rect 34161 18785 34195 18819
rect 34253 18785 34287 18819
rect 3249 18717 3283 18751
rect 3433 18717 3467 18751
rect 4077 18717 4111 18751
rect 4353 18717 4387 18751
rect 4629 18717 4663 18751
rect 4721 18717 4755 18751
rect 6653 18717 6687 18751
rect 8493 18717 8527 18751
rect 8677 18717 8711 18751
rect 9137 18717 9171 18751
rect 12449 18717 12483 18751
rect 12633 18717 12667 18751
rect 12909 18717 12943 18751
rect 13369 18717 13403 18751
rect 13645 18717 13679 18751
rect 13829 18717 13863 18751
rect 14105 18717 14139 18751
rect 14289 18717 14323 18751
rect 15025 18717 15059 18751
rect 15209 18717 15243 18751
rect 15669 18717 15703 18751
rect 17325 18717 17359 18751
rect 17509 18717 17543 18751
rect 17693 18717 17727 18751
rect 18521 18717 18555 18751
rect 19441 18717 19475 18751
rect 21557 18717 21591 18751
rect 21741 18717 21775 18751
rect 22109 18717 22143 18751
rect 22569 18717 22603 18751
rect 23029 18717 23063 18751
rect 23857 18717 23891 18751
rect 24041 18717 24075 18751
rect 24133 18717 24167 18751
rect 24869 18717 24903 18751
rect 25329 18717 25363 18751
rect 25421 18717 25455 18751
rect 26893 18717 26927 18751
rect 27077 18717 27111 18751
rect 27353 18717 27387 18751
rect 27629 18717 27663 18751
rect 27997 18717 28031 18751
rect 28181 18717 28215 18751
rect 28273 18717 28307 18751
rect 28549 18717 28583 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 29193 18717 29227 18751
rect 29561 18717 29595 18751
rect 29745 18717 29779 18751
rect 32137 18717 32171 18751
rect 32413 18717 32447 18751
rect 32781 18717 32815 18751
rect 33425 18717 33459 18751
rect 33977 18717 34011 18751
rect 34345 18717 34379 18751
rect 34529 18717 34563 18751
rect 35909 18717 35943 18751
rect 36093 18717 36127 18751
rect 36553 18717 36587 18751
rect 36645 18717 36679 18751
rect 9413 18649 9447 18683
rect 15117 18649 15151 18683
rect 16865 18649 16899 18683
rect 17065 18649 17099 18683
rect 17601 18649 17635 18683
rect 17969 18649 18003 18683
rect 21465 18649 21499 18683
rect 22017 18649 22051 18683
rect 23397 18649 23431 18683
rect 23597 18649 23631 18683
rect 24961 18649 24995 18683
rect 26985 18649 27019 18683
rect 27215 18649 27249 18683
rect 27813 18649 27847 18683
rect 29101 18649 29135 18683
rect 31401 18649 31435 18683
rect 31585 18649 31619 18683
rect 33701 18649 33735 18683
rect 34865 18649 34899 18683
rect 35081 18649 35115 18683
rect 36369 18649 36403 18683
rect 37105 18649 37139 18683
rect 4445 18581 4479 18615
rect 4997 18581 5031 18615
rect 8401 18581 8435 18615
rect 10885 18581 10919 18615
rect 14197 18581 14231 18615
rect 15301 18581 15335 18615
rect 15761 18581 15795 18615
rect 17877 18581 17911 18615
rect 23765 18581 23799 18615
rect 24133 18581 24167 18615
rect 26709 18581 26743 18615
rect 29377 18581 29411 18615
rect 29653 18581 29687 18615
rect 33517 18581 33551 18615
rect 33793 18581 33827 18615
rect 4537 18377 4571 18411
rect 7849 18377 7883 18411
rect 9137 18377 9171 18411
rect 10057 18377 10091 18411
rect 10517 18377 10551 18411
rect 13737 18377 13771 18411
rect 14289 18377 14323 18411
rect 16497 18377 16531 18411
rect 22569 18377 22603 18411
rect 24409 18377 24443 18411
rect 25421 18377 25455 18411
rect 28181 18377 28215 18411
rect 28457 18377 28491 18411
rect 31769 18377 31803 18411
rect 7481 18309 7515 18343
rect 7697 18309 7731 18343
rect 15025 18309 15059 18343
rect 17141 18309 17175 18343
rect 17371 18309 17405 18343
rect 18245 18309 18279 18343
rect 27813 18309 27847 18343
rect 31401 18309 31435 18343
rect 35081 18309 35115 18343
rect 3525 18241 3559 18275
rect 3985 18241 4019 18275
rect 4353 18241 4387 18275
rect 4905 18241 4939 18275
rect 4997 18241 5031 18275
rect 5181 18241 5215 18275
rect 5273 18241 5307 18275
rect 6009 18241 6043 18275
rect 6193 18241 6227 18275
rect 8125 18241 8159 18275
rect 8309 18241 8343 18275
rect 8493 18241 8527 18275
rect 9229 18241 9263 18275
rect 9413 18241 9447 18275
rect 10425 18241 10459 18275
rect 12633 18241 12667 18275
rect 12909 18241 12943 18275
rect 13277 18241 13311 18275
rect 13553 18241 13587 18275
rect 13829 18241 13863 18275
rect 14105 18241 14139 18275
rect 14657 18241 14691 18275
rect 14749 18241 14783 18275
rect 17049 18241 17083 18275
rect 17233 18241 17267 18275
rect 17509 18241 17543 18275
rect 17969 18241 18003 18275
rect 19993 18241 20027 18275
rect 22201 18241 22235 18275
rect 23581 18241 23615 18275
rect 24225 18241 24259 18275
rect 24961 18241 24995 18275
rect 25605 18241 25639 18275
rect 25697 18241 25731 18275
rect 27629 18241 27663 18275
rect 28089 18241 28123 18275
rect 28365 18241 28399 18275
rect 28549 18241 28583 18275
rect 29009 18241 29043 18275
rect 29837 18241 29871 18275
rect 30021 18241 30055 18275
rect 30205 18241 30239 18275
rect 30389 18241 30423 18275
rect 30573 18241 30607 18275
rect 31125 18241 31159 18275
rect 31218 18241 31252 18275
rect 31493 18241 31527 18275
rect 31631 18241 31665 18275
rect 33425 18241 33459 18275
rect 33517 18241 33551 18275
rect 34345 18241 34379 18275
rect 34621 18241 34655 18275
rect 34989 18241 35023 18275
rect 35265 18241 35299 18275
rect 1501 18173 1535 18207
rect 1777 18173 1811 18207
rect 3249 18173 3283 18207
rect 3709 18173 3743 18207
rect 3893 18173 3927 18207
rect 5825 18173 5859 18207
rect 7941 18173 7975 18207
rect 9321 18173 9355 18207
rect 10701 18173 10735 18207
rect 12081 18173 12115 18207
rect 12817 18173 12851 18207
rect 14013 18173 14047 18207
rect 14381 18173 14415 18207
rect 17877 18173 17911 18207
rect 22293 18173 22327 18207
rect 23949 18173 23983 18207
rect 25053 18173 25087 18207
rect 25421 18173 25455 18207
rect 29101 18173 29135 18207
rect 30113 18173 30147 18207
rect 33241 18173 33275 18207
rect 33609 18173 33643 18207
rect 3341 18105 3375 18139
rect 5181 18105 5215 18139
rect 12725 18105 12759 18139
rect 13093 18105 13127 18139
rect 13369 18105 13403 18139
rect 13461 18105 13495 18139
rect 14473 18105 14507 18139
rect 33333 18105 33367 18139
rect 33885 18105 33919 18139
rect 4261 18037 4295 18071
rect 6193 18037 6227 18071
rect 7665 18037 7699 18071
rect 11529 18037 11563 18071
rect 13829 18037 13863 18071
rect 14565 18037 14599 18071
rect 16865 18037 16899 18071
rect 22201 18037 22235 18071
rect 23673 18037 23707 18071
rect 24041 18037 24075 18071
rect 25145 18037 25179 18071
rect 25329 18037 25363 18071
rect 27997 18037 28031 18071
rect 35449 18037 35483 18071
rect 2421 17833 2455 17867
rect 2789 17833 2823 17867
rect 4629 17833 4663 17867
rect 4813 17833 4847 17867
rect 8769 17833 8803 17867
rect 10793 17833 10827 17867
rect 12817 17833 12851 17867
rect 15853 17833 15887 17867
rect 18429 17833 18463 17867
rect 19809 17833 19843 17867
rect 24501 17833 24535 17867
rect 27261 17833 27295 17867
rect 30941 17833 30975 17867
rect 33241 17833 33275 17867
rect 33517 17833 33551 17867
rect 34161 17833 34195 17867
rect 37243 17833 37277 17867
rect 5089 17765 5123 17799
rect 7297 17765 7331 17799
rect 3065 17697 3099 17731
rect 6561 17697 6595 17731
rect 6837 17697 6871 17731
rect 7941 17697 7975 17731
rect 8125 17697 8159 17731
rect 10885 17697 10919 17731
rect 12633 17697 12667 17731
rect 13369 17697 13403 17731
rect 14105 17697 14139 17731
rect 16681 17697 16715 17731
rect 21281 17697 21315 17731
rect 23029 17697 23063 17731
rect 23673 17697 23707 17731
rect 32137 17697 32171 17731
rect 32229 17697 32263 17731
rect 35817 17697 35851 17731
rect 2605 17629 2639 17663
rect 2881 17629 2915 17663
rect 2973 17629 3007 17663
rect 3157 17629 3191 17663
rect 4445 17629 4479 17663
rect 7021 17629 7055 17663
rect 9045 17629 9079 17663
rect 12817 17629 12851 17663
rect 13001 17629 13035 17663
rect 13461 17629 13495 17663
rect 19257 17629 19291 17663
rect 19625 17629 19659 17663
rect 23949 17629 23983 17663
rect 24041 17629 24075 17663
rect 24777 17629 24811 17663
rect 24869 17629 24903 17663
rect 24961 17629 24995 17663
rect 25145 17629 25179 17663
rect 25973 17629 26007 17663
rect 26157 17629 26191 17663
rect 26617 17629 26651 17663
rect 26801 17629 26835 17663
rect 27077 17629 27111 17663
rect 27261 17629 27295 17663
rect 27905 17629 27939 17663
rect 28089 17629 28123 17663
rect 28181 17629 28215 17663
rect 28273 17629 28307 17663
rect 28457 17629 28491 17663
rect 28733 17629 28767 17663
rect 28917 17629 28951 17663
rect 29009 17629 29043 17663
rect 29101 17629 29135 17663
rect 30021 17629 30055 17663
rect 30205 17629 30239 17663
rect 30297 17629 30331 17663
rect 30389 17629 30423 17663
rect 30573 17629 30607 17663
rect 30849 17629 30883 17663
rect 31861 17629 31895 17663
rect 32045 17629 32079 17663
rect 32413 17629 32447 17663
rect 32814 17629 32848 17663
rect 33333 17629 33367 17663
rect 33701 17629 33735 17663
rect 34345 17629 34379 17663
rect 35449 17629 35483 17663
rect 3801 17561 3835 17595
rect 4997 17561 5031 17595
rect 7297 17561 7331 17595
rect 7389 17561 7423 17595
rect 9321 17561 9355 17595
rect 11161 17561 11195 17595
rect 14381 17561 14415 17595
rect 16957 17561 16991 17595
rect 19441 17561 19475 17595
rect 19533 17561 19567 17595
rect 21557 17561 21591 17595
rect 23121 17561 23155 17595
rect 24225 17561 24259 17595
rect 26433 17561 26467 17595
rect 26525 17561 26559 17595
rect 26985 17561 27019 17595
rect 32597 17561 32631 17595
rect 34529 17561 34563 17595
rect 4797 17493 4831 17527
rect 7113 17493 7147 17527
rect 13553 17493 13587 17527
rect 13921 17493 13955 17527
rect 28641 17493 28675 17527
rect 29285 17493 29319 17527
rect 30757 17493 30791 17527
rect 32689 17493 32723 17527
rect 32873 17493 32907 17527
rect 7665 17289 7699 17323
rect 10425 17289 10459 17323
rect 10885 17289 10919 17323
rect 11529 17289 11563 17323
rect 11989 17289 12023 17323
rect 13185 17289 13219 17323
rect 13829 17289 13863 17323
rect 15117 17289 15151 17323
rect 22017 17289 22051 17323
rect 22385 17289 22419 17323
rect 23673 17289 23707 17323
rect 25881 17289 25915 17323
rect 27721 17289 27755 17323
rect 32965 17289 32999 17323
rect 36369 17289 36403 17323
rect 2789 17221 2823 17255
rect 4445 17221 4479 17255
rect 9137 17221 9171 17255
rect 10793 17221 10827 17255
rect 14105 17221 14139 17255
rect 18797 17221 18831 17255
rect 18997 17221 19031 17255
rect 28733 17221 28767 17255
rect 30113 17221 30147 17255
rect 30573 17221 30607 17255
rect 32137 17221 32171 17255
rect 33793 17221 33827 17255
rect 34529 17221 34563 17255
rect 34897 17221 34931 17255
rect 33563 17187 33597 17221
rect 2237 17153 2271 17187
rect 2421 17153 2455 17187
rect 2513 17153 2547 17187
rect 2605 17153 2639 17187
rect 4077 17153 4111 17187
rect 4905 17153 4939 17187
rect 6837 17153 6871 17187
rect 9413 17153 9447 17187
rect 11897 17153 11931 17187
rect 12541 17153 12575 17187
rect 12725 17153 12759 17187
rect 13001 17153 13035 17187
rect 15025 17153 15059 17187
rect 15209 17153 15243 17187
rect 18429 17153 18463 17187
rect 19901 17153 19935 17187
rect 22477 17153 22511 17187
rect 23305 17153 23339 17187
rect 23949 17153 23983 17187
rect 24041 17153 24075 17187
rect 24225 17153 24259 17187
rect 24501 17153 24535 17187
rect 24777 17153 24811 17187
rect 24961 17153 24995 17187
rect 25237 17153 25271 17187
rect 25421 17153 25455 17187
rect 25605 17153 25639 17187
rect 25789 17153 25823 17187
rect 25973 17153 26007 17187
rect 26249 17153 26283 17187
rect 27261 17153 27295 17187
rect 27537 17153 27571 17187
rect 27721 17153 27755 17187
rect 28917 17153 28951 17187
rect 29101 17153 29135 17187
rect 29285 17153 29319 17187
rect 29469 17153 29503 17187
rect 29837 17153 29871 17187
rect 29930 17153 29964 17187
rect 30205 17153 30239 17187
rect 30302 17153 30336 17187
rect 30665 17153 30699 17187
rect 30941 17153 30975 17187
rect 31217 17153 31251 17187
rect 31953 17153 31987 17187
rect 32321 17153 32355 17187
rect 32597 17153 32631 17187
rect 32689 17153 32723 17187
rect 32873 17153 32907 17187
rect 33149 17153 33183 17187
rect 33977 17153 34011 17187
rect 34253 17153 34287 17187
rect 34345 17153 34379 17187
rect 3433 17085 3467 17119
rect 4813 17085 4847 17119
rect 5365 17085 5399 17119
rect 7573 17085 7607 17119
rect 9505 17085 9539 17119
rect 10977 17085 11011 17119
rect 12081 17085 12115 17119
rect 20177 17085 20211 17119
rect 20637 17085 20671 17119
rect 21189 17085 21223 17119
rect 22661 17085 22695 17119
rect 23673 17085 23707 17119
rect 25513 17085 25547 17119
rect 26985 17085 27019 17119
rect 29193 17085 29227 17119
rect 31033 17085 31067 17119
rect 32505 17085 32539 17119
rect 33333 17085 33367 17119
rect 34621 17085 34655 17119
rect 10149 17017 10183 17051
rect 19349 17017 19383 17051
rect 23397 17017 23431 17051
rect 23857 17017 23891 17051
rect 24593 17017 24627 17051
rect 27077 17017 27111 17051
rect 27445 17017 27479 17051
rect 30481 17017 30515 17051
rect 33425 17017 33459 17051
rect 34069 17017 34103 17051
rect 2421 16949 2455 16983
rect 2789 16949 2823 16983
rect 2881 16949 2915 16983
rect 4537 16949 4571 16983
rect 5089 16949 5123 16983
rect 5917 16949 5951 16983
rect 6745 16949 6779 16983
rect 6929 16949 6963 16983
rect 18613 16949 18647 16983
rect 18981 16949 19015 16983
rect 19165 16949 19199 16983
rect 19717 16949 19751 16983
rect 20085 16949 20119 16983
rect 24409 16949 24443 16983
rect 31401 16949 31435 16983
rect 31769 16949 31803 16983
rect 33609 16949 33643 16983
rect 3433 16745 3467 16779
rect 7021 16745 7055 16779
rect 12817 16745 12851 16779
rect 15117 16745 15151 16779
rect 16221 16745 16255 16779
rect 17496 16745 17530 16779
rect 18981 16745 19015 16779
rect 25145 16745 25179 16779
rect 29745 16745 29779 16779
rect 32229 16745 32263 16779
rect 34529 16745 34563 16779
rect 5181 16677 5215 16711
rect 10977 16677 11011 16711
rect 16129 16677 16163 16711
rect 24869 16677 24903 16711
rect 30941 16677 30975 16711
rect 32137 16677 32171 16711
rect 32505 16677 32539 16711
rect 1409 16609 1443 16643
rect 4261 16609 4295 16643
rect 6929 16609 6963 16643
rect 8493 16609 8527 16643
rect 9689 16609 9723 16643
rect 11253 16609 11287 16643
rect 15991 16609 16025 16643
rect 17233 16609 17267 16643
rect 19533 16609 19567 16643
rect 26801 16609 26835 16643
rect 27261 16609 27295 16643
rect 27537 16609 27571 16643
rect 30113 16609 30147 16643
rect 31033 16609 31067 16643
rect 31125 16609 31159 16643
rect 32321 16609 32355 16643
rect 33057 16609 33091 16643
rect 8769 16541 8803 16575
rect 10701 16541 10735 16575
rect 11345 16541 11379 16575
rect 13001 16541 13035 16575
rect 13277 16541 13311 16575
rect 13461 16541 13495 16575
rect 15301 16541 15335 16575
rect 15577 16541 15611 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 16313 16541 16347 16575
rect 19257 16541 19291 16575
rect 21097 16541 21131 16575
rect 22293 16541 22327 16575
rect 25145 16541 25179 16575
rect 25329 16541 25363 16575
rect 30021 16541 30055 16575
rect 30570 16541 30604 16575
rect 31309 16541 31343 16575
rect 31401 16541 31435 16575
rect 32045 16541 32079 16575
rect 32597 16541 32631 16575
rect 32781 16541 32815 16575
rect 1685 16473 1719 16507
rect 3249 16473 3283 16507
rect 3449 16473 3483 16507
rect 4997 16473 5031 16507
rect 6653 16473 6687 16507
rect 9965 16473 9999 16507
rect 22569 16473 22603 16507
rect 26065 16473 26099 16507
rect 27077 16473 27111 16507
rect 29285 16473 29319 16507
rect 31125 16473 31159 16507
rect 3157 16405 3191 16439
rect 3617 16405 3651 16439
rect 9137 16405 9171 16439
rect 9505 16405 9539 16439
rect 9597 16405 9631 16439
rect 11621 16405 11655 16439
rect 21005 16405 21039 16439
rect 21189 16405 21223 16439
rect 24041 16405 24075 16439
rect 30389 16405 30423 16439
rect 30573 16405 30607 16439
rect 2605 16201 2639 16235
rect 8309 16201 8343 16235
rect 10977 16201 11011 16235
rect 13645 16201 13679 16235
rect 15577 16201 15611 16235
rect 17325 16201 17359 16235
rect 18613 16201 18647 16235
rect 20085 16201 20119 16235
rect 20177 16201 20211 16235
rect 20571 16201 20605 16235
rect 23029 16201 23063 16235
rect 23397 16201 23431 16235
rect 26709 16201 26743 16235
rect 28089 16201 28123 16235
rect 28273 16201 28307 16235
rect 31907 16201 31941 16235
rect 2237 16133 2271 16167
rect 2697 16133 2731 16167
rect 9505 16133 9539 16167
rect 13185 16133 13219 16167
rect 15393 16133 15427 16167
rect 20361 16133 20395 16167
rect 23489 16133 23523 16167
rect 29101 16133 29135 16167
rect 2421 16065 2455 16099
rect 3341 16065 3375 16099
rect 3433 16065 3467 16099
rect 3525 16065 3559 16099
rect 5549 16065 5583 16099
rect 6561 16065 6595 16099
rect 8493 16065 8527 16099
rect 13461 16065 13495 16099
rect 13737 16065 13771 16099
rect 13921 16065 13955 16099
rect 14749 16065 14783 16099
rect 15301 16065 15335 16099
rect 15485 16065 15519 16099
rect 15761 16065 15795 16099
rect 16037 16065 16071 16099
rect 16221 16065 16255 16099
rect 16681 16065 16715 16099
rect 16865 16065 16899 16099
rect 17141 16065 17175 16099
rect 17969 16065 18003 16099
rect 18153 16065 18187 16099
rect 18245 16065 18279 16099
rect 18337 16065 18371 16099
rect 18705 16065 18739 16099
rect 19257 16065 19291 16099
rect 20269 16065 20303 16099
rect 20821 16065 20855 16099
rect 21005 16065 21039 16099
rect 21465 16065 21499 16099
rect 21557 16065 21591 16099
rect 24961 16065 24995 16099
rect 27537 16065 27571 16099
rect 28270 16065 28304 16099
rect 29377 16065 29411 16099
rect 29469 16065 29503 16099
rect 32505 16065 32539 16099
rect 33149 16065 33183 16099
rect 2329 15997 2363 16031
rect 3157 15997 3191 16031
rect 3801 15997 3835 16031
rect 5457 15997 5491 16031
rect 5917 15997 5951 16031
rect 6837 15997 6871 16031
rect 8677 15997 8711 16031
rect 9229 15997 9263 16031
rect 13369 15997 13403 16031
rect 14841 15997 14875 16031
rect 15025 15997 15059 16031
rect 19809 15997 19843 16031
rect 23581 15997 23615 16031
rect 25237 15997 25271 16031
rect 28733 15997 28767 16031
rect 29101 15997 29135 16031
rect 30113 15997 30147 16031
rect 30481 15997 30515 16031
rect 33977 15997 34011 16031
rect 3433 15929 3467 15963
rect 21189 15929 21223 15963
rect 28641 15929 28675 15963
rect 32781 15929 32815 15963
rect 5273 15861 5307 15895
rect 13185 15861 13219 15895
rect 13921 15861 13955 15895
rect 14381 15861 14415 15895
rect 20545 15861 20579 15895
rect 20729 15861 20763 15895
rect 21281 15861 21315 15895
rect 26985 15861 27019 15895
rect 29285 15861 29319 15895
rect 32873 15861 32907 15895
rect 2881 15657 2915 15691
rect 4169 15657 4203 15691
rect 5181 15657 5215 15691
rect 13277 15657 13311 15691
rect 15945 15657 15979 15691
rect 16497 15657 16531 15691
rect 17601 15657 17635 15691
rect 29561 15657 29595 15691
rect 12541 15589 12575 15623
rect 13645 15589 13679 15623
rect 16405 15589 16439 15623
rect 16681 15589 16715 15623
rect 25237 15589 25271 15623
rect 27813 15589 27847 15623
rect 3249 15521 3283 15555
rect 4445 15521 4479 15555
rect 14105 15521 14139 15555
rect 14381 15521 14415 15555
rect 15853 15521 15887 15555
rect 16037 15521 16071 15555
rect 22017 15521 22051 15555
rect 25697 15521 25731 15555
rect 25789 15521 25823 15555
rect 32597 15521 32631 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 3065 15453 3099 15487
rect 4353 15453 4387 15487
rect 4813 15453 4847 15487
rect 10057 15453 10091 15487
rect 10793 15453 10827 15487
rect 12633 15453 12667 15487
rect 12817 15453 12851 15487
rect 13093 15453 13127 15487
rect 13553 15453 13587 15487
rect 13737 15453 13771 15487
rect 13829 15453 13863 15487
rect 15945 15453 15979 15487
rect 16221 15453 16255 15487
rect 17785 15453 17819 15487
rect 17969 15453 18003 15487
rect 18245 15453 18279 15487
rect 18429 15453 18463 15487
rect 18981 15453 19015 15487
rect 19993 15453 20027 15487
rect 22293 15453 22327 15487
rect 22661 15453 22695 15487
rect 24961 15453 24995 15487
rect 25605 15453 25639 15487
rect 26985 15453 27019 15487
rect 29745 15453 29779 15487
rect 37289 15453 37323 15487
rect 4721 15385 4755 15419
rect 11069 15385 11103 15419
rect 13369 15385 13403 15419
rect 16957 15385 16991 15419
rect 18061 15385 18095 15419
rect 19257 15385 19291 15419
rect 28181 15385 28215 15419
rect 32873 15385 32907 15419
rect 35265 15385 35299 15419
rect 35449 15385 35483 15419
rect 2605 15317 2639 15351
rect 4629 15317 4663 15351
rect 20545 15317 20579 15351
rect 23673 15317 23707 15351
rect 24133 15317 24167 15351
rect 24409 15317 24443 15351
rect 27629 15317 27663 15351
rect 27721 15317 27755 15351
rect 31033 15317 31067 15351
rect 31585 15317 31619 15351
rect 34345 15317 34379 15351
rect 36645 15317 36679 15351
rect 38485 15317 38519 15351
rect 10977 15113 11011 15147
rect 11345 15113 11379 15147
rect 14473 15113 14507 15147
rect 14565 15113 14599 15147
rect 18521 15113 18555 15147
rect 19717 15113 19751 15147
rect 23949 15113 23983 15147
rect 28733 15113 28767 15147
rect 30113 15113 30147 15147
rect 4813 15045 4847 15079
rect 11529 15045 11563 15079
rect 18889 15045 18923 15079
rect 19901 15045 19935 15079
rect 20177 15045 20211 15079
rect 33149 15045 33183 15079
rect 1409 14977 1443 15011
rect 5089 14977 5123 15011
rect 5641 14977 5675 15011
rect 5917 14977 5951 15011
rect 6101 14977 6135 15011
rect 6653 14977 6687 15011
rect 8769 14977 8803 15011
rect 12725 14977 12759 15011
rect 17693 14977 17727 15011
rect 17785 14977 17819 15011
rect 18705 14977 18739 15011
rect 18797 14977 18831 15011
rect 19073 14977 19107 15011
rect 19441 14977 19475 15011
rect 19533 14977 19567 15011
rect 19809 14977 19843 15011
rect 19993 14977 20027 15011
rect 20085 14977 20119 15011
rect 20361 14977 20395 15011
rect 24041 14977 24075 15011
rect 24225 14977 24259 15011
rect 26249 14977 26283 15011
rect 26985 14977 27019 15011
rect 30389 14977 30423 15011
rect 30573 14977 30607 15011
rect 32873 14977 32907 15011
rect 36645 14977 36679 15011
rect 1685 14909 1719 14943
rect 3157 14909 3191 14943
rect 3893 14909 3927 14943
rect 4905 14909 4939 14943
rect 6929 14909 6963 14943
rect 8677 14909 8711 14943
rect 9045 14909 9079 14943
rect 10701 14909 10735 14943
rect 10885 14909 10919 14943
rect 12541 14909 12575 14943
rect 13001 14909 13035 14943
rect 15117 14909 15151 14943
rect 17601 14909 17635 14943
rect 22201 14909 22235 14943
rect 22477 14909 22511 14943
rect 24317 14909 24351 14943
rect 25973 14909 26007 14943
rect 27261 14909 27295 14943
rect 34805 14909 34839 14943
rect 35081 14909 35115 14943
rect 5273 14841 5307 14875
rect 5733 14841 5767 14875
rect 19257 14841 19291 14875
rect 36737 14841 36771 14875
rect 3249 14773 3283 14807
rect 4813 14773 4847 14807
rect 6009 14773 6043 14807
rect 10517 14773 10551 14807
rect 18429 14773 18463 14807
rect 20545 14773 20579 14807
rect 24133 14773 24167 14807
rect 24501 14773 24535 14807
rect 30757 14773 30791 14807
rect 34621 14773 34655 14807
rect 36553 14773 36587 14807
rect 2237 14569 2271 14603
rect 4537 14569 4571 14603
rect 5089 14569 5123 14603
rect 5181 14569 5215 14603
rect 9597 14569 9631 14603
rect 11437 14569 11471 14603
rect 17325 14569 17359 14603
rect 20085 14569 20119 14603
rect 23673 14569 23707 14603
rect 24133 14569 24167 14603
rect 25513 14569 25547 14603
rect 26801 14569 26835 14603
rect 33241 14569 33275 14603
rect 34805 14569 34839 14603
rect 35265 14569 35299 14603
rect 2145 14501 2179 14535
rect 4261 14501 4295 14535
rect 9045 14501 9079 14535
rect 13001 14501 13035 14535
rect 16405 14501 16439 14535
rect 24685 14501 24719 14535
rect 31309 14501 31343 14535
rect 34897 14501 34931 14535
rect 36645 14501 36679 14535
rect 2697 14433 2731 14467
rect 3617 14433 3651 14467
rect 4813 14433 4847 14467
rect 5365 14433 5399 14467
rect 5457 14433 5491 14467
rect 5641 14433 5675 14467
rect 10241 14433 10275 14467
rect 13645 14433 13679 14467
rect 18797 14433 18831 14467
rect 24869 14433 24903 14467
rect 25053 14433 25087 14467
rect 26893 14433 26927 14467
rect 27169 14433 27203 14467
rect 29561 14433 29595 14467
rect 31493 14433 31527 14467
rect 34713 14433 34747 14467
rect 37013 14433 37047 14467
rect 1869 14365 1903 14399
rect 2421 14365 2455 14399
rect 2605 14365 2639 14399
rect 3801 14365 3835 14399
rect 3985 14365 4019 14399
rect 4353 14365 4387 14399
rect 4905 14365 4939 14399
rect 5549 14365 5583 14399
rect 5917 14365 5951 14399
rect 10057 14365 10091 14399
rect 11069 14365 11103 14399
rect 13369 14365 13403 14399
rect 13921 14365 13955 14399
rect 16589 14365 16623 14399
rect 19073 14365 19107 14399
rect 19809 14365 19843 14399
rect 21833 14365 21867 14399
rect 22845 14365 22879 14399
rect 23857 14365 23891 14399
rect 23949 14365 23983 14399
rect 24225 14365 24259 14399
rect 24409 14365 24443 14399
rect 26525 14365 26559 14399
rect 29193 14365 29227 14399
rect 29377 14365 29411 14399
rect 34989 14365 35023 14399
rect 35081 14365 35115 14399
rect 35541 14365 35575 14399
rect 36369 14365 36403 14399
rect 36737 14365 36771 14399
rect 2145 14297 2179 14331
rect 2973 14297 3007 14331
rect 4445 14297 4479 14331
rect 6193 14297 6227 14331
rect 9965 14297 9999 14331
rect 12909 14297 12943 14331
rect 14197 14297 14231 14331
rect 15301 14297 15335 14331
rect 21557 14297 21591 14331
rect 23581 14297 23615 14331
rect 24685 14297 24719 14331
rect 25145 14297 25179 14331
rect 26801 14297 26835 14331
rect 29285 14297 29319 14331
rect 29837 14297 29871 14331
rect 31769 14297 31803 14331
rect 35449 14297 35483 14331
rect 36645 14297 36679 14331
rect 1961 14229 1995 14263
rect 3893 14229 3927 14263
rect 7665 14229 7699 14263
rect 10425 14229 10459 14263
rect 13461 14229 13495 14263
rect 15025 14229 15059 14263
rect 16773 14229 16807 14263
rect 19257 14229 19291 14263
rect 24501 14229 24535 14263
rect 26617 14229 26651 14263
rect 28641 14229 28675 14263
rect 36461 14229 36495 14263
rect 38485 14229 38519 14263
rect 3525 14025 3559 14059
rect 5365 14025 5399 14059
rect 6009 14025 6043 14059
rect 9873 14025 9907 14059
rect 12357 14025 12391 14059
rect 13737 14025 13771 14059
rect 17785 14025 17819 14059
rect 19717 14025 19751 14059
rect 20729 14025 20763 14059
rect 24501 14025 24535 14059
rect 25053 14025 25087 14059
rect 27077 14025 27111 14059
rect 27721 14025 27755 14059
rect 30297 14025 30331 14059
rect 31033 14025 31067 14059
rect 31217 14025 31251 14059
rect 32965 14025 32999 14059
rect 33701 14025 33735 14059
rect 35341 14025 35375 14059
rect 36001 14025 36035 14059
rect 36829 14025 36863 14059
rect 37565 14025 37599 14059
rect 3709 13957 3743 13991
rect 4981 13957 5015 13991
rect 5181 13957 5215 13991
rect 5641 13957 5675 13991
rect 5857 13957 5891 13991
rect 7481 13957 7515 13991
rect 11253 13957 11287 13991
rect 18245 13957 18279 13991
rect 19257 13957 19291 13991
rect 19457 13957 19491 13991
rect 20361 13957 20395 13991
rect 20577 13957 20611 13991
rect 20913 13957 20947 13991
rect 24685 13957 24719 13991
rect 29837 13957 29871 13991
rect 33149 13957 33183 13991
rect 33241 13957 33275 13991
rect 35541 13957 35575 13991
rect 35909 13957 35943 13991
rect 36277 13957 36311 13991
rect 1777 13889 1811 13923
rect 5273 13889 5307 13923
rect 5549 13889 5583 13923
rect 6377 13889 6411 13923
rect 7113 13889 7147 13923
rect 7297 13889 7331 13923
rect 8125 13889 8159 13923
rect 10333 13889 10367 13923
rect 10425 13889 10459 13923
rect 11161 13889 11195 13923
rect 11345 13889 11379 13923
rect 11713 13889 11747 13923
rect 11897 13889 11931 13923
rect 12173 13889 12207 13923
rect 12633 13889 12667 13923
rect 12909 13889 12943 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 13553 13889 13587 13923
rect 16957 13889 16991 13923
rect 17233 13889 17267 13923
rect 17877 13889 17911 13923
rect 18981 13889 19015 13923
rect 19165 13889 19199 13923
rect 19901 13889 19935 13923
rect 19993 13889 20027 13923
rect 20177 13889 20211 13923
rect 21005 13889 21039 13923
rect 21833 13889 21867 13923
rect 23765 13889 23799 13923
rect 24041 13889 24075 13923
rect 24133 13889 24167 13923
rect 24225 13889 24259 13923
rect 24409 13889 24443 13923
rect 24961 13889 24995 13923
rect 27353 13889 27387 13923
rect 28365 13889 28399 13923
rect 30021 13889 30055 13923
rect 30205 13889 30239 13923
rect 30573 13889 30607 13923
rect 31585 13889 31619 13923
rect 32873 13889 32907 13923
rect 33425 13889 33459 13923
rect 33517 13889 33551 13923
rect 34253 13889 34287 13923
rect 35725 13889 35759 13923
rect 36001 13889 36035 13923
rect 36093 13889 36127 13923
rect 37013 13889 37047 13923
rect 37105 13889 37139 13923
rect 38209 13889 38243 13923
rect 3985 13821 4019 13855
rect 6929 13821 6963 13855
rect 10609 13821 10643 13855
rect 12449 13821 12483 13855
rect 13461 13821 13495 13855
rect 15485 13821 15519 13855
rect 15761 13821 15795 13855
rect 16681 13821 16715 13855
rect 17969 13821 18003 13855
rect 18797 13821 18831 13855
rect 19073 13821 19107 13855
rect 22109 13821 22143 13855
rect 27077 13821 27111 13855
rect 30297 13821 30331 13855
rect 33241 13821 33275 13855
rect 36829 13821 36863 13855
rect 9965 13753 9999 13787
rect 13369 13753 13403 13787
rect 20085 13753 20119 13787
rect 23765 13753 23799 13787
rect 24685 13753 24719 13787
rect 27261 13753 27295 13787
rect 30665 13753 30699 13787
rect 2040 13685 2074 13719
rect 4813 13685 4847 13719
rect 4997 13685 5031 13719
rect 5549 13685 5583 13719
rect 5825 13685 5859 13719
rect 8388 13685 8422 13719
rect 14013 13685 14047 13719
rect 16773 13685 16807 13719
rect 16865 13685 16899 13719
rect 17141 13685 17175 13719
rect 17417 13685 17451 13719
rect 19441 13685 19475 13719
rect 19625 13685 19659 13719
rect 20545 13685 20579 13719
rect 23581 13685 23615 13719
rect 24869 13685 24903 13719
rect 30481 13685 30515 13719
rect 31033 13685 31067 13719
rect 31493 13685 31527 13719
rect 33149 13685 33183 13719
rect 35173 13685 35207 13719
rect 35357 13685 35391 13719
rect 3801 13481 3835 13515
rect 3985 13481 4019 13515
rect 6101 13481 6135 13515
rect 13001 13481 13035 13515
rect 13369 13481 13403 13515
rect 15301 13481 15335 13515
rect 17555 13481 17589 13515
rect 19349 13481 19383 13515
rect 20637 13481 20671 13515
rect 21925 13481 21959 13515
rect 22109 13481 22143 13515
rect 23489 13481 23523 13515
rect 25237 13481 25271 13515
rect 36461 13481 36495 13515
rect 7849 13413 7883 13447
rect 13645 13413 13679 13447
rect 21281 13413 21315 13447
rect 27813 13413 27847 13447
rect 2329 13345 2363 13379
rect 2789 13345 2823 13379
rect 3617 13345 3651 13379
rect 7941 13345 7975 13379
rect 9413 13345 9447 13379
rect 11805 13345 11839 13379
rect 12449 13345 12483 13379
rect 12817 13345 12851 13379
rect 14749 13345 14783 13379
rect 15761 13345 15795 13379
rect 16129 13345 16163 13379
rect 20269 13345 20303 13379
rect 21097 13345 21131 13379
rect 22661 13345 22695 13379
rect 23949 13345 23983 13379
rect 25605 13345 25639 13379
rect 28365 13345 28399 13379
rect 28457 13345 28491 13379
rect 30573 13345 30607 13379
rect 32505 13345 32539 13379
rect 34713 13345 34747 13379
rect 36737 13345 36771 13379
rect 2421 13277 2455 13311
rect 2973 13277 3007 13311
rect 4353 13277 4387 13311
rect 7389 13277 7423 13311
rect 7573 13277 7607 13311
rect 8493 13277 8527 13311
rect 9505 13277 9539 13311
rect 12265 13277 12299 13311
rect 13001 13277 13035 13311
rect 13553 13277 13587 13311
rect 13737 13277 13771 13311
rect 13829 13277 13863 13311
rect 14933 13277 14967 13311
rect 18521 13277 18555 13311
rect 19533 13277 19567 13311
rect 20085 13277 20119 13311
rect 21373 13277 21407 13311
rect 22569 13277 22603 13311
rect 23305 13277 23339 13311
rect 23581 13277 23615 13311
rect 23857 13277 23891 13311
rect 24593 13277 24627 13311
rect 24869 13277 24903 13311
rect 25053 13277 25087 13311
rect 25145 13277 25179 13311
rect 25421 13277 25455 13311
rect 26525 13277 26559 13311
rect 26801 13277 26835 13311
rect 28549 13277 28583 13311
rect 28641 13277 28675 13311
rect 4169 13209 4203 13243
rect 4629 13209 4663 13243
rect 7849 13209 7883 13243
rect 11529 13209 11563 13243
rect 12725 13209 12759 13243
rect 20913 13209 20947 13243
rect 22477 13209 22511 13243
rect 24409 13209 24443 13243
rect 26709 13209 26743 13243
rect 27629 13209 27663 13243
rect 29653 13209 29687 13243
rect 29929 13209 29963 13243
rect 30849 13209 30883 13243
rect 32781 13209 32815 13243
rect 34529 13209 34563 13243
rect 34989 13209 35023 13243
rect 37013 13209 37047 13243
rect 3969 13141 4003 13175
rect 7297 13141 7331 13175
rect 7665 13141 7699 13175
rect 9597 13141 9631 13175
rect 9965 13141 9999 13175
rect 10057 13141 10091 13175
rect 11897 13141 11931 13175
rect 12357 13141 12391 13175
rect 13185 13141 13219 13175
rect 14841 13141 14875 13175
rect 18705 13141 18739 13175
rect 19901 13141 19935 13175
rect 21097 13141 21131 13175
rect 23121 13141 23155 13175
rect 24225 13141 24259 13175
rect 26801 13141 26835 13175
rect 28181 13141 28215 13175
rect 29745 13141 29779 13175
rect 32321 13141 32355 13175
rect 38485 13141 38519 13175
rect 4261 12937 4295 12971
rect 4813 12937 4847 12971
rect 4997 12937 5031 12971
rect 11161 12937 11195 12971
rect 12173 12937 12207 12971
rect 12633 12937 12667 12971
rect 18797 12937 18831 12971
rect 21557 12937 21591 12971
rect 28825 12937 28859 12971
rect 30665 12937 30699 12971
rect 31125 12937 31159 12971
rect 35725 12937 35759 12971
rect 36461 12937 36495 12971
rect 37013 12937 37047 12971
rect 2789 12869 2823 12903
rect 6929 12869 6963 12903
rect 9689 12869 9723 12903
rect 17325 12869 17359 12903
rect 26433 12869 26467 12903
rect 33057 12869 33091 12903
rect 37289 12869 37323 12903
rect 4537 12801 4571 12835
rect 4721 12801 4755 12835
rect 4905 12801 4939 12835
rect 6653 12801 6687 12835
rect 9413 12801 9447 12835
rect 11529 12801 11563 12835
rect 12817 12801 12851 12835
rect 13093 12801 13127 12835
rect 13277 12801 13311 12835
rect 15945 12801 15979 12835
rect 17049 12801 17083 12835
rect 19533 12801 19567 12835
rect 19717 12801 19751 12835
rect 19901 12801 19935 12835
rect 20085 12801 20119 12835
rect 23765 12801 23799 12835
rect 24041 12801 24075 12835
rect 24225 12801 24259 12835
rect 26341 12801 26375 12835
rect 26617 12801 26651 12835
rect 30573 12801 30607 12835
rect 30849 12801 30883 12835
rect 31401 12801 31435 12835
rect 31493 12801 31527 12835
rect 31585 12801 31619 12835
rect 31769 12801 31803 12835
rect 36001 12801 36035 12835
rect 36093 12801 36127 12835
rect 36185 12801 36219 12835
rect 36645 12801 36679 12835
rect 36921 12801 36955 12835
rect 37105 12801 37139 12835
rect 37565 12801 37599 12835
rect 2513 12733 2547 12767
rect 4353 12733 4387 12767
rect 9229 12733 9263 12767
rect 14105 12733 14139 12767
rect 14197 12733 14231 12767
rect 15669 12733 15703 12767
rect 19809 12733 19843 12767
rect 20177 12733 20211 12767
rect 20729 12733 20763 12767
rect 20913 12733 20947 12767
rect 26985 12733 27019 12767
rect 27261 12733 27295 12767
rect 30297 12733 30331 12767
rect 31033 12733 31067 12767
rect 35909 12733 35943 12767
rect 36829 12733 36863 12767
rect 37289 12733 37323 12767
rect 8401 12665 8435 12699
rect 20085 12665 20119 12699
rect 32689 12665 32723 12699
rect 8677 12597 8711 12631
rect 13461 12597 13495 12631
rect 19349 12597 19383 12631
rect 23581 12597 23615 12631
rect 26801 12597 26835 12631
rect 28733 12597 28767 12631
rect 33057 12597 33091 12631
rect 33241 12597 33275 12631
rect 37473 12597 37507 12631
rect 4813 12393 4847 12427
rect 9229 12393 9263 12427
rect 10149 12393 10183 12427
rect 13185 12393 13219 12427
rect 14105 12393 14139 12427
rect 14565 12393 14599 12427
rect 15393 12393 15427 12427
rect 21097 12393 21131 12427
rect 24869 12393 24903 12427
rect 26801 12393 26835 12427
rect 26985 12393 27019 12427
rect 28365 12393 28399 12427
rect 29377 12393 29411 12427
rect 31033 12393 31067 12427
rect 31309 12393 31343 12427
rect 32505 12393 32539 12427
rect 36645 12393 36679 12427
rect 5825 12325 5859 12359
rect 23029 12325 23063 12359
rect 25053 12325 25087 12359
rect 28181 12325 28215 12359
rect 28825 12325 28859 12359
rect 29837 12325 29871 12359
rect 31585 12325 31619 12359
rect 32689 12325 32723 12359
rect 34897 12325 34931 12359
rect 7941 12257 7975 12291
rect 12541 12257 12575 12291
rect 12633 12257 12667 12291
rect 14197 12257 14231 12291
rect 14841 12257 14875 12291
rect 14933 12257 14967 12291
rect 15761 12257 15795 12291
rect 18245 12257 18279 12291
rect 19625 12257 19659 12291
rect 22293 12257 22327 12291
rect 23121 12257 23155 12291
rect 23213 12257 23247 12291
rect 25421 12257 25455 12291
rect 32781 12257 32815 12291
rect 33057 12257 33091 12291
rect 3617 12189 3651 12223
rect 5089 12189 5123 12223
rect 6101 12189 6135 12223
rect 6193 12189 6227 12223
rect 8585 12189 8619 12223
rect 8769 12189 8803 12223
rect 9781 12189 9815 12223
rect 13369 12189 13403 12223
rect 13645 12189 13679 12223
rect 13829 12189 13863 12223
rect 14105 12189 14139 12223
rect 14381 12189 14415 12223
rect 17509 12189 17543 12223
rect 17969 12189 18003 12223
rect 18889 12189 18923 12223
rect 19349 12189 19383 12223
rect 22201 12189 22235 12223
rect 22937 12189 22971 12223
rect 23397 12189 23431 12223
rect 23673 12189 23707 12223
rect 23949 12189 23983 12223
rect 24041 12189 24075 12223
rect 24409 12189 24443 12223
rect 24685 12189 24719 12223
rect 25513 12189 25547 12223
rect 28733 12189 28767 12223
rect 29009 12189 29043 12223
rect 29653 12189 29687 12223
rect 30389 12189 30423 12223
rect 30573 12189 30607 12223
rect 30757 12189 30791 12223
rect 30849 12189 30883 12223
rect 31585 12189 31619 12223
rect 31769 12189 31803 12223
rect 35081 12189 35115 12223
rect 36277 12189 36311 12223
rect 36645 12189 36679 12223
rect 36737 12189 36771 12223
rect 4169 12121 4203 12155
rect 4797 12121 4831 12155
rect 4997 12121 5031 12155
rect 5733 12121 5767 12155
rect 5825 12121 5859 12155
rect 6469 12121 6503 12155
rect 8125 12121 8159 12155
rect 10117 12121 10151 12155
rect 10333 12121 10367 12155
rect 11805 12121 11839 12155
rect 17233 12121 17267 12155
rect 24133 12121 24167 12155
rect 26617 12121 26651 12155
rect 26817 12121 26851 12155
rect 29193 12121 29227 12155
rect 31125 12121 31159 12155
rect 31325 12121 31359 12155
rect 32321 12121 32355 12155
rect 36921 12121 36955 12155
rect 3893 12053 3927 12087
rect 4353 12053 4387 12087
rect 4629 12053 4663 12087
rect 6009 12053 6043 12087
rect 8217 12053 8251 12087
rect 8677 12053 8711 12087
rect 9965 12053 9999 12087
rect 11621 12053 11655 12087
rect 11897 12053 11931 12087
rect 12725 12053 12759 12087
rect 13093 12053 13127 12087
rect 15025 12053 15059 12087
rect 17601 12053 17635 12087
rect 18061 12053 18095 12087
rect 18981 12053 19015 12087
rect 21833 12053 21867 12087
rect 22753 12053 22787 12087
rect 23765 12053 23799 12087
rect 24501 12053 24535 12087
rect 24961 12053 24995 12087
rect 25697 12053 25731 12087
rect 28365 12053 28399 12087
rect 29101 12053 29135 12087
rect 30481 12053 30515 12087
rect 31493 12053 31527 12087
rect 32521 12053 32555 12087
rect 34529 12053 34563 12087
rect 35725 12053 35759 12087
rect 36461 12053 36495 12087
rect 4445 11849 4479 11883
rect 9597 11849 9631 11883
rect 10885 11849 10919 11883
rect 18429 11849 18463 11883
rect 20361 11849 20395 11883
rect 23029 11849 23063 11883
rect 33241 11849 33275 11883
rect 35081 11849 35115 11883
rect 6377 11781 6411 11815
rect 7389 11781 7423 11815
rect 8125 11781 8159 11815
rect 11161 11781 11195 11815
rect 13277 11781 13311 11815
rect 27077 11781 27111 11815
rect 37473 11781 37507 11815
rect 2973 11713 3007 11747
rect 3249 11713 3283 11747
rect 4077 11713 4111 11747
rect 13645 11713 13679 11747
rect 13829 11713 13863 11747
rect 16221 11713 16255 11747
rect 20453 11713 20487 11747
rect 22017 11713 22051 11747
rect 22569 11713 22603 11747
rect 23581 11713 23615 11747
rect 23765 11713 23799 11747
rect 24685 11713 24719 11747
rect 24869 11713 24903 11747
rect 25973 11713 26007 11747
rect 26157 11713 26191 11747
rect 26249 11713 26283 11747
rect 26525 11713 26559 11747
rect 26985 11713 27019 11747
rect 27261 11713 27295 11747
rect 30849 11713 30883 11747
rect 33057 11713 33091 11747
rect 35265 11713 35299 11747
rect 35449 11713 35483 11747
rect 35541 11713 35575 11747
rect 35725 11713 35759 11747
rect 35817 11713 35851 11747
rect 4353 11645 4387 11679
rect 5917 11645 5951 11679
rect 6193 11645 6227 11679
rect 7205 11645 7239 11679
rect 7849 11645 7883 11679
rect 11805 11645 11839 11679
rect 13553 11645 13587 11679
rect 16681 11645 16715 11679
rect 16957 11645 16991 11679
rect 18613 11645 18647 11679
rect 18889 11645 18923 11679
rect 22109 11645 22143 11679
rect 26341 11645 26375 11679
rect 26709 11645 26743 11679
rect 30941 11645 30975 11679
rect 32781 11645 32815 11679
rect 32873 11645 32907 11679
rect 32965 11645 32999 11679
rect 36645 11645 36679 11679
rect 3433 11577 3467 11611
rect 13829 11577 13863 11611
rect 22937 11577 22971 11611
rect 31217 11577 31251 11611
rect 35357 11577 35391 11611
rect 37841 11577 37875 11611
rect 2881 11509 2915 11543
rect 11253 11509 11287 11543
rect 11621 11509 11655 11543
rect 20637 11509 20671 11543
rect 22293 11509 22327 11543
rect 23581 11509 23615 11543
rect 24869 11509 24903 11543
rect 27445 11509 27479 11543
rect 37289 11509 37323 11543
rect 37473 11509 37507 11543
rect 2881 11305 2915 11339
rect 5549 11305 5583 11339
rect 6929 11305 6963 11339
rect 12265 11305 12299 11339
rect 17417 11305 17451 11339
rect 18337 11305 18371 11339
rect 21649 11305 21683 11339
rect 22017 11305 22051 11339
rect 22293 11305 22327 11339
rect 25973 11305 26007 11339
rect 28549 11305 28583 11339
rect 32781 11305 32815 11339
rect 33333 11305 33367 11339
rect 36093 11305 36127 11339
rect 36185 11305 36219 11339
rect 36277 11305 36311 11339
rect 12357 11237 12391 11271
rect 27629 11237 27663 11271
rect 28365 11237 28399 11271
rect 28641 11237 28675 11271
rect 2605 11169 2639 11203
rect 2973 11169 3007 11203
rect 3617 11169 3651 11203
rect 4077 11169 4111 11203
rect 5825 11169 5859 11203
rect 6561 11169 6595 11203
rect 7389 11169 7423 11203
rect 8217 11169 8251 11203
rect 10793 11169 10827 11203
rect 12817 11169 12851 11203
rect 13001 11169 13035 11203
rect 15853 11169 15887 11203
rect 17141 11169 17175 11203
rect 17969 11169 18003 11203
rect 28273 11169 28307 11203
rect 28549 11169 28583 11203
rect 29929 11169 29963 11203
rect 35173 11169 35207 11203
rect 36921 11169 36955 11203
rect 38393 11169 38427 11203
rect 1409 11101 1443 11135
rect 1685 11101 1719 11135
rect 2513 11101 2547 11135
rect 3801 11101 3835 11135
rect 6377 11101 6411 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 7297 11101 7331 11135
rect 7665 11101 7699 11135
rect 8401 11101 8435 11135
rect 8585 11101 8619 11135
rect 10517 11101 10551 11135
rect 12725 11101 12759 11135
rect 14105 11101 14139 11135
rect 18613 11101 18647 11135
rect 18797 11101 18831 11135
rect 21281 11101 21315 11135
rect 21465 11101 21499 11135
rect 21833 11101 21867 11135
rect 24409 11101 24443 11135
rect 24593 11101 24627 11135
rect 24869 11101 24903 11135
rect 26157 11101 26191 11135
rect 26249 11101 26283 11135
rect 26433 11101 26467 11135
rect 26525 11101 26559 11135
rect 27813 11101 27847 11135
rect 27905 11101 27939 11135
rect 28181 11101 28215 11135
rect 28733 11101 28767 11135
rect 29009 11101 29043 11135
rect 30021 11101 30055 11135
rect 30113 11101 30147 11135
rect 30205 11101 30239 11135
rect 30481 11101 30515 11135
rect 30665 11101 30699 11135
rect 32873 11101 32907 11135
rect 32965 11101 32999 11135
rect 33057 11101 33091 11135
rect 33241 11101 33275 11135
rect 33333 11101 33367 11135
rect 35357 11101 35391 11135
rect 35449 11101 35483 11135
rect 35633 11101 35667 11135
rect 35725 11101 35759 11135
rect 35817 11101 35851 11135
rect 36001 11101 36035 11135
rect 36645 11101 36679 11135
rect 14381 11033 14415 11067
rect 16313 11033 16347 11067
rect 16405 11033 16439 11067
rect 20913 11033 20947 11067
rect 24777 11033 24811 11067
rect 29193 11033 29227 11067
rect 1593 10965 1627 10999
rect 8493 10965 8527 10999
rect 17785 10965 17819 10999
rect 17877 10965 17911 10999
rect 29377 10965 29411 10999
rect 30389 10965 30423 10999
rect 30849 10965 30883 10999
rect 32597 10965 32631 10999
rect 33517 10965 33551 10999
rect 36277 10965 36311 10999
rect 1593 10761 1627 10795
rect 4445 10761 4479 10795
rect 10885 10761 10919 10795
rect 13369 10761 13403 10795
rect 14381 10761 14415 10795
rect 14841 10761 14875 10795
rect 22293 10761 22327 10795
rect 23029 10761 23063 10795
rect 24961 10761 24995 10795
rect 29193 10761 29227 10795
rect 34069 10761 34103 10795
rect 34437 10761 34471 10795
rect 34897 10761 34931 10795
rect 36645 10761 36679 10795
rect 2789 10693 2823 10727
rect 6837 10693 6871 10727
rect 12633 10693 12667 10727
rect 23857 10693 23891 10727
rect 24593 10693 24627 10727
rect 25605 10693 25639 10727
rect 27813 10693 27847 10727
rect 36905 10693 36939 10727
rect 37105 10693 37139 10727
rect 37473 10693 37507 10727
rect 37841 10693 37875 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 1869 10625 1903 10659
rect 2513 10625 2547 10659
rect 5089 10625 5123 10659
rect 6561 10625 6595 10659
rect 8585 10625 8619 10659
rect 9045 10625 9079 10659
rect 11069 10625 11103 10659
rect 13553 10625 13587 10659
rect 13829 10625 13863 10659
rect 14013 10625 14047 10659
rect 14749 10625 14783 10659
rect 17141 10625 17175 10659
rect 17785 10625 17819 10659
rect 22201 10625 22235 10659
rect 22661 10625 22695 10659
rect 22937 10625 22971 10659
rect 23121 10625 23155 10659
rect 23213 10625 23247 10659
rect 23397 10625 23431 10659
rect 24225 10625 24259 10659
rect 24317 10625 24351 10659
rect 24777 10625 24811 10659
rect 25789 10625 25823 10659
rect 26341 10625 26375 10659
rect 26433 10625 26467 10659
rect 26617 10625 26651 10659
rect 27169 10625 27203 10659
rect 27629 10625 27663 10659
rect 29009 10625 29043 10659
rect 29285 10625 29319 10659
rect 29469 10625 29503 10659
rect 30205 10625 30239 10659
rect 30481 10625 30515 10659
rect 30665 10625 30699 10659
rect 30757 10625 30791 10659
rect 30849 10625 30883 10659
rect 31033 10625 31067 10659
rect 32413 10625 32447 10659
rect 33057 10625 33091 10659
rect 33333 10625 33367 10659
rect 33517 10625 33551 10659
rect 33609 10625 33643 10659
rect 33885 10625 33919 10659
rect 34529 10625 34563 10659
rect 34621 10625 34655 10659
rect 36369 10625 36403 10659
rect 36461 10625 36495 10659
rect 37289 10625 37323 10659
rect 37565 10625 37599 10659
rect 2053 10557 2087 10591
rect 2237 10557 2271 10591
rect 4261 10557 4295 10591
rect 8401 10557 8435 10591
rect 9321 10557 9355 10591
rect 10793 10557 10827 10591
rect 12081 10557 12115 10591
rect 15025 10557 15059 10591
rect 18061 10557 18095 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 22477 10557 22511 10591
rect 23305 10557 23339 10591
rect 23949 10557 23983 10591
rect 25973 10557 26007 10591
rect 26801 10557 26835 10591
rect 27077 10557 27111 10591
rect 28825 10557 28859 10591
rect 29377 10557 29411 10591
rect 30021 10557 30055 10591
rect 32505 10557 32539 10591
rect 34161 10557 34195 10591
rect 36185 10557 36219 10591
rect 36277 10557 36311 10591
rect 38393 10557 38427 10591
rect 11529 10489 11563 10523
rect 22753 10489 22787 10523
rect 27537 10489 27571 10523
rect 33701 10489 33735 10523
rect 36737 10489 36771 10523
rect 8309 10421 8343 10455
rect 8769 10421 8803 10455
rect 11253 10421 11287 10455
rect 12909 10421 12943 10455
rect 17233 10421 17267 10455
rect 19533 10421 19567 10455
rect 21465 10421 21499 10455
rect 21833 10421 21867 10455
rect 24501 10421 24535 10455
rect 27997 10421 28031 10455
rect 30389 10421 30423 10455
rect 31217 10421 31251 10455
rect 32781 10421 32815 10455
rect 32873 10421 32907 10455
rect 34253 10421 34287 10455
rect 36921 10421 36955 10455
rect 37289 10421 37323 10455
rect 1685 10217 1719 10251
rect 8125 10217 8159 10251
rect 8769 10217 8803 10251
rect 14105 10217 14139 10251
rect 14841 10217 14875 10251
rect 16957 10217 16991 10251
rect 17601 10217 17635 10251
rect 18153 10217 18187 10251
rect 20729 10217 20763 10251
rect 23305 10217 23339 10251
rect 23673 10217 23707 10251
rect 24041 10217 24075 10251
rect 26341 10217 26375 10251
rect 28089 10217 28123 10251
rect 28825 10217 28859 10251
rect 30113 10217 30147 10251
rect 30757 10217 30791 10251
rect 34345 10217 34379 10251
rect 36461 10217 36495 10251
rect 15117 10149 15151 10183
rect 17693 10149 17727 10183
rect 25237 10149 25271 10183
rect 27905 10149 27939 10183
rect 28641 10149 28675 10183
rect 31769 10149 31803 10183
rect 4997 10081 5031 10115
rect 8493 10081 8527 10115
rect 9505 10081 9539 10115
rect 10517 10081 10551 10115
rect 11345 10081 11379 10115
rect 13737 10081 13771 10115
rect 15209 10081 15243 10115
rect 16405 10081 16439 10115
rect 17049 10081 17083 10115
rect 18705 10081 18739 10115
rect 21189 10081 21223 10115
rect 21373 10081 21407 10115
rect 22109 10081 22143 10115
rect 22753 10081 22787 10115
rect 23121 10081 23155 10115
rect 24685 10081 24719 10115
rect 24777 10081 24811 10115
rect 25697 10081 25731 10115
rect 26157 10081 26191 10115
rect 29653 10081 29687 10115
rect 31125 10081 31159 10115
rect 34713 10081 34747 10115
rect 36921 10081 36955 10115
rect 7389 10013 7423 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 8401 10013 8435 10047
rect 10701 10013 10735 10047
rect 14289 10013 14323 10047
rect 14565 10013 14599 10047
rect 14749 10013 14783 10047
rect 15025 10013 15059 10047
rect 15301 10013 15335 10047
rect 16313 10013 16347 10047
rect 16497 10013 16531 10047
rect 16773 10013 16807 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 17693 10013 17727 10047
rect 17877 10013 17911 10047
rect 17969 10013 18003 10047
rect 18521 10013 18555 10047
rect 21097 10013 21131 10047
rect 22569 10013 22603 10047
rect 22937 10013 22971 10047
rect 23305 10013 23339 10047
rect 23397 10013 23431 10047
rect 23581 10013 23615 10047
rect 23673 10013 23707 10047
rect 23851 10013 23885 10047
rect 23949 10013 23983 10047
rect 24133 10013 24167 10047
rect 24409 10013 24443 10047
rect 24593 10013 24627 10047
rect 24961 10013 24995 10047
rect 25605 10013 25639 10047
rect 26065 10013 26099 10047
rect 28273 10013 28307 10047
rect 28733 10013 28767 10047
rect 28917 10013 28951 10047
rect 29745 10013 29779 10047
rect 30297 10013 30331 10047
rect 30481 10013 30515 10047
rect 30757 10013 30791 10047
rect 30935 10013 30969 10047
rect 31585 10013 31619 10047
rect 31861 10013 31895 10047
rect 32137 10013 32171 10047
rect 33977 10013 34011 10047
rect 36645 10013 36679 10047
rect 5273 9945 5307 9979
rect 8953 9945 8987 9979
rect 11621 9945 11655 9979
rect 13645 9945 13679 9979
rect 17601 9945 17635 9979
rect 18613 9945 18647 9979
rect 22385 9945 22419 9979
rect 27629 9945 27663 9979
rect 28457 9945 28491 9979
rect 30389 9945 30423 9979
rect 31263 9945 31297 9979
rect 31401 9945 31435 9979
rect 31493 9945 31527 9979
rect 34989 9945 35023 9979
rect 1409 9877 1443 9911
rect 6745 9877 6779 9911
rect 6837 9877 6871 9911
rect 9873 9877 9907 9911
rect 11253 9877 11287 9911
rect 13093 9877 13127 9911
rect 13185 9877 13219 9911
rect 13553 9877 13587 9911
rect 16589 9877 16623 9911
rect 17141 9877 17175 9911
rect 21557 9877 21591 9911
rect 21925 9877 21959 9911
rect 22017 9877 22051 9911
rect 23029 9877 23063 9911
rect 23581 9877 23615 9911
rect 25145 9877 25179 9911
rect 31953 9877 31987 9911
rect 32321 9877 32355 9911
rect 34345 9877 34379 9911
rect 34529 9877 34563 9911
rect 38393 9877 38427 9911
rect 11069 9673 11103 9707
rect 11989 9673 12023 9707
rect 12449 9673 12483 9707
rect 13645 9673 13679 9707
rect 15393 9673 15427 9707
rect 23857 9673 23891 9707
rect 28181 9673 28215 9707
rect 29469 9673 29503 9707
rect 31309 9673 31343 9707
rect 31677 9673 31711 9707
rect 34437 9673 34471 9707
rect 36277 9673 36311 9707
rect 7573 9605 7607 9639
rect 7849 9605 7883 9639
rect 11253 9605 11287 9639
rect 12357 9605 12391 9639
rect 14013 9605 14047 9639
rect 21281 9605 21315 9639
rect 22201 9605 22235 9639
rect 25697 9605 25731 9639
rect 25881 9605 25915 9639
rect 26065 9605 26099 9639
rect 32873 9605 32907 9639
rect 35449 9605 35483 9639
rect 35909 9605 35943 9639
rect 36125 9605 36159 9639
rect 36369 9605 36403 9639
rect 37105 9605 37139 9639
rect 35219 9571 35253 9605
rect 4905 9537 4939 9571
rect 7389 9537 7423 9571
rect 7665 9537 7699 9571
rect 10977 9537 11011 9571
rect 13553 9537 13587 9571
rect 14749 9537 14783 9571
rect 15025 9537 15059 9571
rect 15577 9537 15611 9571
rect 15761 9537 15795 9571
rect 15853 9537 15887 9571
rect 16037 9537 16071 9571
rect 16405 9537 16439 9571
rect 16865 9537 16899 9571
rect 17141 9537 17175 9571
rect 17325 9537 17359 9571
rect 17601 9537 17635 9571
rect 22385 9537 22419 9571
rect 22477 9537 22511 9571
rect 22753 9537 22787 9571
rect 23121 9537 23155 9571
rect 23213 9537 23247 9571
rect 23305 9537 23339 9571
rect 23673 9537 23707 9571
rect 23857 9537 23891 9571
rect 25053 9537 25087 9571
rect 25973 9537 26007 9571
rect 26157 9537 26191 9571
rect 28089 9537 28123 9571
rect 28273 9537 28307 9571
rect 29285 9537 29319 9571
rect 29469 9537 29503 9571
rect 29561 9537 29595 9571
rect 29745 9537 29779 9571
rect 30941 9537 30975 9571
rect 31401 9537 31435 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 32413 9537 32447 9571
rect 32689 9537 32723 9571
rect 32965 9537 32999 9571
rect 33057 9537 33091 9571
rect 33241 9537 33275 9571
rect 34713 9537 34747 9571
rect 34897 9537 34931 9571
rect 35541 9537 35575 9571
rect 36553 9537 36587 9571
rect 36829 9537 36863 9571
rect 36921 9537 36955 9571
rect 4813 9469 4847 9503
rect 5273 9469 5307 9503
rect 8401 9469 8435 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 12633 9469 12667 9503
rect 13737 9469 13771 9503
rect 14565 9469 14599 9503
rect 14841 9469 14875 9503
rect 16129 9469 16163 9503
rect 17877 9469 17911 9503
rect 19441 9469 19475 9503
rect 19809 9469 19843 9503
rect 22845 9469 22879 9503
rect 23029 9469 23063 9503
rect 25513 9469 25547 9503
rect 29653 9469 29687 9503
rect 31033 9469 31067 9503
rect 31677 9469 31711 9503
rect 32505 9469 32539 9503
rect 34621 9469 34655 9503
rect 34805 9469 34839 9503
rect 35633 9469 35667 9503
rect 35817 9469 35851 9503
rect 36737 9469 36771 9503
rect 37105 9469 37139 9503
rect 11253 9401 11287 9435
rect 15209 9401 15243 9435
rect 15669 9401 15703 9435
rect 19349 9401 19383 9435
rect 31493 9401 31527 9435
rect 7205 9333 7239 9367
rect 10885 9333 10919 9367
rect 13185 9333 13219 9367
rect 15025 9333 15059 9367
rect 16221 9333 16255 9367
rect 16313 9333 16347 9367
rect 16681 9333 16715 9367
rect 22661 9333 22695 9367
rect 25145 9333 25179 9367
rect 30941 9333 30975 9367
rect 33425 9333 33459 9367
rect 35081 9333 35115 9367
rect 35265 9333 35299 9367
rect 35725 9333 35759 9367
rect 36093 9333 36127 9367
rect 8125 9129 8159 9163
rect 9689 9129 9723 9163
rect 10241 9129 10275 9163
rect 15025 9129 15059 9163
rect 16405 9129 16439 9163
rect 16773 9129 16807 9163
rect 16957 9129 16991 9163
rect 17969 9129 18003 9163
rect 26249 9129 26283 9163
rect 28181 9129 28215 9163
rect 28365 9129 28399 9163
rect 30021 9129 30055 9163
rect 30941 9129 30975 9163
rect 31861 9129 31895 9163
rect 38393 9129 38427 9163
rect 14289 9061 14323 9095
rect 21649 9061 21683 9095
rect 25881 9061 25915 9095
rect 30389 9061 30423 9095
rect 6653 8993 6687 9027
rect 11897 8993 11931 9027
rect 13369 8993 13403 9027
rect 18613 8993 18647 9027
rect 29929 8993 29963 9027
rect 30573 8993 30607 9027
rect 34805 8993 34839 9027
rect 35081 8993 35115 9027
rect 36645 8993 36679 9027
rect 6377 8925 6411 8959
rect 8677 8925 8711 8959
rect 9689 8925 9723 8959
rect 9873 8925 9907 8959
rect 9965 8925 9999 8959
rect 11621 8925 11655 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 14933 8925 14967 8959
rect 15209 8925 15243 8959
rect 15301 8925 15335 8959
rect 16129 8925 16163 8959
rect 16497 8925 16531 8959
rect 16589 8925 16623 8959
rect 16865 8925 16899 8959
rect 18337 8925 18371 8959
rect 21925 8925 21959 8959
rect 25053 8925 25087 8959
rect 25237 8925 25271 8959
rect 25329 8925 25363 8959
rect 26157 8925 26191 8959
rect 26249 8925 26283 8959
rect 26433 8925 26467 8959
rect 27813 8925 27847 8959
rect 28273 8925 28307 8959
rect 28457 8925 28491 8959
rect 29653 8925 29687 8959
rect 29745 8925 29779 8959
rect 30021 8925 30055 8959
rect 30113 8925 30147 8959
rect 30757 8925 30791 8959
rect 31677 8925 31711 8959
rect 31861 8925 31895 8959
rect 34897 8925 34931 8959
rect 34989 8925 35023 8959
rect 36461 8925 36495 8959
rect 8309 8857 8343 8891
rect 10425 8857 10459 8891
rect 15025 8857 15059 8891
rect 16313 8857 16347 8891
rect 21649 8857 21683 8891
rect 25881 8857 25915 8891
rect 26065 8857 26099 8891
rect 27997 8857 28031 8891
rect 29929 8857 29963 8891
rect 36921 8857 36955 8891
rect 10241 8789 10275 8823
rect 14841 8789 14875 8823
rect 15577 8789 15611 8823
rect 18429 8789 18463 8823
rect 21833 8789 21867 8823
rect 25237 8789 25271 8823
rect 25513 8789 25547 8823
rect 35265 8789 35299 8823
rect 36277 8789 36311 8823
rect 5457 8585 5491 8619
rect 15209 8585 15243 8619
rect 16129 8585 16163 8619
rect 17693 8585 17727 8619
rect 23213 8585 23247 8619
rect 25789 8585 25823 8619
rect 27537 8585 27571 8619
rect 29193 8585 29227 8619
rect 31309 8585 31343 8619
rect 31693 8585 31727 8619
rect 31861 8585 31895 8619
rect 35265 8585 35299 8619
rect 36737 8585 36771 8619
rect 5620 8517 5654 8551
rect 5825 8517 5859 8551
rect 8033 8517 8067 8551
rect 12817 8517 12851 8551
rect 15301 8517 15335 8551
rect 16037 8517 16071 8551
rect 21465 8517 21499 8551
rect 28181 8517 28215 8551
rect 29009 8517 29043 8551
rect 31493 8517 31527 8551
rect 33885 8517 33919 8551
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 5917 8449 5951 8483
rect 6009 8449 6043 8483
rect 6193 8449 6227 8483
rect 6561 8449 6595 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 7757 8449 7791 8483
rect 12541 8449 12575 8483
rect 22477 8449 22511 8483
rect 22845 8449 22879 8483
rect 23397 8449 23431 8483
rect 23489 8449 23523 8483
rect 23673 8449 23707 8483
rect 23857 8449 23891 8483
rect 23949 8449 23983 8483
rect 24041 8449 24075 8483
rect 24409 8449 24443 8483
rect 25237 8449 25271 8483
rect 25421 8449 25455 8483
rect 25513 8449 25547 8483
rect 25697 8449 25731 8483
rect 25881 8449 25915 8483
rect 25973 8449 26007 8483
rect 26065 8449 26099 8483
rect 27169 8449 27203 8483
rect 28089 8449 28123 8483
rect 28273 8449 28307 8483
rect 28549 8449 28583 8483
rect 28733 8449 28767 8483
rect 28825 8449 28859 8483
rect 31125 8449 31159 8483
rect 31401 8449 31435 8483
rect 34069 8449 34103 8483
rect 34345 8449 34379 8483
rect 34529 8449 34563 8483
rect 34897 8449 34931 8483
rect 36645 8449 36679 8483
rect 36829 8449 36863 8483
rect 7665 8381 7699 8415
rect 9597 8381 9631 8415
rect 9873 8381 9907 8415
rect 11345 8381 11379 8415
rect 12081 8381 12115 8415
rect 14289 8381 14323 8415
rect 15485 8381 15519 8415
rect 16221 8381 16255 8415
rect 17785 8381 17819 8415
rect 17969 8381 18003 8415
rect 19625 8381 19659 8415
rect 19993 8381 20027 8415
rect 21925 8381 21959 8415
rect 27077 8381 27111 8415
rect 28365 8381 28399 8415
rect 34621 8381 34655 8415
rect 34805 8381 34839 8415
rect 6193 8313 6227 8347
rect 24501 8313 24535 8347
rect 31125 8313 31159 8347
rect 34253 8313 34287 8347
rect 3985 8245 4019 8279
rect 5365 8245 5399 8279
rect 5641 8245 5675 8279
rect 9505 8245 9539 8279
rect 11529 8245 11563 8279
rect 14841 8245 14875 8279
rect 15669 8245 15703 8279
rect 17325 8245 17359 8279
rect 24317 8245 24351 8279
rect 31677 8245 31711 8279
rect 34437 8245 34471 8279
rect 3893 8041 3927 8075
rect 6837 8041 6871 8075
rect 7113 8041 7147 8075
rect 7297 8041 7331 8075
rect 7757 8041 7791 8075
rect 8309 8041 8343 8075
rect 9689 8041 9723 8075
rect 15853 8041 15887 8075
rect 18705 8041 18739 8075
rect 26893 8041 26927 8075
rect 27169 8041 27203 8075
rect 31125 8041 31159 8075
rect 37749 8041 37783 8075
rect 8217 7973 8251 8007
rect 21649 7973 21683 8007
rect 25145 7973 25179 8007
rect 28181 7973 28215 8007
rect 30113 7973 30147 8007
rect 36369 7973 36403 8007
rect 5089 7905 5123 7939
rect 7665 7905 7699 7939
rect 7941 7905 7975 7939
rect 9045 7905 9079 7939
rect 9965 7905 9999 7939
rect 14105 7905 14139 7939
rect 14381 7905 14415 7939
rect 16221 7905 16255 7939
rect 16405 7905 16439 7939
rect 17233 7905 17267 7939
rect 27537 7905 27571 7939
rect 27905 7905 27939 7939
rect 28917 7905 28951 7939
rect 29653 7905 29687 7939
rect 30941 7905 30975 7939
rect 33885 7905 33919 7939
rect 34345 7905 34379 7939
rect 37013 7905 37047 7939
rect 37841 7905 37875 7939
rect 4077 7837 4111 7871
rect 4261 7837 4295 7871
rect 4445 7837 4479 7871
rect 8033 7837 8067 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 10057 7837 10091 7871
rect 10517 7837 10551 7871
rect 16957 7837 16991 7871
rect 21373 7837 21407 7871
rect 21465 7837 21499 7871
rect 21741 7837 21775 7871
rect 22385 7837 22419 7871
rect 22477 7837 22511 7871
rect 22753 7837 22787 7871
rect 23029 7837 23063 7871
rect 23305 7837 23339 7871
rect 23765 7837 23799 7871
rect 23857 7837 23891 7871
rect 24041 7837 24075 7871
rect 24133 7837 24167 7871
rect 24416 7837 24450 7871
rect 24557 7837 24591 7871
rect 24777 7837 24811 7871
rect 24874 7837 24908 7871
rect 25145 7837 25179 7871
rect 25329 7837 25363 7871
rect 26801 7837 26835 7871
rect 26985 7837 27019 7871
rect 27077 7837 27111 7871
rect 27353 7837 27387 7871
rect 27813 7837 27847 7871
rect 28273 7837 28307 7871
rect 28457 7837 28491 7871
rect 28733 7837 28767 7871
rect 29745 7837 29779 7871
rect 30205 7837 30239 7871
rect 30573 7837 30607 7871
rect 30849 7837 30883 7871
rect 31309 7837 31343 7871
rect 31493 7837 31527 7871
rect 31769 7837 31803 7871
rect 34253 7837 34287 7871
rect 34713 7837 34747 7871
rect 34897 7837 34931 7871
rect 35173 7837 35207 7871
rect 35357 7837 35391 7871
rect 35633 7837 35667 7871
rect 36093 7837 36127 7871
rect 36369 7837 36403 7871
rect 36829 7837 36863 7871
rect 37289 7837 37323 7871
rect 37565 7837 37599 7871
rect 37933 7837 37967 7871
rect 38209 7837 38243 7871
rect 5365 7769 5399 7803
rect 7757 7769 7791 7803
rect 10793 7769 10827 7803
rect 21649 7769 21683 7803
rect 21925 7769 21959 7803
rect 22569 7769 22603 7803
rect 22845 7769 22879 7803
rect 23213 7769 23247 7803
rect 24685 7769 24719 7803
rect 30389 7769 30423 7803
rect 35449 7769 35483 7803
rect 37197 7769 37231 7803
rect 4997 7701 5031 7735
rect 7297 7701 7331 7735
rect 12265 7701 12299 7735
rect 16497 7701 16531 7735
rect 16865 7701 16899 7735
rect 22109 7701 22143 7735
rect 22201 7701 22235 7735
rect 23581 7701 23615 7735
rect 25053 7701 25087 7735
rect 31953 7701 31987 7735
rect 34713 7701 34747 7735
rect 35357 7701 35391 7735
rect 35817 7701 35851 7735
rect 36185 7701 36219 7735
rect 37381 7701 37415 7735
rect 38117 7701 38151 7735
rect 38393 7701 38427 7735
rect 4721 7497 4755 7531
rect 10333 7497 10367 7531
rect 11529 7497 11563 7531
rect 16221 7497 16255 7531
rect 18429 7497 18463 7531
rect 26985 7497 27019 7531
rect 27445 7497 27479 7531
rect 36829 7497 36863 7531
rect 2881 7429 2915 7463
rect 9965 7429 9999 7463
rect 10165 7429 10199 7463
rect 10425 7429 10459 7463
rect 14749 7429 14783 7463
rect 16957 7429 16991 7463
rect 22569 7429 22603 7463
rect 27169 7429 27203 7463
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 4905 7361 4939 7395
rect 5089 7361 5123 7395
rect 8217 7361 8251 7395
rect 14473 7361 14507 7395
rect 20913 7361 20947 7395
rect 21189 7361 21223 7395
rect 21373 7361 21407 7395
rect 21833 7361 21867 7395
rect 22845 7361 22879 7395
rect 22937 7361 22971 7395
rect 23029 7361 23063 7395
rect 23213 7361 23247 7395
rect 24041 7361 24075 7395
rect 24225 7361 24259 7395
rect 24317 7361 24351 7395
rect 24409 7361 24443 7395
rect 24593 7361 24627 7395
rect 24685 7361 24719 7395
rect 24778 7361 24812 7395
rect 24961 7361 24995 7395
rect 25053 7361 25087 7395
rect 25150 7361 25184 7395
rect 27353 7361 27387 7395
rect 27445 7361 27479 7395
rect 27629 7361 27663 7395
rect 32321 7361 32355 7395
rect 32781 7361 32815 7395
rect 32965 7361 32999 7395
rect 33149 7361 33183 7395
rect 33333 7361 33367 7395
rect 33425 7361 33459 7395
rect 33517 7361 33551 7395
rect 33701 7361 33735 7395
rect 35725 7361 35759 7395
rect 36185 7361 36219 7395
rect 36369 7361 36403 7395
rect 36461 7361 36495 7395
rect 36553 7361 36587 7395
rect 1409 7293 1443 7327
rect 2605 7293 2639 7327
rect 8401 7293 8435 7327
rect 11161 7293 11195 7327
rect 16681 7293 16715 7327
rect 22385 7293 22419 7327
rect 32229 7293 32263 7327
rect 32873 7293 32907 7327
rect 35817 7293 35851 7327
rect 32689 7225 32723 7259
rect 4353 7157 4387 7191
rect 4905 7157 4939 7191
rect 8033 7157 8067 7191
rect 10149 7157 10183 7191
rect 20729 7157 20763 7191
rect 23857 7157 23891 7191
rect 25329 7157 25363 7191
rect 33885 7157 33919 7191
rect 35449 7157 35483 7191
rect 3433 6953 3467 6987
rect 3985 6953 4019 6987
rect 5469 6953 5503 6987
rect 6456 6953 6490 6987
rect 19980 6953 20014 6987
rect 21465 6953 21499 6987
rect 27813 6953 27847 6987
rect 30389 6953 30423 6987
rect 36724 6953 36758 6987
rect 3617 6885 3651 6919
rect 1409 6817 1443 6851
rect 5733 6817 5767 6851
rect 6193 6817 6227 6851
rect 8953 6817 8987 6851
rect 12173 6817 12207 6851
rect 26249 6817 26283 6851
rect 27445 6817 27479 6851
rect 32781 6817 32815 6851
rect 34713 6817 34747 6851
rect 35817 6817 35851 6851
rect 36369 6817 36403 6851
rect 36461 6817 36495 6851
rect 38485 6817 38519 6851
rect 8585 6749 8619 6783
rect 11345 6749 11379 6783
rect 11529 6749 11563 6783
rect 11713 6749 11747 6783
rect 11805 6749 11839 6783
rect 14657 6749 14691 6783
rect 17693 6749 17727 6783
rect 17785 6749 17819 6783
rect 19717 6749 19751 6783
rect 22845 6749 22879 6783
rect 24869 6749 24903 6783
rect 25697 6749 25731 6783
rect 25881 6749 25915 6783
rect 26065 6749 26099 6783
rect 26157 6749 26191 6783
rect 26341 6749 26375 6783
rect 27537 6749 27571 6783
rect 29101 6749 29135 6783
rect 29285 6749 29319 6783
rect 29561 6749 29595 6783
rect 29745 6749 29779 6783
rect 32137 6749 32171 6783
rect 32689 6749 32723 6783
rect 32873 6749 32907 6783
rect 33425 6749 33459 6783
rect 33518 6749 33552 6783
rect 33793 6749 33827 6783
rect 33931 6749 33965 6783
rect 34805 6749 34839 6783
rect 34989 6749 35023 6783
rect 35633 6749 35667 6783
rect 1685 6681 1719 6715
rect 3249 6681 3283 6715
rect 9229 6681 9263 6715
rect 10885 6681 10919 6715
rect 12449 6681 12483 6715
rect 18521 6681 18555 6715
rect 29929 6681 29963 6715
rect 30021 6681 30055 6715
rect 30205 6681 30239 6715
rect 32321 6681 32355 6715
rect 33701 6681 33735 6715
rect 3157 6613 3191 6647
rect 3459 6613 3493 6647
rect 7941 6613 7975 6647
rect 8033 6613 8067 6647
rect 10701 6613 10735 6647
rect 13921 6613 13955 6647
rect 14105 6613 14139 6647
rect 22753 6613 22787 6647
rect 24777 6613 24811 6647
rect 29193 6613 29227 6647
rect 32505 6613 32539 6647
rect 34069 6613 34103 6647
rect 35173 6613 35207 6647
rect 35449 6613 35483 6647
rect 7205 6409 7239 6443
rect 8033 6409 8067 6443
rect 10333 6409 10367 6443
rect 23213 6409 23247 6443
rect 24409 6409 24443 6443
rect 26157 6409 26191 6443
rect 27261 6409 27295 6443
rect 28825 6409 28859 6443
rect 30849 6409 30883 6443
rect 33333 6409 33367 6443
rect 36093 6409 36127 6443
rect 4629 6341 4663 6375
rect 5273 6341 5307 6375
rect 7849 6341 7883 6375
rect 10701 6341 10735 6375
rect 12173 6341 12207 6375
rect 12449 6341 12483 6375
rect 13277 6341 13311 6375
rect 22937 6341 22971 6375
rect 25789 6341 25823 6375
rect 27905 6341 27939 6375
rect 31309 6341 31343 6375
rect 31953 6341 31987 6375
rect 32505 6341 32539 6375
rect 1409 6273 1443 6307
rect 2697 6273 2731 6307
rect 2973 6273 3007 6307
rect 3985 6273 4019 6307
rect 4721 6273 4755 6307
rect 4997 6273 5031 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 7389 6273 7423 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 7941 6273 7975 6307
rect 8309 6273 8343 6307
rect 8401 6273 8435 6307
rect 8493 6273 8527 6307
rect 8677 6273 8711 6307
rect 8769 6273 8803 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 11253 6273 11287 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 12357 6273 12391 6307
rect 12633 6273 12667 6307
rect 12725 6273 12759 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 13369 6273 13403 6307
rect 17969 6273 18003 6307
rect 22109 6273 22143 6307
rect 23305 6273 23339 6307
rect 23489 6273 23523 6307
rect 24317 6273 24351 6307
rect 24961 6273 24995 6307
rect 25145 6273 25179 6307
rect 25237 6273 25271 6307
rect 25329 6273 25363 6307
rect 25513 6273 25547 6307
rect 25973 6273 26007 6307
rect 26617 6273 26651 6307
rect 26801 6273 26835 6307
rect 27813 6273 27847 6307
rect 28089 6273 28123 6307
rect 28457 6273 28491 6307
rect 28917 6273 28951 6307
rect 29101 6273 29135 6307
rect 29377 6273 29411 6307
rect 29561 6273 29595 6307
rect 30481 6273 30515 6307
rect 30665 6273 30699 6307
rect 30941 6273 30975 6307
rect 31125 6273 31159 6307
rect 31217 6273 31251 6307
rect 31401 6273 31435 6307
rect 31585 6273 31619 6307
rect 31769 6273 31803 6307
rect 32137 6273 32171 6307
rect 32321 6273 32355 6307
rect 32413 6273 32447 6307
rect 32689 6273 32723 6307
rect 33149 6273 33183 6307
rect 34621 6273 34655 6307
rect 34769 6273 34803 6307
rect 34897 6273 34931 6307
rect 34989 6273 35023 6307
rect 35086 6273 35120 6307
rect 35541 6273 35575 6307
rect 35725 6273 35759 6307
rect 35817 6273 35851 6307
rect 35909 6273 35943 6307
rect 2329 6205 2363 6239
rect 2789 6205 2823 6239
rect 3617 6205 3651 6239
rect 4813 6205 4847 6239
rect 7665 6205 7699 6239
rect 8861 6205 8895 6239
rect 10124 6205 10158 6239
rect 10241 6205 10275 6239
rect 10609 6205 10643 6239
rect 22293 6205 22327 6239
rect 24593 6205 24627 6239
rect 27721 6205 27755 6239
rect 28365 6205 28399 6239
rect 31033 6205 31067 6239
rect 32873 6205 32907 6239
rect 32965 6205 32999 6239
rect 5273 6137 5307 6171
rect 10793 6137 10827 6171
rect 12633 6137 12667 6171
rect 23949 6137 23983 6171
rect 27353 6137 27387 6171
rect 28089 6137 28123 6171
rect 35265 6137 35299 6171
rect 4721 6069 4755 6103
rect 5181 6069 5215 6103
rect 9965 6069 9999 6103
rect 11161 6069 11195 6103
rect 11529 6069 11563 6103
rect 11989 6069 12023 6103
rect 23029 6069 23063 6103
rect 24777 6069 24811 6103
rect 26617 6069 26651 6103
rect 32229 6069 32263 6103
rect 5181 5865 5215 5899
rect 8217 5865 8251 5899
rect 8401 5865 8435 5899
rect 9597 5865 9631 5899
rect 10149 5865 10183 5899
rect 10517 5865 10551 5899
rect 11437 5865 11471 5899
rect 23489 5865 23523 5899
rect 26801 5865 26835 5899
rect 27629 5865 27663 5899
rect 30113 5865 30147 5899
rect 31953 5865 31987 5899
rect 32781 5865 32815 5899
rect 33793 5865 33827 5899
rect 34437 5865 34471 5899
rect 34713 5865 34747 5899
rect 35173 5865 35207 5899
rect 35633 5865 35667 5899
rect 10057 5797 10091 5831
rect 10793 5797 10827 5831
rect 11713 5797 11747 5831
rect 22937 5797 22971 5831
rect 25145 5797 25179 5831
rect 1869 5729 1903 5763
rect 3617 5729 3651 5763
rect 4629 5729 4663 5763
rect 4813 5729 4847 5763
rect 7757 5729 7791 5763
rect 7849 5729 7883 5763
rect 9505 5729 9539 5763
rect 9689 5729 9723 5763
rect 10425 5729 10459 5763
rect 10977 5729 11011 5763
rect 11437 5729 11471 5763
rect 12081 5729 12115 5763
rect 12357 5729 12391 5763
rect 12909 5729 12943 5763
rect 13185 5729 13219 5763
rect 15577 5729 15611 5763
rect 21741 5729 21775 5763
rect 22569 5729 22603 5763
rect 22753 5729 22787 5763
rect 23305 5729 23339 5763
rect 26341 5729 26375 5763
rect 1409 5661 1443 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 4077 5661 4111 5695
rect 4997 5661 5031 5695
rect 5641 5661 5675 5695
rect 5825 5661 5859 5695
rect 6653 5661 6687 5695
rect 7941 5661 7975 5695
rect 8033 5661 8067 5695
rect 9045 5661 9079 5695
rect 9137 5661 9171 5695
rect 9873 5661 9907 5695
rect 10517 5661 10551 5695
rect 10885 5661 10919 5695
rect 11529 5661 11563 5695
rect 11989 5661 12023 5695
rect 12173 5661 12207 5695
rect 12265 5661 12299 5695
rect 12449 5661 12483 5695
rect 12817 5661 12851 5695
rect 13277 5661 13311 5695
rect 13829 5661 13863 5695
rect 15853 5661 15887 5695
rect 22477 5661 22511 5695
rect 22937 5661 22971 5695
rect 23213 5661 23247 5695
rect 23581 5661 23615 5695
rect 24409 5661 24443 5695
rect 24557 5661 24591 5695
rect 24913 5661 24947 5695
rect 25145 5661 25179 5695
rect 25421 5661 25455 5695
rect 25881 5661 25915 5695
rect 25973 5661 26007 5695
rect 26157 5661 26191 5695
rect 26249 5661 26283 5695
rect 26433 5661 26467 5695
rect 27261 5661 27295 5695
rect 27445 5661 27479 5695
rect 31861 5661 31895 5695
rect 32045 5661 32079 5695
rect 32505 5661 32539 5695
rect 32781 5661 32815 5695
rect 33793 5661 33827 5695
rect 33977 5661 34011 5695
rect 34345 5661 34379 5695
rect 34529 5661 34563 5695
rect 34713 5661 34747 5695
rect 34897 5661 34931 5695
rect 35081 5661 35115 5695
rect 35357 5661 35391 5695
rect 35449 5661 35483 5695
rect 2145 5593 2179 5627
rect 8369 5593 8403 5627
rect 8585 5593 8619 5627
rect 9229 5593 9263 5627
rect 9321 5593 9355 5627
rect 9597 5593 9631 5627
rect 10609 5593 10643 5627
rect 11069 5593 11103 5627
rect 21557 5593 21591 5627
rect 23121 5593 23155 5627
rect 24685 5593 24719 5627
rect 24777 5593 24811 5627
rect 25329 5593 25363 5627
rect 26985 5593 27019 5627
rect 27169 5593 27203 5627
rect 29745 5593 29779 5627
rect 29929 5593 29963 5627
rect 32689 5593 32723 5627
rect 3893 5525 3927 5559
rect 5733 5525 5767 5559
rect 6101 5525 6135 5559
rect 7573 5525 7607 5559
rect 10701 5525 10735 5559
rect 14105 5525 14139 5559
rect 21189 5525 21223 5559
rect 21649 5525 21683 5559
rect 22109 5525 22143 5559
rect 23305 5525 23339 5559
rect 25053 5525 25087 5559
rect 2973 5321 3007 5355
rect 6377 5321 6411 5355
rect 6545 5321 6579 5355
rect 9597 5321 9631 5355
rect 13369 5321 13403 5355
rect 22017 5321 22051 5355
rect 22937 5321 22971 5355
rect 29561 5321 29595 5355
rect 31217 5321 31251 5355
rect 31953 5321 31987 5355
rect 32689 5321 32723 5355
rect 33349 5321 33383 5355
rect 33517 5321 33551 5355
rect 34621 5321 34655 5355
rect 35357 5321 35391 5355
rect 3893 5253 3927 5287
rect 6745 5253 6779 5287
rect 11989 5253 12023 5287
rect 12205 5253 12239 5287
rect 24869 5253 24903 5287
rect 25329 5253 25363 5287
rect 25421 5253 25455 5287
rect 25605 5253 25639 5287
rect 32413 5253 32447 5287
rect 33149 5253 33183 5287
rect 33885 5253 33919 5287
rect 2881 5185 2915 5219
rect 3065 5185 3099 5219
rect 4445 5185 4479 5219
rect 7113 5185 7147 5219
rect 7389 5185 7423 5219
rect 7573 5185 7607 5219
rect 9137 5185 9171 5219
rect 9413 5185 9447 5219
rect 11161 5185 11195 5219
rect 11897 5185 11931 5219
rect 13093 5185 13127 5219
rect 13185 5185 13219 5219
rect 13461 5185 13495 5219
rect 19809 5185 19843 5219
rect 21603 5185 21637 5219
rect 21833 5185 21867 5219
rect 22385 5185 22419 5219
rect 22477 5185 22511 5219
rect 22753 5185 22787 5219
rect 23029 5185 23063 5219
rect 25053 5185 25087 5219
rect 25237 5185 25271 5219
rect 29377 5185 29411 5219
rect 29653 5185 29687 5219
rect 29837 5185 29871 5219
rect 29929 5185 29963 5219
rect 30113 5185 30147 5219
rect 30849 5185 30883 5219
rect 31585 5185 31619 5219
rect 32137 5185 32171 5219
rect 32505 5185 32539 5219
rect 32689 5185 32723 5219
rect 33609 5185 33643 5219
rect 33701 5185 33735 5219
rect 34253 5185 34287 5219
rect 34437 5185 34471 5219
rect 34713 5185 34747 5219
rect 34897 5185 34931 5219
rect 35173 5185 35207 5219
rect 1409 5117 1443 5151
rect 4721 5117 4755 5151
rect 9229 5117 9263 5151
rect 12449 5117 12483 5151
rect 20177 5117 20211 5151
rect 28641 5117 28675 5151
rect 29193 5117 29227 5151
rect 30021 5117 30055 5151
rect 30757 5117 30791 5151
rect 31677 5117 31711 5151
rect 32413 5117 32447 5151
rect 6193 5049 6227 5083
rect 11345 5049 11379 5083
rect 22661 5049 22695 5083
rect 28917 5049 28951 5083
rect 29101 5049 29135 5083
rect 29837 5049 29871 5083
rect 32229 5049 32263 5083
rect 33885 5049 33919 5083
rect 6561 4981 6595 5015
rect 6929 4981 6963 5015
rect 9413 4981 9447 5015
rect 11713 4981 11747 5015
rect 12173 4981 12207 5015
rect 12357 4981 12391 5015
rect 13185 4981 13219 5015
rect 22201 4981 22235 5015
rect 25789 4981 25823 5015
rect 31585 4981 31619 5015
rect 33333 4981 33367 5015
rect 6009 4777 6043 4811
rect 8309 4777 8343 4811
rect 9413 4777 9447 4811
rect 9689 4777 9723 4811
rect 10885 4777 10919 4811
rect 11161 4777 11195 4811
rect 23305 4777 23339 4811
rect 25789 4777 25823 4811
rect 27721 4777 27755 4811
rect 28917 4777 28951 4811
rect 33701 4777 33735 4811
rect 34069 4777 34103 4811
rect 34161 4777 34195 4811
rect 35357 4777 35391 4811
rect 4169 4709 4203 4743
rect 22753 4709 22787 4743
rect 23581 4709 23615 4743
rect 27077 4709 27111 4743
rect 34253 4709 34287 4743
rect 4997 4641 5031 4675
rect 6561 4641 6595 4675
rect 6837 4641 6871 4675
rect 9045 4641 9079 4675
rect 12173 4641 12207 4675
rect 13921 4641 13955 4675
rect 19257 4641 19291 4675
rect 21281 4641 21315 4675
rect 26433 4641 26467 4675
rect 27537 4641 27571 4675
rect 28641 4641 28675 4675
rect 33609 4641 33643 4675
rect 34437 4641 34471 4675
rect 3893 4573 3927 4607
rect 4169 4573 4203 4607
rect 5273 4573 5307 4607
rect 5825 4573 5859 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 6285 4573 6319 4607
rect 9137 4573 9171 4607
rect 9505 4573 9539 4607
rect 10517 4573 10551 4607
rect 10609 4573 10643 4607
rect 10977 4573 11011 4607
rect 22477 4573 22511 4607
rect 22937 4573 22971 4607
rect 23397 4573 23431 4607
rect 23949 4573 23983 4607
rect 24133 4573 24167 4607
rect 26157 4573 26191 4607
rect 26801 4573 26835 4607
rect 27445 4573 27479 4607
rect 28549 4573 28583 4607
rect 33885 4573 33919 4607
rect 34161 4573 34195 4607
rect 35081 4573 35115 4607
rect 35173 4573 35207 4607
rect 4261 4505 4295 4539
rect 13645 4505 13679 4539
rect 19533 4505 19567 4539
rect 22753 4505 22787 4539
rect 23121 4505 23155 4539
rect 27077 4505 27111 4539
rect 1409 4437 1443 4471
rect 3985 4437 4019 4471
rect 22569 4437 22603 4471
rect 24041 4437 24075 4471
rect 26249 4437 26283 4471
rect 26893 4437 26927 4471
rect 34713 4437 34747 4471
rect 5365 4233 5399 4267
rect 10961 4233 10995 4267
rect 12541 4233 12575 4267
rect 22401 4233 22435 4267
rect 22569 4233 22603 4267
rect 26157 4233 26191 4267
rect 27353 4233 27387 4267
rect 28181 4233 28215 4267
rect 28917 4233 28951 4267
rect 31677 4233 31711 4267
rect 33517 4233 33551 4267
rect 11161 4165 11195 4199
rect 22201 4165 22235 4199
rect 23857 4165 23891 4199
rect 25145 4165 25179 4199
rect 26433 4165 26467 4199
rect 26649 4165 26683 4199
rect 27813 4165 27847 4199
rect 3249 4097 3283 4131
rect 5733 4097 5767 4131
rect 5917 4097 5951 4131
rect 6377 4097 6411 4131
rect 6653 4097 6687 4131
rect 7665 4097 7699 4131
rect 7849 4097 7883 4131
rect 8585 4097 8619 4131
rect 8769 4097 8803 4131
rect 10333 4097 10367 4131
rect 10517 4097 10551 4131
rect 11529 4097 11563 4131
rect 11713 4097 11747 4131
rect 12449 4097 12483 4131
rect 12633 4097 12667 4131
rect 22109 4097 22143 4131
rect 23305 4097 23339 4131
rect 23673 4097 23707 4131
rect 23765 4097 23799 4131
rect 24041 4097 24075 4131
rect 24317 4097 24351 4131
rect 24777 4097 24811 4131
rect 25329 4097 25363 4131
rect 25513 4097 25547 4131
rect 26157 4097 26191 4131
rect 26341 4097 26375 4131
rect 27997 4097 28031 4131
rect 29561 4097 29595 4131
rect 29653 4097 29687 4131
rect 29837 4097 29871 4131
rect 31033 4097 31067 4131
rect 31309 4097 31343 4131
rect 31493 4097 31527 4131
rect 31585 4097 31619 4131
rect 31769 4097 31803 4131
rect 32628 4097 32662 4131
rect 33057 4097 33091 4131
rect 3525 4029 3559 4063
rect 6469 4029 6503 4063
rect 11621 4029 11655 4063
rect 22017 4029 22051 4063
rect 24869 4029 24903 4063
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 27445 4029 27479 4063
rect 27537 4029 27571 4063
rect 29101 4029 29135 4063
rect 29193 4029 29227 4063
rect 30757 4029 30791 4063
rect 31217 4029 31251 4063
rect 32505 4029 32539 4063
rect 32965 4029 32999 4063
rect 6837 3961 6871 3995
rect 10793 3961 10827 3995
rect 24133 3961 24167 3995
rect 24593 3961 24627 3995
rect 25513 3961 25547 3995
rect 26801 3961 26835 3995
rect 29745 3961 29779 3995
rect 31401 3961 31435 3995
rect 33333 3961 33367 3995
rect 4997 3893 5031 3927
rect 5733 3893 5767 3927
rect 6561 3893 6595 3927
rect 7849 3893 7883 3927
rect 8769 3893 8803 3927
rect 10517 3893 10551 3927
rect 10977 3893 11011 3927
rect 22385 3893 22419 3927
rect 23489 3893 23523 3927
rect 26617 3893 26651 3927
rect 26985 3893 27019 3927
rect 30849 3893 30883 3927
rect 3801 3689 3835 3723
rect 4077 3689 4111 3723
rect 4261 3689 4295 3723
rect 7113 3689 7147 3723
rect 7941 3689 7975 3723
rect 8493 3689 8527 3723
rect 9965 3689 9999 3723
rect 10885 3689 10919 3723
rect 22845 3689 22879 3723
rect 23949 3689 23983 3723
rect 25053 3689 25087 3723
rect 25421 3689 25455 3723
rect 27905 3689 27939 3723
rect 29193 3689 29227 3723
rect 30297 3689 30331 3723
rect 31125 3689 31159 3723
rect 31677 3689 31711 3723
rect 32045 3689 32079 3723
rect 32321 3689 32355 3723
rect 1409 3621 1443 3655
rect 8309 3621 8343 3655
rect 25973 3621 26007 3655
rect 27629 3621 27663 3655
rect 28641 3621 28675 3655
rect 30021 3621 30055 3655
rect 5365 3553 5399 3587
rect 5641 3553 5675 3587
rect 10149 3553 10183 3587
rect 10241 3553 10275 3587
rect 11161 3553 11195 3587
rect 11805 3553 11839 3587
rect 12357 3553 12391 3587
rect 21097 3553 21131 3587
rect 24585 3553 24619 3587
rect 24777 3553 24811 3587
rect 26893 3553 26927 3587
rect 24869 3519 24903 3553
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 5089 3485 5123 3519
rect 7757 3485 7791 3519
rect 8217 3485 8251 3519
rect 8953 3485 8987 3519
rect 9689 3485 9723 3519
rect 10057 3485 10091 3519
rect 11069 3485 11103 3519
rect 11253 3485 11287 3519
rect 11529 3485 11563 3519
rect 11713 3485 11747 3519
rect 12081 3485 12115 3519
rect 12173 3485 12207 3519
rect 13001 3485 13035 3519
rect 23857 3485 23891 3519
rect 24685 3485 24719 3519
rect 25237 3485 25271 3519
rect 25513 3485 25547 3519
rect 25789 3485 25823 3519
rect 26065 3485 26099 3519
rect 26249 3485 26283 3519
rect 26433 3485 26467 3519
rect 26985 3485 27019 3519
rect 27353 3485 27387 3519
rect 27445 3485 27479 3519
rect 27629 3485 27663 3519
rect 27721 3485 27755 3519
rect 27905 3485 27939 3519
rect 28549 3485 28583 3519
rect 28733 3485 28767 3519
rect 29009 3485 29043 3519
rect 29745 3485 29779 3519
rect 29837 3485 29871 3519
rect 30665 3485 30699 3519
rect 30757 3485 30791 3519
rect 30941 3485 30975 3519
rect 31217 3485 31251 3519
rect 31401 3485 31435 3519
rect 31585 3485 31619 3519
rect 31677 3485 31711 3519
rect 31769 3485 31803 3519
rect 32137 3485 32171 3519
rect 32321 3485 32355 3519
rect 38485 3485 38519 3519
rect 4445 3417 4479 3451
rect 7941 3417 7975 3451
rect 8677 3417 8711 3451
rect 11897 3417 11931 3451
rect 21373 3417 21407 3451
rect 23121 3417 23155 3451
rect 25605 3417 25639 3451
rect 26543 3417 26577 3451
rect 26709 3417 26743 3451
rect 28825 3417 28859 3451
rect 30021 3417 30055 3451
rect 30113 3417 30147 3451
rect 4235 3349 4269 3383
rect 4537 3349 4571 3383
rect 7205 3349 7239 3383
rect 8125 3349 8159 3383
rect 8477 3349 8511 3383
rect 9597 3349 9631 3383
rect 9781 3349 9815 3383
rect 11345 3349 11379 3383
rect 24409 3349 24443 3383
rect 27169 3349 27203 3383
rect 30313 3349 30347 3383
rect 30481 3349 30515 3383
rect 5641 3145 5675 3179
rect 6009 3145 6043 3179
rect 7757 3145 7791 3179
rect 13277 3145 13311 3179
rect 24225 3145 24259 3179
rect 26525 3145 26559 3179
rect 27077 3145 27111 3179
rect 30113 3145 30147 3179
rect 31033 3145 31067 3179
rect 31401 3145 31435 3179
rect 9229 3077 9263 3111
rect 11805 3077 11839 3111
rect 22477 3077 22511 3111
rect 31125 3077 31159 3111
rect 3433 3009 3467 3043
rect 3893 3009 3927 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 6561 3009 6595 3043
rect 6745 3009 6779 3043
rect 11345 3009 11379 3043
rect 11529 3009 11563 3043
rect 22201 3009 22235 3043
rect 24133 3009 24167 3043
rect 24317 3009 24351 3043
rect 24501 3009 24535 3043
rect 24869 3009 24903 3043
rect 26433 3009 26467 3043
rect 26617 3009 26651 3043
rect 26985 3009 27019 3043
rect 27181 3009 27215 3043
rect 28089 3009 28123 3043
rect 30021 3009 30055 3043
rect 30757 3009 30791 3043
rect 30849 3009 30883 3043
rect 31309 3009 31343 3043
rect 31401 3009 31435 3043
rect 1409 2941 1443 2975
rect 3525 2941 3559 2975
rect 3801 2941 3835 2975
rect 4169 2941 4203 2975
rect 9505 2941 9539 2975
rect 9597 2941 9631 2975
rect 11069 2941 11103 2975
rect 28181 2941 28215 2975
rect 28457 2941 28491 2975
rect 31033 2941 31067 2975
rect 38485 2941 38519 2975
rect 6377 2873 6411 2907
rect 26295 2873 26329 2907
rect 7205 2805 7239 2839
rect 23949 2805 23983 2839
rect 8953 2601 8987 2635
rect 15117 2601 15151 2635
rect 6929 2465 6963 2499
rect 7205 2465 7239 2499
rect 8677 2465 8711 2499
rect 9505 2465 9539 2499
rect 5273 2397 5307 2431
rect 14933 2397 14967 2431
rect 21373 2397 21407 2431
rect 23949 2397 23983 2431
rect 29745 2397 29779 2431
rect 30389 2397 30423 2431
rect 35541 2397 35575 2431
rect 36185 2397 36219 2431
rect 14841 2261 14875 2295
rect 21557 2261 21591 2295
rect 24593 2261 24627 2295
rect 27169 2261 27203 2295
rect 27813 2261 27847 2295
rect 29101 2261 29135 2295
rect 38485 2261 38519 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1302 37408 1308 37460
rect 1360 37448 1366 37460
rect 1673 37451 1731 37457
rect 1673 37448 1685 37451
rect 1360 37420 1685 37448
rect 1360 37408 1366 37420
rect 1673 37417 1685 37420
rect 1719 37417 1731 37451
rect 1673 37411 1731 37417
rect 3234 37408 3240 37460
rect 3292 37448 3298 37460
rect 3329 37451 3387 37457
rect 3329 37448 3341 37451
rect 3292 37420 3341 37448
rect 3292 37408 3298 37420
rect 3329 37417 3341 37420
rect 3375 37417 3387 37451
rect 3329 37411 3387 37417
rect 27706 37408 27712 37460
rect 27764 37448 27770 37460
rect 27801 37451 27859 37457
rect 27801 37448 27813 37451
rect 27764 37420 27813 37448
rect 27764 37408 27770 37420
rect 27801 37417 27813 37420
rect 27847 37417 27859 37451
rect 27801 37411 27859 37417
rect 28994 37408 29000 37460
rect 29052 37448 29058 37460
rect 29089 37451 29147 37457
rect 29089 37448 29101 37451
rect 29052 37420 29101 37448
rect 29052 37408 29058 37420
rect 29089 37417 29101 37420
rect 29135 37417 29147 37451
rect 29089 37411 29147 37417
rect 29638 37408 29644 37460
rect 29696 37448 29702 37460
rect 29733 37451 29791 37457
rect 29733 37448 29745 37451
rect 29696 37420 29745 37448
rect 29696 37408 29702 37420
rect 29733 37417 29745 37420
rect 29779 37417 29791 37451
rect 29733 37411 29791 37417
rect 34146 37408 34152 37460
rect 34204 37448 34210 37460
rect 34241 37451 34299 37457
rect 34241 37448 34253 37451
rect 34204 37420 34253 37448
rect 34204 37408 34210 37420
rect 34241 37417 34253 37420
rect 34287 37417 34299 37451
rect 34241 37411 34299 37417
rect 34790 37408 34796 37460
rect 34848 37448 34854 37460
rect 34885 37451 34943 37457
rect 34885 37448 34897 37451
rect 34848 37420 34897 37448
rect 34848 37408 34854 37420
rect 34885 37417 34897 37420
rect 34931 37417 34943 37451
rect 34885 37411 34943 37417
rect 35434 37408 35440 37460
rect 35492 37448 35498 37460
rect 35529 37451 35587 37457
rect 35529 37448 35541 37451
rect 35492 37420 35541 37448
rect 35492 37408 35498 37420
rect 35529 37417 35541 37420
rect 35575 37417 35587 37451
rect 35529 37411 35587 37417
rect 36078 37408 36084 37460
rect 36136 37448 36142 37460
rect 36173 37451 36231 37457
rect 36173 37448 36185 37451
rect 36136 37420 36185 37448
rect 36136 37408 36142 37420
rect 36173 37417 36185 37420
rect 36219 37417 36231 37451
rect 36173 37411 36231 37417
rect 36722 37408 36728 37460
rect 36780 37448 36786 37460
rect 36817 37451 36875 37457
rect 36817 37448 36829 37451
rect 36780 37420 36829 37448
rect 36780 37408 36786 37420
rect 36817 37417 36829 37420
rect 36863 37417 36875 37451
rect 36817 37411 36875 37417
rect 37918 37408 37924 37460
rect 37976 37408 37982 37460
rect 38194 37408 38200 37460
rect 38252 37408 38258 37460
rect 842 37272 848 37324
rect 900 37312 906 37324
rect 1397 37315 1455 37321
rect 1397 37312 1409 37315
rect 900 37284 1409 37312
rect 900 37272 906 37284
rect 1397 37281 1409 37284
rect 1443 37281 1455 37315
rect 1397 37275 1455 37281
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5261 37247 5319 37253
rect 5261 37244 5273 37247
rect 5224 37216 5273 37244
rect 5224 37204 5230 37216
rect 5261 37213 5273 37216
rect 5307 37213 5319 37247
rect 5261 37207 5319 37213
rect 8110 37204 8116 37256
rect 8168 37244 8174 37256
rect 8205 37247 8263 37253
rect 8205 37244 8217 37247
rect 8168 37216 8217 37244
rect 8168 37204 8174 37216
rect 8205 37213 8217 37216
rect 8251 37213 8263 37247
rect 8205 37207 8263 37213
rect 24210 37204 24216 37256
rect 24268 37204 24274 37256
rect 25498 37204 25504 37256
rect 25556 37204 25562 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25700 37216 25881 37244
rect 20806 37136 20812 37188
rect 20864 37136 20870 37188
rect 20993 37179 21051 37185
rect 20993 37145 21005 37179
rect 21039 37176 21051 37179
rect 21174 37176 21180 37188
rect 21039 37148 21180 37176
rect 21039 37145 21051 37148
rect 20993 37139 21051 37145
rect 21174 37136 21180 37148
rect 21232 37136 21238 37188
rect 6822 37068 6828 37120
rect 6880 37108 6886 37120
rect 7653 37111 7711 37117
rect 7653 37108 7665 37111
rect 6880 37080 7665 37108
rect 6880 37068 6886 37080
rect 7653 37077 7665 37080
rect 7699 37077 7711 37111
rect 7653 37071 7711 37077
rect 19610 37068 19616 37120
rect 19668 37108 19674 37120
rect 20625 37111 20683 37117
rect 20625 37108 20637 37111
rect 19668 37080 20637 37108
rect 19668 37068 19674 37080
rect 20625 37077 20637 37080
rect 20671 37077 20683 37111
rect 20625 37071 20683 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 25700 37117 25728 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 26789 37247 26847 37253
rect 26789 37213 26801 37247
rect 26835 37244 26847 37247
rect 26970 37244 26976 37256
rect 26835 37216 26976 37244
rect 26835 37213 26847 37216
rect 26789 37207 26847 37213
rect 26970 37204 26976 37216
rect 27028 37204 27034 37256
rect 27062 37204 27068 37256
rect 27120 37244 27126 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 27120 37216 27169 37244
rect 27120 37204 27126 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 28350 37204 28356 37256
rect 28408 37244 28414 37256
rect 28445 37247 28503 37253
rect 28445 37244 28457 37247
rect 28408 37216 28457 37244
rect 28408 37204 28414 37216
rect 28445 37213 28457 37216
rect 28491 37213 28503 37247
rect 28445 37207 28503 37213
rect 30282 37204 30288 37256
rect 30340 37244 30346 37256
rect 30377 37247 30435 37253
rect 30377 37244 30389 37247
rect 30340 37216 30389 37244
rect 30340 37204 30346 37216
rect 30377 37213 30389 37216
rect 30423 37213 30435 37247
rect 30377 37207 30435 37213
rect 30926 37204 30932 37256
rect 30984 37244 30990 37256
rect 31021 37247 31079 37253
rect 31021 37244 31033 37247
rect 30984 37216 31033 37244
rect 30984 37204 30990 37216
rect 31021 37213 31033 37216
rect 31067 37213 31079 37247
rect 31021 37207 31079 37213
rect 31570 37204 31576 37256
rect 31628 37244 31634 37256
rect 31665 37247 31723 37253
rect 31665 37244 31677 37247
rect 31628 37216 31677 37244
rect 31628 37204 31634 37216
rect 31665 37213 31677 37216
rect 31711 37213 31723 37247
rect 31665 37207 31723 37213
rect 32214 37204 32220 37256
rect 32272 37244 32278 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 32272 37216 32321 37244
rect 32272 37204 32278 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 32309 37207 32367 37213
rect 32858 37204 32864 37256
rect 32916 37244 32922 37256
rect 32953 37247 33011 37253
rect 32953 37244 32965 37247
rect 32916 37216 32965 37244
rect 32916 37204 32922 37216
rect 32953 37213 32965 37216
rect 32999 37213 33011 37247
rect 32953 37207 33011 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33597 37247 33655 37253
rect 33597 37244 33609 37247
rect 33560 37216 33609 37244
rect 33560 37204 33566 37216
rect 33597 37213 33609 37216
rect 33643 37213 33655 37247
rect 33597 37207 33655 37213
rect 24029 37111 24087 37117
rect 24029 37108 24041 37111
rect 23900 37080 24041 37108
rect 23900 37068 23906 37080
rect 24029 37077 24041 37080
rect 24075 37077 24087 37111
rect 24029 37071 24087 37077
rect 25685 37111 25743 37117
rect 25685 37077 25697 37111
rect 25731 37077 25743 37111
rect 25685 37071 25743 37077
rect 25774 37068 25780 37120
rect 25832 37108 25838 37120
rect 26053 37111 26111 37117
rect 26053 37108 26065 37111
rect 25832 37080 26065 37108
rect 25832 37068 25838 37080
rect 26053 37077 26065 37080
rect 26099 37077 26111 37111
rect 26053 37071 26111 37077
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 26605 37111 26663 37117
rect 26605 37108 26617 37111
rect 26476 37080 26617 37108
rect 26476 37068 26482 37080
rect 26605 37077 26617 37080
rect 26651 37077 26663 37111
rect 26605 37071 26663 37077
rect 38470 37068 38476 37120
rect 38528 37068 38534 37120
rect 1104 37018 38824 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 38824 37018
rect 1104 36944 38824 36966
rect 19797 36907 19855 36913
rect 19797 36873 19809 36907
rect 19843 36904 19855 36907
rect 19843 36876 20208 36904
rect 19843 36873 19855 36876
rect 19797 36867 19855 36873
rect 5718 36796 5724 36848
rect 5776 36796 5782 36848
rect 19426 36796 19432 36848
rect 19484 36796 19490 36848
rect 19645 36839 19703 36845
rect 19645 36805 19657 36839
rect 19691 36836 19703 36839
rect 20070 36836 20076 36848
rect 19691 36808 20076 36836
rect 19691 36805 19703 36808
rect 19645 36799 19703 36805
rect 20070 36796 20076 36808
rect 20128 36796 20134 36848
rect 20180 36845 20208 36876
rect 20806 36864 20812 36916
rect 20864 36904 20870 36916
rect 21637 36907 21695 36913
rect 21637 36904 21649 36907
rect 20864 36876 21649 36904
rect 20864 36864 20870 36876
rect 21637 36873 21649 36876
rect 21683 36904 21695 36907
rect 21726 36904 21732 36916
rect 21683 36876 21732 36904
rect 21683 36873 21695 36876
rect 21637 36867 21695 36873
rect 21726 36864 21732 36876
rect 21784 36864 21790 36916
rect 24210 36864 24216 36916
rect 24268 36864 24274 36916
rect 26970 36864 26976 36916
rect 27028 36864 27034 36916
rect 29365 36907 29423 36913
rect 29365 36873 29377 36907
rect 29411 36904 29423 36907
rect 30098 36904 30104 36916
rect 29411 36876 30104 36904
rect 29411 36873 29423 36876
rect 29365 36867 29423 36873
rect 30098 36864 30104 36876
rect 30156 36864 30162 36916
rect 20165 36839 20223 36845
rect 20165 36805 20177 36839
rect 20211 36805 20223 36839
rect 23934 36836 23940 36848
rect 23874 36808 23940 36836
rect 20165 36799 20223 36805
rect 23934 36796 23940 36808
rect 23992 36796 23998 36848
rect 27982 36836 27988 36848
rect 26358 36808 27988 36836
rect 27982 36796 27988 36808
rect 28040 36836 28046 36848
rect 31846 36836 31852 36848
rect 28040 36808 28382 36836
rect 30498 36808 31852 36836
rect 28040 36796 28046 36808
rect 31846 36796 31852 36808
rect 31904 36796 31910 36848
rect 8202 36728 8208 36780
rect 8260 36728 8266 36780
rect 8386 36728 8392 36780
rect 8444 36768 8450 36780
rect 8665 36771 8723 36777
rect 8665 36768 8677 36771
rect 8444 36740 8677 36768
rect 8444 36728 8450 36740
rect 8665 36737 8677 36740
rect 8711 36737 8723 36771
rect 8665 36731 8723 36737
rect 8757 36771 8815 36777
rect 8757 36737 8769 36771
rect 8803 36737 8815 36771
rect 8757 36731 8815 36737
rect 4433 36703 4491 36709
rect 4433 36669 4445 36703
rect 4479 36700 4491 36703
rect 4709 36703 4767 36709
rect 4479 36672 4568 36700
rect 4479 36669 4491 36672
rect 4433 36663 4491 36669
rect 4540 36564 4568 36672
rect 4709 36669 4721 36703
rect 4755 36700 4767 36703
rect 5166 36700 5172 36712
rect 4755 36672 5172 36700
rect 4755 36669 4767 36672
rect 4709 36663 4767 36669
rect 5166 36660 5172 36672
rect 5224 36660 5230 36712
rect 6546 36660 6552 36712
rect 6604 36700 6610 36712
rect 6825 36703 6883 36709
rect 6825 36700 6837 36703
rect 6604 36672 6837 36700
rect 6604 36660 6610 36672
rect 6825 36669 6837 36672
rect 6871 36669 6883 36703
rect 6825 36663 6883 36669
rect 7101 36703 7159 36709
rect 7101 36669 7113 36703
rect 7147 36700 7159 36703
rect 7190 36700 7196 36712
rect 7147 36672 7196 36700
rect 7147 36669 7159 36672
rect 7101 36663 7159 36669
rect 7190 36660 7196 36672
rect 7248 36660 7254 36712
rect 6564 36632 6592 36660
rect 8772 36632 8800 36731
rect 8938 36728 8944 36780
rect 8996 36728 9002 36780
rect 19242 36660 19248 36712
rect 19300 36700 19306 36712
rect 19889 36703 19947 36709
rect 19889 36700 19901 36703
rect 19300 36672 19901 36700
rect 19300 36660 19306 36672
rect 19889 36669 19901 36672
rect 19935 36669 19947 36703
rect 21284 36700 21312 36754
rect 24394 36728 24400 36780
rect 24452 36728 24458 36780
rect 27154 36728 27160 36780
rect 27212 36728 27218 36780
rect 38197 36771 38255 36777
rect 38197 36737 38209 36771
rect 38243 36768 38255 36771
rect 38286 36768 38292 36780
rect 38243 36740 38292 36768
rect 38243 36737 38255 36740
rect 38197 36731 38255 36737
rect 38286 36728 38292 36740
rect 38344 36728 38350 36780
rect 38473 36771 38531 36777
rect 38473 36737 38485 36771
rect 38519 36768 38531 36771
rect 38562 36768 38568 36780
rect 38519 36740 38568 36768
rect 38519 36737 38531 36740
rect 38473 36731 38531 36737
rect 38562 36728 38568 36740
rect 38620 36728 38626 36780
rect 21358 36700 21364 36712
rect 21284 36672 21364 36700
rect 19889 36663 19947 36669
rect 21358 36660 21364 36672
rect 21416 36660 21422 36712
rect 22373 36703 22431 36709
rect 22373 36669 22385 36703
rect 22419 36700 22431 36703
rect 22419 36672 22508 36700
rect 22419 36669 22431 36672
rect 22373 36663 22431 36669
rect 5736 36604 6592 36632
rect 8588 36604 8800 36632
rect 5736 36564 5764 36604
rect 4540 36536 5764 36564
rect 6178 36524 6184 36576
rect 6236 36524 6242 36576
rect 7282 36524 7288 36576
rect 7340 36564 7346 36576
rect 8110 36564 8116 36576
rect 7340 36536 8116 36564
rect 7340 36524 7346 36536
rect 8110 36524 8116 36536
rect 8168 36564 8174 36576
rect 8588 36573 8616 36604
rect 8573 36567 8631 36573
rect 8573 36564 8585 36567
rect 8168 36536 8585 36564
rect 8168 36524 8174 36536
rect 8573 36533 8585 36536
rect 8619 36533 8631 36567
rect 8573 36527 8631 36533
rect 8662 36524 8668 36576
rect 8720 36564 8726 36576
rect 8941 36567 8999 36573
rect 8941 36564 8953 36567
rect 8720 36536 8953 36564
rect 8720 36524 8726 36536
rect 8941 36533 8953 36536
rect 8987 36533 8999 36567
rect 8941 36527 8999 36533
rect 19610 36524 19616 36576
rect 19668 36524 19674 36576
rect 22480 36564 22508 36672
rect 22646 36660 22652 36712
rect 22704 36660 22710 36712
rect 24854 36660 24860 36712
rect 24912 36660 24918 36712
rect 25130 36660 25136 36712
rect 25188 36660 25194 36712
rect 27522 36660 27528 36712
rect 27580 36700 27586 36712
rect 27617 36703 27675 36709
rect 27617 36700 27629 36703
rect 27580 36672 27629 36700
rect 27580 36660 27586 36672
rect 27617 36669 27629 36672
rect 27663 36669 27675 36703
rect 27617 36663 27675 36669
rect 27893 36703 27951 36709
rect 27893 36669 27905 36703
rect 27939 36700 27951 36703
rect 28350 36700 28356 36712
rect 27939 36672 28356 36700
rect 27939 36669 27951 36672
rect 27893 36663 27951 36669
rect 28350 36660 28356 36672
rect 28408 36660 28414 36712
rect 29362 36660 29368 36712
rect 29420 36700 29426 36712
rect 30929 36703 30987 36709
rect 30929 36700 30941 36703
rect 29420 36672 30941 36700
rect 29420 36660 29426 36672
rect 30929 36669 30941 36672
rect 30975 36669 30987 36703
rect 30929 36663 30987 36669
rect 31205 36703 31263 36709
rect 31205 36669 31217 36703
rect 31251 36700 31263 36703
rect 33134 36700 33140 36712
rect 31251 36672 33140 36700
rect 31251 36669 31263 36672
rect 31205 36663 31263 36669
rect 33134 36660 33140 36672
rect 33192 36660 33198 36712
rect 24872 36632 24900 36660
rect 23676 36604 24900 36632
rect 23676 36564 23704 36604
rect 22480 36536 23704 36564
rect 24118 36524 24124 36576
rect 24176 36524 24182 36576
rect 26602 36524 26608 36576
rect 26660 36524 26666 36576
rect 29454 36524 29460 36576
rect 29512 36524 29518 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 4433 36363 4491 36369
rect 4433 36329 4445 36363
rect 4479 36360 4491 36363
rect 4479 36332 4936 36360
rect 4479 36329 4491 36332
rect 4433 36323 4491 36329
rect 842 36252 848 36304
rect 900 36292 906 36304
rect 1397 36295 1455 36301
rect 1397 36292 1409 36295
rect 900 36264 1409 36292
rect 900 36252 906 36264
rect 1397 36261 1409 36264
rect 1443 36261 1455 36295
rect 1397 36255 1455 36261
rect 3326 36184 3332 36236
rect 3384 36224 3390 36236
rect 3384 36196 4752 36224
rect 3384 36184 3390 36196
rect 4430 36116 4436 36168
rect 4488 36116 4494 36168
rect 4724 36165 4752 36196
rect 4617 36159 4675 36165
rect 4617 36158 4629 36159
rect 4540 36130 4629 36158
rect 4540 36088 4568 36130
rect 4617 36125 4629 36130
rect 4663 36125 4675 36159
rect 4617 36119 4675 36125
rect 4709 36159 4767 36165
rect 4709 36125 4721 36159
rect 4755 36125 4767 36159
rect 4908 36156 4936 36332
rect 5166 36320 5172 36372
rect 5224 36320 5230 36372
rect 7190 36320 7196 36372
rect 7248 36320 7254 36372
rect 7466 36320 7472 36372
rect 7524 36360 7530 36372
rect 8110 36360 8116 36372
rect 7524 36332 8116 36360
rect 7524 36320 7530 36332
rect 8110 36320 8116 36332
rect 8168 36320 8174 36372
rect 8938 36320 8944 36372
rect 8996 36320 9002 36372
rect 20070 36320 20076 36372
rect 20128 36360 20134 36372
rect 21177 36363 21235 36369
rect 21177 36360 21189 36363
rect 20128 36332 21189 36360
rect 20128 36320 20134 36332
rect 21177 36329 21189 36332
rect 21223 36360 21235 36363
rect 21223 36332 21395 36360
rect 21223 36329 21235 36332
rect 21177 36323 21235 36329
rect 4985 36295 5043 36301
rect 4985 36261 4997 36295
rect 5031 36292 5043 36295
rect 5258 36292 5264 36304
rect 5031 36264 5264 36292
rect 5031 36261 5043 36264
rect 4985 36255 5043 36261
rect 5258 36252 5264 36264
rect 5316 36252 5322 36304
rect 5445 36227 5503 36233
rect 5445 36193 5457 36227
rect 5491 36224 5503 36227
rect 6917 36227 6975 36233
rect 6917 36224 6929 36227
rect 5491 36196 6929 36224
rect 5491 36193 5503 36196
rect 5445 36187 5503 36193
rect 6917 36193 6929 36196
rect 6963 36224 6975 36227
rect 8386 36224 8392 36236
rect 6963 36196 8392 36224
rect 6963 36193 6975 36196
rect 6917 36187 6975 36193
rect 5169 36159 5227 36165
rect 5169 36156 5181 36159
rect 4908 36128 5181 36156
rect 4709 36119 4767 36125
rect 5169 36125 5181 36128
rect 5215 36125 5227 36159
rect 5169 36119 5227 36125
rect 5353 36159 5411 36165
rect 5353 36125 5365 36159
rect 5399 36156 5411 36159
rect 5460 36156 5488 36187
rect 5399 36128 5488 36156
rect 5399 36125 5411 36128
rect 5353 36119 5411 36125
rect 5626 36116 5632 36168
rect 5684 36116 5690 36168
rect 5813 36159 5871 36165
rect 5813 36125 5825 36159
rect 5859 36156 5871 36159
rect 6178 36156 6184 36168
rect 5859 36128 6184 36156
rect 5859 36125 5871 36128
rect 5813 36119 5871 36125
rect 6178 36116 6184 36128
rect 6236 36156 6242 36168
rect 6549 36159 6607 36165
rect 6549 36156 6561 36159
rect 6236 36128 6561 36156
rect 6236 36116 6242 36128
rect 6549 36125 6561 36128
rect 6595 36156 6607 36159
rect 6638 36156 6644 36168
rect 6595 36128 6644 36156
rect 6595 36125 6607 36128
rect 6549 36119 6607 36125
rect 6638 36116 6644 36128
rect 6696 36116 6702 36168
rect 6822 36116 6828 36168
rect 6880 36116 6886 36168
rect 4985 36091 5043 36097
rect 4540 36060 4936 36088
rect 4706 35980 4712 36032
rect 4764 36020 4770 36032
rect 4801 36023 4859 36029
rect 4801 36020 4813 36023
rect 4764 35992 4813 36020
rect 4764 35980 4770 35992
rect 4801 35989 4813 35992
rect 4847 35989 4859 36023
rect 4908 36020 4936 36060
rect 4985 36057 4997 36091
rect 5031 36088 5043 36091
rect 5534 36088 5540 36100
rect 5031 36060 5540 36088
rect 5031 36057 5043 36060
rect 4985 36051 5043 36057
rect 5534 36048 5540 36060
rect 5592 36048 5598 36100
rect 7190 36048 7196 36100
rect 7248 36088 7254 36100
rect 7484 36097 7512 36196
rect 8386 36184 8392 36196
rect 8444 36184 8450 36236
rect 8662 36184 8668 36236
rect 8720 36184 8726 36236
rect 7745 36159 7803 36165
rect 7745 36125 7757 36159
rect 7791 36125 7803 36159
rect 7745 36119 7803 36125
rect 7929 36159 7987 36165
rect 7929 36125 7941 36159
rect 7975 36156 7987 36159
rect 8021 36159 8079 36165
rect 8021 36156 8033 36159
rect 7975 36128 8033 36156
rect 7975 36125 7987 36128
rect 7929 36119 7987 36125
rect 8021 36125 8033 36128
rect 8067 36125 8079 36159
rect 8021 36119 8079 36125
rect 7285 36091 7343 36097
rect 7285 36088 7297 36091
rect 7248 36060 7297 36088
rect 7248 36048 7254 36060
rect 7285 36057 7297 36060
rect 7331 36057 7343 36091
rect 7484 36091 7543 36097
rect 7484 36060 7497 36091
rect 7285 36051 7343 36057
rect 7485 36057 7497 36060
rect 7531 36057 7543 36091
rect 7485 36051 7543 36057
rect 7760 36032 7788 36119
rect 8110 36116 8116 36168
rect 8168 36156 8174 36168
rect 9493 36159 9551 36165
rect 9493 36156 9505 36159
rect 8168 36128 9505 36156
rect 8168 36116 8174 36128
rect 9493 36125 9505 36128
rect 9539 36125 9551 36159
rect 9493 36119 9551 36125
rect 19242 36116 19248 36168
rect 19300 36116 19306 36168
rect 20806 36116 20812 36168
rect 20864 36156 20870 36168
rect 21085 36159 21143 36165
rect 21085 36156 21097 36159
rect 20864 36128 21097 36156
rect 20864 36116 20870 36128
rect 21085 36125 21097 36128
rect 21131 36125 21143 36159
rect 21085 36119 21143 36125
rect 21266 36116 21272 36168
rect 21324 36116 21330 36168
rect 21367 36165 21395 36332
rect 21726 36320 21732 36372
rect 21784 36320 21790 36372
rect 22646 36320 22652 36372
rect 22704 36360 22710 36372
rect 23477 36363 23535 36369
rect 23477 36360 23489 36363
rect 22704 36332 23489 36360
rect 22704 36320 22710 36332
rect 23477 36329 23489 36332
rect 23523 36329 23535 36363
rect 23477 36323 23535 36329
rect 24394 36320 24400 36372
rect 24452 36320 24458 36372
rect 24765 36363 24823 36369
rect 24765 36329 24777 36363
rect 24811 36360 24823 36363
rect 25130 36360 25136 36372
rect 24811 36332 25136 36360
rect 24811 36329 24823 36332
rect 24765 36323 24823 36329
rect 25130 36320 25136 36332
rect 25188 36320 25194 36372
rect 27154 36320 27160 36372
rect 27212 36360 27218 36372
rect 27893 36363 27951 36369
rect 27893 36360 27905 36363
rect 27212 36332 27905 36360
rect 27212 36320 27218 36332
rect 27893 36329 27905 36332
rect 27939 36329 27951 36363
rect 27893 36323 27951 36329
rect 28350 36320 28356 36372
rect 28408 36320 28414 36372
rect 28813 36363 28871 36369
rect 28813 36329 28825 36363
rect 28859 36360 28871 36363
rect 29181 36363 29239 36369
rect 29181 36360 29193 36363
rect 28859 36332 29193 36360
rect 28859 36329 28871 36332
rect 28813 36323 28871 36329
rect 29181 36329 29193 36332
rect 29227 36360 29239 36363
rect 29270 36360 29276 36372
rect 29227 36332 29276 36360
rect 29227 36329 29239 36332
rect 29181 36323 29239 36329
rect 29270 36320 29276 36332
rect 29328 36320 29334 36372
rect 29362 36320 29368 36372
rect 29420 36320 29426 36372
rect 22189 36295 22247 36301
rect 22189 36261 22201 36295
rect 22235 36292 22247 36295
rect 22235 36264 22324 36292
rect 22235 36261 22247 36264
rect 22189 36255 22247 36261
rect 21361 36159 21419 36165
rect 21361 36125 21373 36159
rect 21407 36125 21419 36159
rect 21361 36119 21419 36125
rect 21545 36159 21603 36165
rect 21545 36125 21557 36159
rect 21591 36156 21603 36159
rect 21637 36159 21695 36165
rect 21637 36156 21649 36159
rect 21591 36128 21649 36156
rect 21591 36125 21603 36128
rect 21545 36119 21603 36125
rect 21637 36125 21649 36128
rect 21683 36125 21695 36159
rect 21637 36119 21695 36125
rect 22005 36159 22063 36165
rect 22005 36125 22017 36159
rect 22051 36156 22063 36159
rect 22186 36156 22192 36168
rect 22051 36128 22192 36156
rect 22051 36125 22063 36128
rect 22005 36119 22063 36125
rect 19518 36048 19524 36100
rect 19576 36048 19582 36100
rect 19978 36048 19984 36100
rect 20036 36048 20042 36100
rect 21560 36088 21588 36119
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 22296 36165 22324 36264
rect 24044 36264 24900 36292
rect 23658 36184 23664 36236
rect 23716 36224 23722 36236
rect 24044 36233 24072 36264
rect 24029 36227 24087 36233
rect 23716 36196 23888 36224
rect 23716 36184 23722 36196
rect 22281 36159 22339 36165
rect 22281 36125 22293 36159
rect 22327 36156 22339 36159
rect 22370 36156 22376 36168
rect 22327 36128 22376 36156
rect 22327 36125 22339 36128
rect 22281 36119 22339 36125
rect 22370 36116 22376 36128
rect 22428 36116 22434 36168
rect 22465 36159 22523 36165
rect 22465 36125 22477 36159
rect 22511 36125 22523 36159
rect 22465 36119 22523 36125
rect 22833 36159 22891 36165
rect 22833 36125 22845 36159
rect 22879 36156 22891 36159
rect 23750 36156 23756 36168
rect 22879 36128 23756 36156
rect 22879 36125 22891 36128
rect 22833 36119 22891 36125
rect 22480 36088 22508 36119
rect 23750 36116 23756 36128
rect 23808 36116 23814 36168
rect 23860 36165 23888 36196
rect 24029 36193 24041 36227
rect 24075 36193 24087 36227
rect 24762 36224 24768 36236
rect 24029 36187 24087 36193
rect 24136 36196 24768 36224
rect 24136 36168 24164 36196
rect 24762 36184 24768 36196
rect 24820 36184 24826 36236
rect 24872 36224 24900 36264
rect 27614 36252 27620 36304
rect 27672 36292 27678 36304
rect 27672 36264 30512 36292
rect 27672 36252 27678 36264
rect 25038 36224 25044 36236
rect 24872 36196 25044 36224
rect 25038 36184 25044 36196
rect 25096 36224 25102 36236
rect 25317 36227 25375 36233
rect 25317 36224 25329 36227
rect 25096 36196 25329 36224
rect 25096 36184 25102 36196
rect 25317 36193 25329 36196
rect 25363 36193 25375 36227
rect 25317 36187 25375 36193
rect 25961 36227 26019 36233
rect 25961 36193 25973 36227
rect 26007 36224 26019 36227
rect 26602 36224 26608 36236
rect 26007 36196 26608 36224
rect 26007 36193 26019 36196
rect 25961 36187 26019 36193
rect 23845 36159 23903 36165
rect 23845 36125 23857 36159
rect 23891 36156 23903 36159
rect 24118 36156 24124 36168
rect 23891 36128 24124 36156
rect 23891 36125 23903 36128
rect 23845 36119 23903 36125
rect 24118 36116 24124 36128
rect 24176 36116 24182 36168
rect 24210 36116 24216 36168
rect 24268 36156 24274 36168
rect 24397 36159 24455 36165
rect 24397 36156 24409 36159
rect 24268 36128 24409 36156
rect 24268 36116 24274 36128
rect 24397 36125 24409 36128
rect 24443 36125 24455 36159
rect 24581 36159 24639 36165
rect 24581 36156 24593 36159
rect 24397 36119 24455 36125
rect 24504 36128 24593 36156
rect 21008 36060 22508 36088
rect 23937 36091 23995 36097
rect 21008 36032 21036 36060
rect 23937 36057 23949 36091
rect 23983 36088 23995 36091
rect 24504 36088 24532 36128
rect 24581 36125 24593 36128
rect 24627 36156 24639 36159
rect 25133 36159 25191 36165
rect 24627 36128 25085 36156
rect 24627 36125 24639 36128
rect 24581 36119 24639 36125
rect 23983 36060 24532 36088
rect 25057 36088 25085 36128
rect 25133 36125 25145 36159
rect 25179 36156 25191 36159
rect 25976 36156 26004 36187
rect 26602 36184 26608 36196
rect 26660 36184 26666 36236
rect 30484 36233 30512 36264
rect 30469 36227 30527 36233
rect 28736 36196 30144 36224
rect 25179 36128 26004 36156
rect 25179 36125 25191 36128
rect 25133 36119 25191 36125
rect 26142 36116 26148 36168
rect 26200 36156 26206 36168
rect 28736 36165 28764 36196
rect 30116 36168 30144 36196
rect 30469 36193 30481 36227
rect 30515 36193 30527 36227
rect 30469 36187 30527 36193
rect 28077 36159 28135 36165
rect 28077 36156 28089 36159
rect 26200 36128 26245 36156
rect 27632 36128 28089 36156
rect 26200 36116 26206 36128
rect 27632 36100 27660 36128
rect 28077 36125 28089 36128
rect 28123 36125 28135 36159
rect 28077 36119 28135 36125
rect 28353 36159 28411 36165
rect 28353 36125 28365 36159
rect 28399 36125 28411 36159
rect 28353 36119 28411 36125
rect 28537 36159 28595 36165
rect 28537 36125 28549 36159
rect 28583 36125 28595 36159
rect 28537 36119 28595 36125
rect 28721 36159 28779 36165
rect 28721 36125 28733 36159
rect 28767 36125 28779 36159
rect 28721 36119 28779 36125
rect 28905 36159 28963 36165
rect 28905 36125 28917 36159
rect 28951 36156 28963 36159
rect 29454 36156 29460 36168
rect 28951 36128 29460 36156
rect 28951 36125 28963 36128
rect 28905 36119 28963 36125
rect 26329 36091 26387 36097
rect 26329 36088 26341 36091
rect 25057 36060 26341 36088
rect 23983 36057 23995 36060
rect 23937 36051 23995 36057
rect 26329 36057 26341 36060
rect 26375 36088 26387 36091
rect 26970 36088 26976 36100
rect 26375 36060 26976 36088
rect 26375 36057 26387 36060
rect 26329 36051 26387 36057
rect 26970 36048 26976 36060
rect 27028 36088 27034 36100
rect 27028 36060 27568 36088
rect 27028 36048 27034 36060
rect 5905 36023 5963 36029
rect 5905 36020 5917 36023
rect 4908 35992 5917 36020
rect 4801 35983 4859 35989
rect 5905 35989 5917 35992
rect 5951 35989 5963 36023
rect 5905 35983 5963 35989
rect 7653 36023 7711 36029
rect 7653 35989 7665 36023
rect 7699 36020 7711 36023
rect 7742 36020 7748 36032
rect 7699 35992 7748 36020
rect 7699 35989 7711 35992
rect 7653 35983 7711 35989
rect 7742 35980 7748 35992
rect 7800 35980 7806 36032
rect 7834 35980 7840 36032
rect 7892 35980 7898 36032
rect 20990 35980 20996 36032
rect 21048 35980 21054 36032
rect 21450 35980 21456 36032
rect 21508 35980 21514 36032
rect 22278 35980 22284 36032
rect 22336 36020 22342 36032
rect 22465 36023 22523 36029
rect 22465 36020 22477 36023
rect 22336 35992 22477 36020
rect 22336 35980 22342 35992
rect 22465 35989 22477 35992
rect 22511 35989 22523 36023
rect 22465 35983 22523 35989
rect 25222 35980 25228 36032
rect 25280 35980 25286 36032
rect 27338 35980 27344 36032
rect 27396 36020 27402 36032
rect 27433 36023 27491 36029
rect 27433 36020 27445 36023
rect 27396 35992 27445 36020
rect 27396 35980 27402 35992
rect 27433 35989 27445 35992
rect 27479 35989 27491 36023
rect 27540 36020 27568 36060
rect 27614 36048 27620 36100
rect 27672 36048 27678 36100
rect 27798 36048 27804 36100
rect 27856 36048 27862 36100
rect 28166 36048 28172 36100
rect 28224 36088 28230 36100
rect 28261 36091 28319 36097
rect 28261 36088 28273 36091
rect 28224 36060 28273 36088
rect 28224 36048 28230 36060
rect 28261 36057 28273 36060
rect 28307 36088 28319 36091
rect 28368 36088 28396 36119
rect 28307 36060 28396 36088
rect 28552 36088 28580 36119
rect 29454 36116 29460 36128
rect 29512 36116 29518 36168
rect 30098 36116 30104 36168
rect 30156 36116 30162 36168
rect 31846 36116 31852 36168
rect 31904 36116 31910 36168
rect 28552 36060 28948 36088
rect 28307 36057 28319 36060
rect 28261 36051 28319 36057
rect 28810 36020 28816 36032
rect 27540 35992 28816 36020
rect 27433 35983 27491 35989
rect 28810 35980 28816 35992
rect 28868 35980 28874 36032
rect 28920 36020 28948 36060
rect 28994 36048 29000 36100
rect 29052 36048 29058 36100
rect 29549 36091 29607 36097
rect 29549 36088 29561 36091
rect 29104 36060 29561 36088
rect 29104 36020 29132 36060
rect 29549 36057 29561 36060
rect 29595 36057 29607 36091
rect 29549 36051 29607 36057
rect 30742 36048 30748 36100
rect 30800 36048 30806 36100
rect 38470 36048 38476 36100
rect 38528 36048 38534 36100
rect 28920 35992 29132 36020
rect 29178 35980 29184 36032
rect 29236 36029 29242 36032
rect 29236 36023 29255 36029
rect 29243 35989 29255 36023
rect 29236 35983 29255 35989
rect 29236 35980 29242 35983
rect 32214 35980 32220 36032
rect 32272 35980 32278 36032
rect 1104 35930 38824 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 38824 35930
rect 1104 35856 38824 35878
rect 4430 35776 4436 35828
rect 4488 35816 4494 35828
rect 5442 35816 5448 35828
rect 4488 35788 5448 35816
rect 4488 35776 4494 35788
rect 5442 35776 5448 35788
rect 5500 35776 5506 35828
rect 5534 35776 5540 35828
rect 5592 35776 5598 35828
rect 7208 35788 7972 35816
rect 7208 35748 7236 35788
rect 7282 35748 7288 35760
rect 7208 35720 7288 35748
rect 7282 35708 7288 35720
rect 7340 35708 7346 35760
rect 5258 35640 5264 35692
rect 5316 35640 5322 35692
rect 6546 35640 6552 35692
rect 6604 35640 6610 35692
rect 7944 35680 7972 35788
rect 8110 35776 8116 35828
rect 8168 35816 8174 35828
rect 8297 35819 8355 35825
rect 8297 35816 8309 35819
rect 8168 35788 8309 35816
rect 8168 35776 8174 35788
rect 8297 35785 8309 35788
rect 8343 35785 8355 35819
rect 8297 35779 8355 35785
rect 19429 35819 19487 35825
rect 19429 35785 19441 35819
rect 19475 35816 19487 35819
rect 19518 35816 19524 35828
rect 19475 35788 19524 35816
rect 19475 35785 19487 35788
rect 19429 35779 19487 35785
rect 19518 35776 19524 35788
rect 19576 35776 19582 35828
rect 23750 35776 23756 35828
rect 23808 35776 23814 35828
rect 23952 35788 24716 35816
rect 20717 35751 20775 35757
rect 20717 35717 20729 35751
rect 20763 35748 20775 35751
rect 21818 35748 21824 35760
rect 20763 35720 21824 35748
rect 20763 35717 20775 35720
rect 20717 35711 20775 35717
rect 21818 35708 21824 35720
rect 21876 35708 21882 35760
rect 8754 35680 8760 35692
rect 7944 35666 8760 35680
rect 7958 35652 8760 35666
rect 8754 35640 8760 35652
rect 8812 35640 8818 35692
rect 13078 35640 13084 35692
rect 13136 35640 13142 35692
rect 19426 35640 19432 35692
rect 19484 35680 19490 35692
rect 19613 35683 19671 35689
rect 19613 35680 19625 35683
rect 19484 35652 19625 35680
rect 19484 35640 19490 35652
rect 19613 35649 19625 35652
rect 19659 35649 19671 35683
rect 19613 35643 19671 35649
rect 842 35572 848 35624
rect 900 35612 906 35624
rect 1397 35615 1455 35621
rect 1397 35612 1409 35615
rect 900 35584 1409 35612
rect 900 35572 906 35584
rect 1397 35581 1409 35584
rect 1443 35581 1455 35615
rect 1397 35575 1455 35581
rect 4525 35615 4583 35621
rect 4525 35581 4537 35615
rect 4571 35612 4583 35615
rect 4706 35612 4712 35624
rect 4571 35584 4712 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 4706 35572 4712 35584
rect 4764 35572 4770 35624
rect 6086 35572 6092 35624
rect 6144 35572 6150 35624
rect 6825 35615 6883 35621
rect 6825 35581 6837 35615
rect 6871 35612 6883 35615
rect 7834 35612 7840 35624
rect 6871 35584 7840 35612
rect 6871 35581 6883 35584
rect 6825 35575 6883 35581
rect 7834 35572 7840 35584
rect 7892 35572 7898 35624
rect 8018 35572 8024 35624
rect 8076 35612 8082 35624
rect 9861 35615 9919 35621
rect 9861 35612 9873 35615
rect 8076 35584 9873 35612
rect 8076 35572 8082 35584
rect 9861 35581 9873 35584
rect 9907 35581 9919 35615
rect 9861 35575 9919 35581
rect 10137 35615 10195 35621
rect 10137 35581 10149 35615
rect 10183 35612 10195 35615
rect 11054 35612 11060 35624
rect 10183 35584 11060 35612
rect 10183 35581 10195 35584
rect 10137 35575 10195 35581
rect 11054 35572 11060 35584
rect 11112 35572 11118 35624
rect 13357 35615 13415 35621
rect 13357 35581 13369 35615
rect 13403 35612 13415 35615
rect 13630 35612 13636 35624
rect 13403 35584 13636 35612
rect 13403 35581 13415 35584
rect 13357 35575 13415 35581
rect 13630 35572 13636 35584
rect 13688 35572 13694 35624
rect 10870 35504 10876 35556
rect 10928 35544 10934 35556
rect 13173 35547 13231 35553
rect 13173 35544 13185 35547
rect 10928 35516 13185 35544
rect 10928 35504 10934 35516
rect 13173 35513 13185 35516
rect 13219 35513 13231 35547
rect 19628 35544 19656 35643
rect 20070 35640 20076 35692
rect 20128 35680 20134 35692
rect 20165 35683 20223 35689
rect 20165 35680 20177 35683
rect 20128 35652 20177 35680
rect 20128 35640 20134 35652
rect 20165 35649 20177 35652
rect 20211 35649 20223 35683
rect 21450 35680 21456 35692
rect 20165 35643 20223 35649
rect 20272 35652 21456 35680
rect 19889 35615 19947 35621
rect 19889 35581 19901 35615
rect 19935 35612 19947 35615
rect 20272 35612 20300 35652
rect 21450 35640 21456 35652
rect 21508 35640 21514 35692
rect 23658 35640 23664 35692
rect 23716 35640 23722 35692
rect 23842 35640 23848 35692
rect 23900 35680 23906 35692
rect 23952 35689 23980 35788
rect 24026 35708 24032 35760
rect 24084 35748 24090 35760
rect 24581 35751 24639 35757
rect 24581 35748 24593 35751
rect 24084 35720 24593 35748
rect 24084 35708 24090 35720
rect 24581 35717 24593 35720
rect 24627 35717 24639 35751
rect 24581 35711 24639 35717
rect 24688 35748 24716 35788
rect 24762 35776 24768 35828
rect 24820 35816 24826 35828
rect 24820 35788 25084 35816
rect 24820 35776 24826 35788
rect 24949 35751 25007 35757
rect 24949 35748 24961 35751
rect 24688 35720 24961 35748
rect 23937 35683 23995 35689
rect 23937 35680 23949 35683
rect 23900 35652 23949 35680
rect 23900 35640 23906 35652
rect 23937 35649 23949 35652
rect 23983 35649 23995 35683
rect 23937 35643 23995 35649
rect 24121 35683 24179 35689
rect 24121 35649 24133 35683
rect 24167 35649 24179 35683
rect 24121 35643 24179 35649
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 24489 35683 24547 35689
rect 24489 35649 24501 35683
rect 24535 35680 24547 35683
rect 24688 35680 24716 35720
rect 24949 35717 24961 35720
rect 24995 35717 25007 35751
rect 25056 35748 25084 35788
rect 25222 35776 25228 35828
rect 25280 35816 25286 35828
rect 25317 35819 25375 35825
rect 25317 35816 25329 35819
rect 25280 35788 25329 35816
rect 25280 35776 25286 35788
rect 25317 35785 25329 35788
rect 25363 35785 25375 35819
rect 25317 35779 25375 35785
rect 29178 35776 29184 35828
rect 29236 35816 29242 35828
rect 29549 35819 29607 35825
rect 29549 35816 29561 35819
rect 29236 35788 29561 35816
rect 29236 35776 29242 35788
rect 29549 35785 29561 35788
rect 29595 35785 29607 35819
rect 29549 35779 29607 35785
rect 30561 35819 30619 35825
rect 30561 35785 30573 35819
rect 30607 35816 30619 35819
rect 30742 35816 30748 35828
rect 30607 35788 30748 35816
rect 30607 35785 30619 35788
rect 30561 35779 30619 35785
rect 30742 35776 30748 35788
rect 30800 35776 30806 35828
rect 25869 35751 25927 35757
rect 25869 35748 25881 35751
rect 25056 35720 25881 35748
rect 24949 35711 25007 35717
rect 25869 35717 25881 35720
rect 25915 35717 25927 35751
rect 27522 35748 27528 35760
rect 25869 35711 25927 35717
rect 26988 35720 27528 35748
rect 24535 35652 24716 35680
rect 24535 35649 24547 35652
rect 24489 35643 24547 35649
rect 19935 35584 20300 35612
rect 20349 35615 20407 35621
rect 19935 35581 19947 35584
rect 19889 35575 19947 35581
rect 20349 35581 20361 35615
rect 20395 35612 20407 35615
rect 20990 35612 20996 35624
rect 20395 35584 20996 35612
rect 20395 35581 20407 35584
rect 20349 35575 20407 35581
rect 20990 35572 20996 35584
rect 21048 35572 21054 35624
rect 20438 35544 20444 35556
rect 19628 35516 20444 35544
rect 13173 35507 13231 35513
rect 20438 35504 20444 35516
rect 20496 35544 20502 35556
rect 21085 35547 21143 35553
rect 20496 35516 20760 35544
rect 20496 35504 20502 35516
rect 3234 35436 3240 35488
rect 3292 35476 3298 35488
rect 3881 35479 3939 35485
rect 3881 35476 3893 35479
rect 3292 35448 3893 35476
rect 3292 35436 3298 35448
rect 3881 35445 3893 35448
rect 3927 35445 3939 35479
rect 3881 35439 3939 35445
rect 4614 35436 4620 35488
rect 4672 35436 4678 35488
rect 8386 35436 8392 35488
rect 8444 35436 8450 35488
rect 12434 35436 12440 35488
rect 12492 35476 12498 35488
rect 13081 35479 13139 35485
rect 13081 35476 13093 35479
rect 12492 35448 13093 35476
rect 12492 35436 12498 35448
rect 13081 35445 13093 35448
rect 13127 35445 13139 35479
rect 13081 35439 13139 35445
rect 19797 35479 19855 35485
rect 19797 35445 19809 35479
rect 19843 35476 19855 35479
rect 19981 35479 20039 35485
rect 19981 35476 19993 35479
rect 19843 35448 19993 35476
rect 19843 35445 19855 35448
rect 19797 35439 19855 35445
rect 19981 35445 19993 35448
rect 20027 35445 20039 35479
rect 19981 35439 20039 35445
rect 20530 35436 20536 35488
rect 20588 35436 20594 35488
rect 20732 35485 20760 35516
rect 21085 35513 21097 35547
rect 21131 35544 21143 35547
rect 21266 35544 21272 35556
rect 21131 35516 21272 35544
rect 21131 35513 21143 35516
rect 21085 35507 21143 35513
rect 21266 35504 21272 35516
rect 21324 35544 21330 35556
rect 21910 35544 21916 35556
rect 21324 35516 21916 35544
rect 21324 35504 21330 35516
rect 21910 35504 21916 35516
rect 21968 35504 21974 35556
rect 24136 35544 24164 35643
rect 24412 35612 24440 35643
rect 24762 35640 24768 35692
rect 24820 35640 24826 35692
rect 24857 35683 24915 35689
rect 24857 35649 24869 35683
rect 24903 35649 24915 35683
rect 24857 35643 24915 35649
rect 24872 35612 24900 35643
rect 25130 35640 25136 35692
rect 25188 35640 25194 35692
rect 26142 35640 26148 35692
rect 26200 35680 26206 35692
rect 26237 35683 26295 35689
rect 26237 35680 26249 35683
rect 26200 35652 26249 35680
rect 26200 35640 26206 35652
rect 26237 35649 26249 35652
rect 26283 35649 26295 35683
rect 26237 35643 26295 35649
rect 26513 35683 26571 35689
rect 26513 35649 26525 35683
rect 26559 35680 26571 35683
rect 26602 35680 26608 35692
rect 26559 35652 26608 35680
rect 26559 35649 26571 35652
rect 26513 35643 26571 35649
rect 25409 35615 25467 35621
rect 25409 35612 25421 35615
rect 24412 35584 25421 35612
rect 25409 35581 25421 35584
rect 25455 35581 25467 35615
rect 25409 35575 25467 35581
rect 25593 35547 25651 35553
rect 25593 35544 25605 35547
rect 24136 35516 25605 35544
rect 25593 35513 25605 35516
rect 25639 35544 25651 35547
rect 26234 35544 26240 35556
rect 25639 35516 26240 35544
rect 25639 35513 25651 35516
rect 25593 35507 25651 35513
rect 26234 35504 26240 35516
rect 26292 35544 26298 35556
rect 26528 35544 26556 35643
rect 26602 35640 26608 35652
rect 26660 35640 26666 35692
rect 26988 35689 27016 35720
rect 27522 35708 27528 35720
rect 27580 35708 27586 35760
rect 27982 35708 27988 35760
rect 28040 35708 28046 35760
rect 29454 35708 29460 35760
rect 29512 35748 29518 35760
rect 29733 35751 29791 35757
rect 29733 35748 29745 35751
rect 29512 35720 29745 35748
rect 29512 35708 29518 35720
rect 29733 35717 29745 35720
rect 29779 35717 29791 35751
rect 29733 35711 29791 35717
rect 30377 35751 30435 35757
rect 30377 35717 30389 35751
rect 30423 35748 30435 35751
rect 30466 35748 30472 35760
rect 30423 35720 30472 35748
rect 30423 35717 30435 35720
rect 30377 35711 30435 35717
rect 26973 35683 27031 35689
rect 26973 35649 26985 35683
rect 27019 35649 27031 35683
rect 26973 35643 27031 35649
rect 27614 35572 27620 35624
rect 27672 35612 27678 35624
rect 28721 35615 28779 35621
rect 28721 35612 28733 35615
rect 27672 35584 28733 35612
rect 27672 35572 27678 35584
rect 28721 35581 28733 35584
rect 28767 35581 28779 35615
rect 29748 35612 29776 35711
rect 30466 35708 30472 35720
rect 30524 35708 30530 35760
rect 30944 35720 31524 35748
rect 29917 35683 29975 35689
rect 29917 35649 29929 35683
rect 29963 35680 29975 35683
rect 30098 35680 30104 35692
rect 29963 35652 30104 35680
rect 29963 35649 29975 35652
rect 29917 35643 29975 35649
rect 30098 35640 30104 35652
rect 30156 35680 30162 35692
rect 30944 35689 30972 35720
rect 31496 35689 31524 35720
rect 30668 35680 30880 35686
rect 30929 35683 30987 35689
rect 30929 35680 30941 35683
rect 30156 35658 30941 35680
rect 30156 35652 30696 35658
rect 30852 35652 30941 35658
rect 30156 35640 30162 35652
rect 30929 35649 30941 35652
rect 30975 35649 30987 35683
rect 30929 35643 30987 35649
rect 31113 35683 31171 35689
rect 31113 35649 31125 35683
rect 31159 35680 31171 35683
rect 31481 35683 31539 35689
rect 31159 35652 31432 35680
rect 31159 35649 31171 35652
rect 31113 35643 31171 35649
rect 29748 35584 30604 35612
rect 28721 35575 28779 35581
rect 26292 35516 26556 35544
rect 30009 35547 30067 35553
rect 26292 35504 26298 35516
rect 30009 35513 30021 35547
rect 30055 35544 30067 35547
rect 30190 35544 30196 35556
rect 30055 35516 30196 35544
rect 30055 35513 30067 35516
rect 30009 35507 30067 35513
rect 30190 35504 30196 35516
rect 30248 35504 30254 35556
rect 30576 35544 30604 35584
rect 30834 35572 30840 35624
rect 30892 35572 30898 35624
rect 31021 35615 31079 35621
rect 31021 35581 31033 35615
rect 31067 35612 31079 35615
rect 31297 35615 31355 35621
rect 31297 35612 31309 35615
rect 31067 35584 31309 35612
rect 31067 35581 31079 35584
rect 31021 35575 31079 35581
rect 31297 35581 31309 35584
rect 31343 35581 31355 35615
rect 31404 35612 31432 35652
rect 31481 35649 31493 35683
rect 31527 35649 31539 35683
rect 31481 35643 31539 35649
rect 31754 35612 31760 35624
rect 31404 35584 31760 35612
rect 31297 35575 31355 35581
rect 31036 35544 31064 35575
rect 31754 35572 31760 35584
rect 31812 35612 31818 35624
rect 32214 35612 32220 35624
rect 31812 35584 32220 35612
rect 31812 35572 31818 35584
rect 32214 35572 32220 35584
rect 32272 35572 32278 35624
rect 30576 35516 31064 35544
rect 20717 35479 20775 35485
rect 20717 35445 20729 35479
rect 20763 35476 20775 35479
rect 22278 35476 22284 35488
rect 20763 35448 22284 35476
rect 20763 35445 20775 35448
rect 20717 35439 20775 35445
rect 22278 35436 22284 35448
rect 22336 35436 22342 35488
rect 24210 35436 24216 35488
rect 24268 35436 24274 35488
rect 24302 35436 24308 35488
rect 24360 35476 24366 35488
rect 25130 35476 25136 35488
rect 24360 35448 25136 35476
rect 24360 35436 24366 35448
rect 25130 35436 25136 35448
rect 25188 35436 25194 35488
rect 26329 35479 26387 35485
rect 26329 35445 26341 35479
rect 26375 35476 26387 35479
rect 27062 35476 27068 35488
rect 26375 35448 27068 35476
rect 26375 35445 26387 35448
rect 26329 35439 26387 35445
rect 27062 35436 27068 35448
rect 27120 35436 27126 35488
rect 27236 35479 27294 35485
rect 27236 35445 27248 35479
rect 27282 35476 27294 35479
rect 27430 35476 27436 35488
rect 27282 35448 27436 35476
rect 27282 35445 27294 35448
rect 27236 35439 27294 35445
rect 27430 35436 27436 35448
rect 27488 35436 27494 35488
rect 28994 35436 29000 35488
rect 29052 35476 29058 35488
rect 30377 35479 30435 35485
rect 30377 35476 30389 35479
rect 29052 35448 30389 35476
rect 29052 35436 29058 35448
rect 30377 35445 30389 35448
rect 30423 35445 30435 35479
rect 30377 35439 30435 35445
rect 30466 35436 30472 35488
rect 30524 35476 30530 35488
rect 30653 35479 30711 35485
rect 30653 35476 30665 35479
rect 30524 35448 30665 35476
rect 30524 35436 30530 35448
rect 30653 35445 30665 35448
rect 30699 35445 30711 35479
rect 30653 35439 30711 35445
rect 31665 35479 31723 35485
rect 31665 35445 31677 35479
rect 31711 35476 31723 35479
rect 32030 35476 32036 35488
rect 31711 35448 32036 35476
rect 31711 35445 31723 35448
rect 31665 35439 31723 35445
rect 32030 35436 32036 35448
rect 32088 35436 32094 35488
rect 38470 35436 38476 35488
rect 38528 35436 38534 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 3970 35232 3976 35284
rect 4028 35272 4034 35284
rect 5718 35272 5724 35284
rect 4028 35244 5724 35272
rect 4028 35232 4034 35244
rect 5718 35232 5724 35244
rect 5776 35232 5782 35284
rect 6086 35232 6092 35284
rect 6144 35232 6150 35284
rect 7193 35275 7251 35281
rect 7193 35241 7205 35275
rect 7239 35272 7251 35275
rect 7466 35272 7472 35284
rect 7239 35244 7472 35272
rect 7239 35241 7251 35244
rect 7193 35235 7251 35241
rect 7466 35232 7472 35244
rect 7524 35232 7530 35284
rect 8018 35232 8024 35284
rect 8076 35232 8082 35284
rect 10778 35232 10784 35284
rect 10836 35272 10842 35284
rect 12529 35275 12587 35281
rect 10836 35244 12434 35272
rect 10836 35232 10842 35244
rect 8386 35204 8392 35216
rect 6748 35176 8392 35204
rect 2866 35096 2872 35148
rect 2924 35096 2930 35148
rect 3326 35096 3332 35148
rect 3384 35096 3390 35148
rect 4614 35136 4620 35148
rect 4264 35108 4620 35136
rect 842 35028 848 35080
rect 900 35068 906 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 900 35040 1409 35068
rect 900 35028 906 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 3234 35028 3240 35080
rect 3292 35028 3298 35080
rect 4264 35077 4292 35108
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 6748 35145 6776 35176
rect 8386 35164 8392 35176
rect 8444 35204 8450 35216
rect 12406 35204 12434 35244
rect 12529 35241 12541 35275
rect 12575 35272 12587 35275
rect 12710 35272 12716 35284
rect 12575 35244 12716 35272
rect 12575 35241 12587 35244
rect 12529 35235 12587 35241
rect 12710 35232 12716 35244
rect 12768 35232 12774 35284
rect 13078 35232 13084 35284
rect 13136 35272 13142 35284
rect 13725 35275 13783 35281
rect 13725 35272 13737 35275
rect 13136 35244 13737 35272
rect 13136 35232 13142 35244
rect 13725 35241 13737 35244
rect 13771 35241 13783 35275
rect 13725 35235 13783 35241
rect 17034 35232 17040 35284
rect 17092 35272 17098 35284
rect 17773 35275 17831 35281
rect 17773 35272 17785 35275
rect 17092 35244 17785 35272
rect 17092 35232 17098 35244
rect 17773 35241 17785 35244
rect 17819 35241 17831 35275
rect 17773 35235 17831 35241
rect 20530 35232 20536 35284
rect 20588 35272 20594 35284
rect 20698 35275 20756 35281
rect 20698 35272 20710 35275
rect 20588 35244 20710 35272
rect 20588 35232 20594 35244
rect 20698 35241 20710 35244
rect 20744 35241 20756 35275
rect 20698 35235 20756 35241
rect 22186 35232 22192 35284
rect 22244 35232 22250 35284
rect 24213 35275 24271 35281
rect 24213 35241 24225 35275
rect 24259 35272 24271 35275
rect 24302 35272 24308 35284
rect 24259 35244 24308 35272
rect 24259 35241 24271 35244
rect 24213 35235 24271 35241
rect 24302 35232 24308 35244
rect 24360 35232 24366 35284
rect 25225 35275 25283 35281
rect 25225 35272 25237 35275
rect 25056 35244 25237 35272
rect 15289 35207 15347 35213
rect 8444 35176 8708 35204
rect 12406 35176 15148 35204
rect 8444 35164 8450 35176
rect 6733 35139 6791 35145
rect 6733 35105 6745 35139
rect 6779 35105 6791 35139
rect 6733 35099 6791 35105
rect 7742 35096 7748 35148
rect 7800 35096 7806 35148
rect 8680 35145 8708 35176
rect 8665 35139 8723 35145
rect 8665 35105 8677 35139
rect 8711 35105 8723 35139
rect 8665 35099 8723 35105
rect 10781 35139 10839 35145
rect 10781 35105 10793 35139
rect 10827 35136 10839 35139
rect 11054 35136 11060 35148
rect 10827 35108 11060 35136
rect 10827 35105 10839 35108
rect 10781 35099 10839 35105
rect 11054 35096 11060 35108
rect 11112 35096 11118 35148
rect 13538 35136 13544 35148
rect 12176 35108 13544 35136
rect 4065 35071 4123 35077
rect 4065 35037 4077 35071
rect 4111 35037 4123 35071
rect 4065 35031 4123 35037
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35037 4307 35071
rect 4249 35031 4307 35037
rect 4080 34932 4108 35031
rect 4338 35028 4344 35080
rect 4396 35028 4402 35080
rect 5718 35028 5724 35080
rect 5776 35028 5782 35080
rect 6638 35028 6644 35080
rect 6696 35068 6702 35080
rect 6825 35071 6883 35077
rect 6825 35068 6837 35071
rect 6696 35040 6837 35068
rect 6696 35028 6702 35040
rect 6825 35037 6837 35040
rect 6871 35037 6883 35071
rect 6825 35031 6883 35037
rect 7190 35028 7196 35080
rect 7248 35028 7254 35080
rect 7653 35071 7711 35077
rect 7653 35037 7665 35071
rect 7699 35068 7711 35071
rect 8113 35071 8171 35077
rect 8113 35068 8125 35071
rect 7699 35040 8125 35068
rect 7699 35037 7711 35040
rect 7653 35031 7711 35037
rect 8113 35037 8125 35040
rect 8159 35037 8171 35071
rect 12176 35054 12204 35108
rect 13538 35096 13544 35108
rect 13596 35096 13602 35148
rect 8113 35031 8171 35037
rect 12710 35028 12716 35080
rect 12768 35068 12774 35080
rect 13265 35071 13323 35077
rect 13265 35068 13277 35071
rect 12768 35040 13277 35068
rect 12768 35028 12774 35040
rect 13265 35037 13277 35040
rect 13311 35068 13323 35071
rect 13446 35068 13452 35080
rect 13311 35040 13452 35068
rect 13311 35037 13323 35040
rect 13265 35031 13323 35037
rect 13446 35028 13452 35040
rect 13504 35028 13510 35080
rect 13906 35028 13912 35080
rect 13964 35068 13970 35080
rect 15120 35077 15148 35176
rect 15289 35173 15301 35207
rect 15335 35204 15347 35207
rect 15565 35207 15623 35213
rect 15565 35204 15577 35207
rect 15335 35176 15577 35204
rect 15335 35173 15347 35176
rect 15289 35167 15347 35173
rect 15565 35173 15577 35176
rect 15611 35204 15623 35207
rect 16298 35204 16304 35216
rect 15611 35176 16304 35204
rect 15611 35173 15623 35176
rect 15565 35167 15623 35173
rect 16298 35164 16304 35176
rect 16356 35204 16362 35216
rect 18233 35207 18291 35213
rect 18233 35204 18245 35207
rect 16356 35176 18245 35204
rect 16356 35164 16362 35176
rect 18233 35173 18245 35176
rect 18279 35173 18291 35207
rect 18233 35167 18291 35173
rect 24026 35164 24032 35216
rect 24084 35204 24090 35216
rect 24084 35176 24808 35204
rect 24084 35164 24090 35176
rect 15933 35139 15991 35145
rect 15933 35136 15945 35139
rect 15212 35108 15945 35136
rect 14645 35071 14703 35077
rect 14645 35068 14657 35071
rect 13964 35040 14657 35068
rect 13964 35028 13970 35040
rect 14645 35037 14657 35040
rect 14691 35037 14703 35071
rect 14645 35031 14703 35037
rect 15105 35071 15163 35077
rect 15105 35037 15117 35071
rect 15151 35037 15163 35071
rect 15105 35031 15163 35037
rect 4157 35003 4215 35009
rect 4157 34969 4169 35003
rect 4203 35000 4215 35003
rect 4617 35003 4675 35009
rect 4617 35000 4629 35003
rect 4203 34972 4629 35000
rect 4203 34969 4215 34972
rect 4157 34963 4215 34969
rect 4617 34969 4629 34972
rect 4663 34969 4675 35003
rect 4617 34963 4675 34969
rect 10962 34960 10968 35012
rect 11020 35000 11026 35012
rect 11057 35003 11115 35009
rect 11057 35000 11069 35003
rect 11020 34972 11069 35000
rect 11020 34960 11026 34972
rect 11057 34969 11069 34972
rect 11103 34969 11115 35003
rect 11057 34963 11115 34969
rect 13725 35003 13783 35009
rect 13725 34969 13737 35003
rect 13771 35000 13783 35003
rect 14093 35003 14151 35009
rect 14093 35000 14105 35003
rect 13771 34972 14105 35000
rect 13771 34969 13783 34972
rect 13725 34963 13783 34969
rect 14093 34969 14105 34972
rect 14139 34969 14151 35003
rect 14093 34963 14151 34969
rect 15010 34960 15016 35012
rect 15068 35000 15074 35012
rect 15212 35000 15240 35108
rect 15933 35105 15945 35108
rect 15979 35105 15991 35139
rect 15933 35099 15991 35105
rect 20441 35139 20499 35145
rect 20441 35105 20453 35139
rect 20487 35136 20499 35139
rect 22186 35136 22192 35148
rect 20487 35108 22192 35136
rect 20487 35105 20499 35108
rect 20441 35099 20499 35105
rect 22186 35096 22192 35108
rect 22244 35096 22250 35148
rect 22925 35139 22983 35145
rect 22925 35105 22937 35139
rect 22971 35136 22983 35139
rect 24210 35136 24216 35148
rect 22971 35108 24216 35136
rect 22971 35105 22983 35108
rect 22925 35099 22983 35105
rect 24210 35096 24216 35108
rect 24268 35096 24274 35148
rect 24780 35136 24808 35176
rect 24857 35139 24915 35145
rect 24857 35136 24869 35139
rect 24780 35108 24869 35136
rect 24857 35105 24869 35108
rect 24903 35105 24915 35139
rect 24857 35099 24915 35105
rect 24946 35096 24952 35148
rect 25004 35096 25010 35148
rect 15654 35028 15660 35080
rect 15712 35028 15718 35080
rect 17494 35028 17500 35080
rect 17552 35068 17558 35080
rect 18049 35071 18107 35077
rect 18049 35068 18061 35071
rect 17552 35040 18061 35068
rect 17552 35028 17558 35040
rect 18049 35037 18061 35040
rect 18095 35037 18107 35071
rect 18049 35031 18107 35037
rect 18322 35028 18328 35080
rect 18380 35028 18386 35080
rect 22370 35028 22376 35080
rect 22428 35068 22434 35080
rect 22649 35071 22707 35077
rect 22649 35068 22661 35071
rect 22428 35040 22661 35068
rect 22428 35028 22434 35040
rect 22649 35037 22661 35040
rect 22695 35037 22707 35071
rect 22649 35031 22707 35037
rect 22741 35071 22799 35077
rect 22741 35037 22753 35071
rect 22787 35068 22799 35071
rect 23290 35068 23296 35080
rect 22787 35040 23296 35068
rect 22787 35037 22799 35040
rect 22741 35031 22799 35037
rect 23290 35028 23296 35040
rect 23348 35028 23354 35080
rect 23658 35028 23664 35080
rect 23716 35068 23722 35080
rect 23753 35071 23811 35077
rect 23753 35068 23765 35071
rect 23716 35040 23765 35068
rect 23716 35028 23722 35040
rect 23753 35037 23765 35040
rect 23799 35037 23811 35071
rect 23753 35031 23811 35037
rect 15068 34972 15240 35000
rect 15068 34960 15074 34972
rect 15286 34960 15292 35012
rect 15344 35000 15350 35012
rect 15381 35003 15439 35009
rect 15381 35000 15393 35003
rect 15344 34972 15393 35000
rect 15344 34960 15350 34972
rect 15381 34969 15393 34972
rect 15427 35000 15439 35003
rect 16114 35000 16120 35012
rect 15427 34972 16120 35000
rect 15427 34969 15439 34972
rect 15381 34963 15439 34969
rect 16114 34960 16120 34972
rect 16172 34960 16178 35012
rect 17402 34960 17408 35012
rect 17460 35000 17466 35012
rect 17957 35003 18015 35009
rect 17957 35000 17969 35003
rect 17460 34972 17969 35000
rect 17460 34960 17466 34972
rect 17957 34969 17969 34972
rect 18003 34969 18015 35003
rect 17957 34963 18015 34969
rect 21358 34960 21364 35012
rect 21416 34960 21422 35012
rect 23768 35000 23796 35031
rect 23842 35028 23848 35080
rect 23900 35068 23906 35080
rect 24765 35071 24823 35077
rect 24765 35068 24777 35071
rect 23900 35040 24777 35068
rect 23900 35028 23906 35040
rect 24765 35037 24777 35040
rect 24811 35068 24823 35071
rect 25056 35068 25084 35244
rect 25225 35241 25237 35244
rect 25271 35241 25283 35275
rect 25225 35235 25283 35241
rect 27246 35232 27252 35284
rect 27304 35232 27310 35284
rect 27430 35232 27436 35284
rect 27488 35232 27494 35284
rect 30834 35232 30840 35284
rect 30892 35272 30898 35284
rect 30929 35275 30987 35281
rect 30929 35272 30941 35275
rect 30892 35244 30941 35272
rect 30892 35232 30898 35244
rect 30929 35241 30941 35244
rect 30975 35272 30987 35275
rect 31202 35272 31208 35284
rect 30975 35244 31208 35272
rect 30975 35241 30987 35244
rect 30929 35235 30987 35241
rect 31202 35232 31208 35244
rect 31260 35272 31266 35284
rect 31941 35275 31999 35281
rect 31941 35272 31953 35275
rect 31260 35244 31953 35272
rect 31260 35232 31266 35244
rect 31941 35241 31953 35244
rect 31987 35272 31999 35275
rect 32398 35272 32404 35284
rect 31987 35244 32404 35272
rect 31987 35241 31999 35244
rect 31941 35235 31999 35241
rect 32398 35232 32404 35244
rect 32456 35232 32462 35284
rect 26142 35164 26148 35216
rect 26200 35204 26206 35216
rect 28261 35207 28319 35213
rect 28261 35204 28273 35207
rect 26200 35176 28273 35204
rect 26200 35164 26206 35176
rect 28261 35173 28273 35176
rect 28307 35204 28319 35207
rect 28307 35176 30144 35204
rect 28307 35173 28319 35176
rect 28261 35167 28319 35173
rect 30116 35148 30144 35176
rect 30190 35164 30196 35216
rect 30248 35204 30254 35216
rect 30745 35207 30803 35213
rect 30745 35204 30757 35207
rect 30248 35176 30757 35204
rect 30248 35164 30254 35176
rect 30745 35173 30757 35176
rect 30791 35173 30803 35207
rect 32122 35204 32128 35216
rect 30745 35167 30803 35173
rect 30852 35176 32128 35204
rect 26234 35136 26240 35148
rect 25240 35108 26240 35136
rect 25240 35077 25268 35108
rect 26234 35096 26240 35108
rect 26292 35096 26298 35148
rect 27798 35136 27804 35148
rect 27724 35108 27804 35136
rect 24811 35040 25084 35068
rect 25225 35071 25283 35077
rect 24811 35037 24823 35040
rect 24765 35031 24823 35037
rect 25225 35037 25237 35071
rect 25271 35037 25283 35071
rect 25225 35031 25283 35037
rect 25317 35071 25375 35077
rect 25317 35037 25329 35071
rect 25363 35037 25375 35071
rect 25317 35031 25375 35037
rect 25332 35000 25360 35031
rect 27154 35028 27160 35080
rect 27212 35068 27218 35080
rect 27525 35071 27583 35077
rect 27212 35040 27476 35068
rect 27212 35028 27218 35040
rect 23768 34972 25360 35000
rect 26970 34960 26976 35012
rect 27028 35000 27034 35012
rect 27338 35009 27344 35012
rect 27065 35003 27123 35009
rect 27065 35000 27077 35003
rect 27028 34972 27077 35000
rect 27028 34960 27034 34972
rect 27065 34969 27077 34972
rect 27111 34969 27123 35003
rect 27065 34963 27123 34969
rect 27281 35003 27344 35009
rect 27281 34969 27293 35003
rect 27327 34969 27344 35003
rect 27281 34963 27344 34969
rect 27338 34960 27344 34963
rect 27396 34960 27402 35012
rect 27448 35000 27476 35040
rect 27525 35037 27537 35071
rect 27571 35068 27583 35071
rect 27614 35068 27620 35080
rect 27571 35040 27620 35068
rect 27571 35037 27583 35040
rect 27525 35031 27583 35037
rect 27614 35028 27620 35040
rect 27672 35028 27678 35080
rect 27724 35077 27752 35108
rect 27798 35096 27804 35108
rect 27856 35136 27862 35148
rect 29641 35139 29699 35145
rect 29641 35136 29653 35139
rect 27856 35108 29653 35136
rect 27856 35096 27862 35108
rect 28276 35077 28304 35108
rect 29641 35105 29653 35108
rect 29687 35105 29699 35139
rect 29641 35099 29699 35105
rect 30098 35096 30104 35148
rect 30156 35136 30162 35148
rect 30852 35136 30880 35176
rect 32122 35164 32128 35176
rect 32180 35164 32186 35216
rect 32030 35136 32036 35148
rect 30156 35108 30880 35136
rect 31036 35108 32036 35136
rect 30156 35096 30162 35108
rect 27709 35071 27767 35077
rect 27709 35037 27721 35071
rect 27755 35037 27767 35071
rect 27709 35031 27767 35037
rect 28077 35071 28135 35077
rect 28077 35037 28089 35071
rect 28123 35037 28135 35071
rect 28077 35031 28135 35037
rect 28261 35071 28319 35077
rect 28261 35037 28273 35071
rect 28307 35037 28319 35071
rect 28261 35031 28319 35037
rect 28092 35000 28120 35031
rect 29270 35028 29276 35080
rect 29328 35068 29334 35080
rect 29549 35071 29607 35077
rect 29549 35068 29561 35071
rect 29328 35040 29561 35068
rect 29328 35028 29334 35040
rect 29549 35037 29561 35040
rect 29595 35037 29607 35071
rect 29549 35031 29607 35037
rect 29730 35028 29736 35080
rect 29788 35028 29794 35080
rect 30190 35028 30196 35080
rect 30248 35028 30254 35080
rect 30377 35071 30435 35077
rect 30377 35037 30389 35071
rect 30423 35068 30435 35071
rect 30650 35068 30656 35080
rect 30423 35040 30656 35068
rect 30423 35037 30435 35040
rect 30377 35031 30435 35037
rect 28166 35000 28172 35012
rect 27448 34972 28172 35000
rect 28166 34960 28172 34972
rect 28224 35000 28230 35012
rect 28718 35000 28724 35012
rect 28224 34972 28724 35000
rect 28224 34960 28230 34972
rect 28718 34960 28724 34972
rect 28776 34960 28782 35012
rect 29914 34960 29920 35012
rect 29972 35000 29978 35012
rect 30392 35000 30420 35031
rect 30650 35028 30656 35040
rect 30708 35028 30714 35080
rect 29972 34972 30420 35000
rect 30913 35003 30971 35009
rect 29972 34960 29978 34972
rect 30913 34969 30925 35003
rect 30959 35000 30971 35003
rect 31036 35000 31064 35108
rect 32030 35096 32036 35108
rect 32088 35096 32094 35148
rect 33318 35096 33324 35148
rect 33376 35136 33382 35148
rect 33689 35139 33747 35145
rect 33689 35136 33701 35139
rect 33376 35108 33701 35136
rect 33376 35096 33382 35108
rect 33689 35105 33701 35108
rect 33735 35105 33747 35139
rect 33689 35099 33747 35105
rect 31202 35028 31208 35080
rect 31260 35028 31266 35080
rect 31846 35028 31852 35080
rect 31904 35068 31910 35080
rect 31904 35040 32338 35068
rect 31904 35028 31910 35040
rect 30959 34972 31064 35000
rect 31113 35003 31171 35009
rect 30959 34969 30971 34972
rect 30913 34963 30971 34969
rect 31113 34969 31125 35003
rect 31159 35000 31171 35003
rect 31754 35000 31760 35012
rect 31159 34972 31760 35000
rect 31159 34969 31171 34972
rect 31113 34963 31171 34969
rect 5258 34932 5264 34944
rect 4080 34904 5264 34932
rect 5258 34892 5264 34904
rect 5316 34892 5322 34944
rect 7374 34892 7380 34944
rect 7432 34892 7438 34944
rect 11698 34892 11704 34944
rect 11756 34932 11762 34944
rect 12621 34935 12679 34941
rect 12621 34932 12633 34935
rect 11756 34904 12633 34932
rect 11756 34892 11762 34904
rect 12621 34901 12633 34904
rect 12667 34901 12679 34935
rect 12621 34895 12679 34901
rect 13078 34892 13084 34944
rect 13136 34932 13142 34944
rect 13541 34935 13599 34941
rect 13541 34932 13553 34935
rect 13136 34904 13553 34932
rect 13136 34892 13142 34904
rect 13541 34901 13553 34904
rect 13587 34901 13599 34935
rect 13541 34895 13599 34901
rect 15470 34892 15476 34944
rect 15528 34932 15534 34944
rect 15657 34935 15715 34941
rect 15657 34932 15669 34935
rect 15528 34904 15669 34932
rect 15528 34892 15534 34904
rect 15657 34901 15669 34904
rect 15703 34901 15715 34935
rect 15657 34895 15715 34901
rect 16022 34892 16028 34944
rect 16080 34932 16086 34944
rect 16577 34935 16635 34941
rect 16577 34932 16589 34935
rect 16080 34904 16589 34932
rect 16080 34892 16086 34904
rect 16577 34901 16589 34904
rect 16623 34901 16635 34935
rect 16577 34895 16635 34901
rect 17494 34892 17500 34944
rect 17552 34932 17558 34944
rect 17589 34935 17647 34941
rect 17589 34932 17601 34935
rect 17552 34904 17601 34932
rect 17552 34892 17558 34904
rect 17589 34901 17601 34904
rect 17635 34901 17647 34935
rect 17589 34895 17647 34901
rect 17757 34935 17815 34941
rect 17757 34901 17769 34935
rect 17803 34932 17815 34935
rect 17862 34932 17868 34944
rect 17803 34904 17868 34932
rect 17803 34901 17815 34904
rect 17757 34895 17815 34901
rect 17862 34892 17868 34904
rect 17920 34892 17926 34944
rect 18325 34935 18383 34941
rect 18325 34901 18337 34935
rect 18371 34932 18383 34935
rect 18874 34932 18880 34944
rect 18371 34904 18880 34932
rect 18371 34901 18383 34904
rect 18325 34895 18383 34901
rect 18874 34892 18880 34904
rect 18932 34892 18938 34944
rect 22922 34892 22928 34944
rect 22980 34892 22986 34944
rect 24397 34935 24455 34941
rect 24397 34901 24409 34935
rect 24443 34932 24455 34935
rect 24578 34932 24584 34944
rect 24443 34904 24584 34932
rect 24443 34901 24455 34904
rect 24397 34895 24455 34901
rect 24578 34892 24584 34904
rect 24636 34892 24642 34944
rect 25222 34892 25228 34944
rect 25280 34932 25286 34944
rect 25593 34935 25651 34941
rect 25593 34932 25605 34935
rect 25280 34904 25605 34932
rect 25280 34892 25286 34904
rect 25593 34901 25605 34904
rect 25639 34901 25651 34935
rect 25593 34895 25651 34901
rect 27430 34892 27436 34944
rect 27488 34932 27494 34944
rect 27525 34935 27583 34941
rect 27525 34932 27537 34935
rect 27488 34904 27537 34932
rect 27488 34892 27494 34904
rect 27525 34901 27537 34904
rect 27571 34901 27583 34935
rect 27525 34895 27583 34901
rect 30374 34892 30380 34944
rect 30432 34892 30438 34944
rect 31018 34892 31024 34944
rect 31076 34932 31082 34944
rect 31128 34932 31156 34963
rect 31754 34960 31760 34972
rect 31812 34960 31818 35012
rect 33413 35003 33471 35009
rect 33413 34969 33425 35003
rect 33459 34969 33471 35003
rect 33413 34963 33471 34969
rect 31076 34904 31156 34932
rect 31076 34892 31082 34904
rect 31662 34892 31668 34944
rect 31720 34932 31726 34944
rect 31849 34935 31907 34941
rect 31849 34932 31861 34935
rect 31720 34904 31861 34932
rect 31720 34892 31726 34904
rect 31849 34901 31861 34904
rect 31895 34901 31907 34935
rect 31849 34895 31907 34901
rect 31938 34892 31944 34944
rect 31996 34932 32002 34944
rect 33428 34932 33456 34963
rect 31996 34904 33456 34932
rect 31996 34892 32002 34904
rect 38470 34892 38476 34944
rect 38528 34892 38534 34944
rect 1104 34842 38824 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 38824 34842
rect 1104 34768 38824 34790
rect 3878 34728 3884 34740
rect 2608 34700 3884 34728
rect 2222 34484 2228 34536
rect 2280 34524 2286 34536
rect 2608 34533 2636 34700
rect 3878 34688 3884 34700
rect 3936 34728 3942 34740
rect 3936 34700 4384 34728
rect 3936 34688 3942 34700
rect 4356 34672 4384 34700
rect 10962 34688 10968 34740
rect 11020 34688 11026 34740
rect 12618 34728 12624 34740
rect 11808 34700 12624 34728
rect 2866 34620 2872 34672
rect 2924 34620 2930 34672
rect 4338 34620 4344 34672
rect 4396 34660 4402 34672
rect 4617 34663 4675 34669
rect 4617 34660 4629 34663
rect 4396 34632 4629 34660
rect 4396 34620 4402 34632
rect 4617 34629 4629 34632
rect 4663 34660 4675 34663
rect 11698 34660 11704 34672
rect 4663 34632 5948 34660
rect 4663 34629 4675 34632
rect 4617 34623 4675 34629
rect 3970 34552 3976 34604
rect 4028 34552 4034 34604
rect 5920 34601 5948 34632
rect 11072 34632 11704 34660
rect 5353 34595 5411 34601
rect 5353 34561 5365 34595
rect 5399 34561 5411 34595
rect 5353 34555 5411 34561
rect 5905 34595 5963 34601
rect 5905 34561 5917 34595
rect 5951 34592 5963 34595
rect 6546 34592 6552 34604
rect 5951 34564 6552 34592
rect 5951 34561 5963 34564
rect 5905 34555 5963 34561
rect 2593 34527 2651 34533
rect 2593 34524 2605 34527
rect 2280 34496 2605 34524
rect 2280 34484 2286 34496
rect 2593 34493 2605 34496
rect 2639 34493 2651 34527
rect 5368 34524 5396 34555
rect 6546 34552 6552 34564
rect 6604 34552 6610 34604
rect 9766 34552 9772 34604
rect 9824 34552 9830 34604
rect 10137 34595 10195 34601
rect 10137 34561 10149 34595
rect 10183 34561 10195 34595
rect 10137 34555 10195 34561
rect 6181 34527 6239 34533
rect 6181 34524 6193 34527
rect 5368 34496 6193 34524
rect 2593 34487 2651 34493
rect 6181 34493 6193 34496
rect 6227 34524 6239 34527
rect 6362 34524 6368 34536
rect 6227 34496 6368 34524
rect 6227 34493 6239 34496
rect 6181 34487 6239 34493
rect 6362 34484 6368 34496
rect 6420 34484 6426 34536
rect 9214 34484 9220 34536
rect 9272 34524 9278 34536
rect 9585 34527 9643 34533
rect 9585 34524 9597 34527
rect 9272 34496 9597 34524
rect 9272 34484 9278 34496
rect 9585 34493 9597 34496
rect 9631 34493 9643 34527
rect 9585 34487 9643 34493
rect 9950 34484 9956 34536
rect 10008 34524 10014 34536
rect 10152 34524 10180 34555
rect 10778 34552 10784 34604
rect 10836 34552 10842 34604
rect 10870 34552 10876 34604
rect 10928 34552 10934 34604
rect 11072 34601 11100 34632
rect 11698 34620 11704 34632
rect 11756 34620 11762 34672
rect 11057 34595 11115 34601
rect 11057 34561 11069 34595
rect 11103 34561 11115 34595
rect 11057 34555 11115 34561
rect 11149 34595 11207 34601
rect 11149 34561 11161 34595
rect 11195 34561 11207 34595
rect 11149 34555 11207 34561
rect 11333 34595 11391 34601
rect 11333 34561 11345 34595
rect 11379 34592 11391 34595
rect 11379 34564 11560 34592
rect 11379 34561 11391 34564
rect 11333 34555 11391 34561
rect 10008 34496 10180 34524
rect 10413 34527 10471 34533
rect 10008 34484 10014 34496
rect 10413 34493 10425 34527
rect 10459 34524 10471 34527
rect 10888 34524 10916 34552
rect 11164 34524 11192 34555
rect 10459 34496 11192 34524
rect 10459 34493 10471 34496
rect 10413 34487 10471 34493
rect 10612 34465 10640 34496
rect 11532 34465 11560 34564
rect 11808 34533 11836 34700
rect 12618 34688 12624 34700
rect 12676 34688 12682 34740
rect 13906 34688 13912 34740
rect 13964 34688 13970 34740
rect 14200 34700 15608 34728
rect 12434 34620 12440 34672
rect 12492 34620 12498 34672
rect 13722 34620 13728 34672
rect 13780 34660 13786 34672
rect 14200 34660 14228 34700
rect 13780 34632 14228 34660
rect 13780 34620 13786 34632
rect 14918 34620 14924 34672
rect 14976 34620 14982 34672
rect 15470 34620 15476 34672
rect 15528 34620 15534 34672
rect 15580 34660 15608 34700
rect 15654 34688 15660 34740
rect 15712 34728 15718 34740
rect 15933 34731 15991 34737
rect 15933 34728 15945 34731
rect 15712 34700 15945 34728
rect 15712 34688 15718 34700
rect 15933 34697 15945 34700
rect 15979 34697 15991 34731
rect 15933 34691 15991 34697
rect 17402 34688 17408 34740
rect 17460 34688 17466 34740
rect 17586 34688 17592 34740
rect 17644 34728 17650 34740
rect 19978 34728 19984 34740
rect 17644 34700 18552 34728
rect 17644 34688 17650 34700
rect 15580 34632 15884 34660
rect 11885 34595 11943 34601
rect 11885 34561 11897 34595
rect 11931 34592 11943 34595
rect 11931 34564 12112 34592
rect 11931 34561 11943 34564
rect 11885 34555 11943 34561
rect 11793 34527 11851 34533
rect 11793 34493 11805 34527
rect 11839 34493 11851 34527
rect 11793 34487 11851 34493
rect 10597 34459 10655 34465
rect 10597 34425 10609 34459
rect 10643 34456 10655 34459
rect 11517 34459 11575 34465
rect 10643 34428 10677 34456
rect 10643 34425 10655 34428
rect 10597 34419 10655 34425
rect 11517 34425 11529 34459
rect 11563 34425 11575 34459
rect 12084 34456 12112 34564
rect 13538 34552 13544 34604
rect 13596 34592 13602 34604
rect 14458 34592 14464 34604
rect 13596 34564 14464 34592
rect 13596 34552 13602 34564
rect 14458 34552 14464 34564
rect 14516 34552 14522 34604
rect 15856 34601 15884 34632
rect 16114 34620 16120 34672
rect 16172 34660 16178 34672
rect 18524 34660 18552 34700
rect 18708 34700 19984 34728
rect 18708 34660 18736 34700
rect 19978 34688 19984 34700
rect 20036 34688 20042 34740
rect 20158 34731 20216 34737
rect 20158 34697 20170 34731
rect 20204 34728 20216 34731
rect 21726 34728 21732 34740
rect 20204 34700 21732 34728
rect 20204 34697 20216 34700
rect 20158 34691 20216 34697
rect 21726 34688 21732 34700
rect 21784 34688 21790 34740
rect 21818 34688 21824 34740
rect 21876 34688 21882 34740
rect 21910 34688 21916 34740
rect 21968 34728 21974 34740
rect 22465 34731 22523 34737
rect 22465 34728 22477 34731
rect 21968 34700 22477 34728
rect 21968 34688 21974 34700
rect 22465 34697 22477 34700
rect 22511 34697 22523 34731
rect 22465 34691 22523 34697
rect 22922 34688 22928 34740
rect 22980 34728 22986 34740
rect 25409 34731 25467 34737
rect 25409 34728 25421 34731
rect 22980 34700 25421 34728
rect 22980 34688 22986 34700
rect 25409 34697 25421 34700
rect 25455 34697 25467 34731
rect 25409 34691 25467 34697
rect 25501 34731 25559 34737
rect 25501 34697 25513 34731
rect 25547 34728 25559 34731
rect 28261 34731 28319 34737
rect 28261 34728 28273 34731
rect 25547 34700 28273 34728
rect 25547 34697 25559 34700
rect 25501 34691 25559 34697
rect 28261 34697 28273 34700
rect 28307 34697 28319 34731
rect 28261 34691 28319 34697
rect 29730 34688 29736 34740
rect 29788 34728 29794 34740
rect 30837 34731 30895 34737
rect 30837 34728 30849 34731
rect 29788 34700 30849 34728
rect 29788 34688 29794 34700
rect 30837 34697 30849 34700
rect 30883 34697 30895 34731
rect 30837 34691 30895 34697
rect 30944 34700 31248 34728
rect 16172 34632 17172 34660
rect 18446 34632 18736 34660
rect 16172 34620 16178 34632
rect 15841 34595 15899 34601
rect 15841 34561 15853 34595
rect 15887 34561 15899 34595
rect 15841 34555 15899 34561
rect 16022 34552 16028 34604
rect 16080 34552 16086 34604
rect 16298 34552 16304 34604
rect 16356 34552 16362 34604
rect 16485 34595 16543 34601
rect 16485 34561 16497 34595
rect 16531 34592 16543 34595
rect 16531 34564 16712 34592
rect 16531 34561 16543 34564
rect 16485 34555 16543 34561
rect 12158 34484 12164 34536
rect 12216 34484 12222 34536
rect 13078 34524 13084 34536
rect 12268 34496 13084 34524
rect 12268 34456 12296 34496
rect 13078 34484 13084 34496
rect 13136 34484 13142 34536
rect 14001 34527 14059 34533
rect 14001 34493 14013 34527
rect 14047 34524 14059 34527
rect 15010 34524 15016 34536
rect 14047 34496 15016 34524
rect 14047 34493 14059 34496
rect 14001 34487 14059 34493
rect 15010 34484 15016 34496
rect 15068 34484 15074 34536
rect 15746 34484 15752 34536
rect 15804 34484 15810 34536
rect 16684 34465 16712 34564
rect 17034 34552 17040 34604
rect 17092 34552 17098 34604
rect 17144 34533 17172 34632
rect 18874 34620 18880 34672
rect 18932 34620 18938 34672
rect 20257 34663 20315 34669
rect 20257 34629 20269 34663
rect 20303 34660 20315 34663
rect 20349 34663 20407 34669
rect 20349 34660 20361 34663
rect 20303 34632 20361 34660
rect 20303 34629 20315 34632
rect 20257 34623 20315 34629
rect 20349 34629 20361 34632
rect 20395 34629 20407 34663
rect 22741 34663 22799 34669
rect 22741 34660 22753 34663
rect 20349 34623 20407 34629
rect 22296 34632 22753 34660
rect 22296 34604 22324 34632
rect 22741 34629 22753 34632
rect 22787 34629 22799 34663
rect 22741 34623 22799 34629
rect 23934 34620 23940 34672
rect 23992 34620 23998 34672
rect 24578 34620 24584 34672
rect 24636 34620 24642 34672
rect 24946 34620 24952 34672
rect 25004 34660 25010 34672
rect 25869 34663 25927 34669
rect 25869 34660 25881 34663
rect 25004 34632 25881 34660
rect 25004 34620 25010 34632
rect 25869 34629 25881 34632
rect 25915 34629 25927 34663
rect 30190 34660 30196 34672
rect 25869 34623 25927 34629
rect 28552 34632 29132 34660
rect 19981 34595 20039 34601
rect 19981 34561 19993 34595
rect 20027 34561 20039 34595
rect 19981 34555 20039 34561
rect 20073 34595 20131 34601
rect 20073 34561 20085 34595
rect 20119 34592 20131 34595
rect 20625 34595 20683 34601
rect 20625 34592 20637 34595
rect 20119 34564 20637 34592
rect 20119 34561 20131 34564
rect 20073 34555 20131 34561
rect 20625 34561 20637 34564
rect 20671 34592 20683 34595
rect 20671 34564 22232 34592
rect 20671 34561 20683 34564
rect 20625 34555 20683 34561
rect 17129 34527 17187 34533
rect 17129 34493 17141 34527
rect 17175 34524 17187 34527
rect 17862 34524 17868 34536
rect 17175 34496 17868 34524
rect 17175 34493 17187 34496
rect 17129 34487 17187 34493
rect 17862 34484 17868 34496
rect 17920 34484 17926 34536
rect 19153 34527 19211 34533
rect 19153 34493 19165 34527
rect 19199 34524 19211 34527
rect 19242 34524 19248 34536
rect 19199 34496 19248 34524
rect 19199 34493 19211 34496
rect 19153 34487 19211 34493
rect 19242 34484 19248 34496
rect 19300 34484 19306 34536
rect 19996 34524 20024 34555
rect 19996 34496 20300 34524
rect 12084 34428 12296 34456
rect 16669 34459 16727 34465
rect 11517 34419 11575 34425
rect 16669 34425 16681 34459
rect 16715 34425 16727 34459
rect 20272 34456 20300 34496
rect 20346 34484 20352 34536
rect 20404 34484 20410 34536
rect 20717 34527 20775 34533
rect 20717 34524 20729 34527
rect 20548 34496 20729 34524
rect 20548 34456 20576 34496
rect 20717 34493 20729 34496
rect 20763 34493 20775 34527
rect 21269 34527 21327 34533
rect 21269 34524 21281 34527
rect 20717 34487 20775 34493
rect 21100 34496 21281 34524
rect 20272 34428 20576 34456
rect 16669 34419 16727 34425
rect 4341 34391 4399 34397
rect 4341 34357 4353 34391
rect 4387 34388 4399 34391
rect 4706 34388 4712 34400
rect 4387 34360 4712 34388
rect 4387 34357 4399 34360
rect 4341 34351 4399 34357
rect 4706 34348 4712 34360
rect 4764 34388 4770 34400
rect 5074 34388 5080 34400
rect 4764 34360 5080 34388
rect 4764 34348 4770 34360
rect 5074 34348 5080 34360
rect 5132 34388 5138 34400
rect 5626 34388 5632 34400
rect 5132 34360 5632 34388
rect 5132 34348 5138 34360
rect 5626 34348 5632 34360
rect 5684 34348 5690 34400
rect 10226 34348 10232 34400
rect 10284 34348 10290 34400
rect 10318 34348 10324 34400
rect 10376 34348 10382 34400
rect 11333 34391 11391 34397
rect 11333 34357 11345 34391
rect 11379 34388 11391 34391
rect 11606 34388 11612 34400
rect 11379 34360 11612 34388
rect 11379 34357 11391 34360
rect 11333 34351 11391 34357
rect 11606 34348 11612 34360
rect 11664 34348 11670 34400
rect 16206 34348 16212 34400
rect 16264 34388 16270 34400
rect 16485 34391 16543 34397
rect 16485 34388 16497 34391
rect 16264 34360 16497 34388
rect 16264 34348 16270 34360
rect 16485 34357 16497 34360
rect 16531 34357 16543 34391
rect 16485 34351 16543 34357
rect 20346 34348 20352 34400
rect 20404 34388 20410 34400
rect 20533 34391 20591 34397
rect 20533 34388 20545 34391
rect 20404 34360 20545 34388
rect 20404 34348 20410 34360
rect 20533 34357 20545 34360
rect 20579 34388 20591 34391
rect 21100 34388 21128 34496
rect 21269 34493 21281 34496
rect 21315 34493 21327 34527
rect 21997 34527 22055 34533
rect 21997 34524 22009 34527
rect 21269 34487 21327 34493
rect 21928 34496 22009 34524
rect 21818 34416 21824 34468
rect 21876 34456 21882 34468
rect 21928 34456 21956 34496
rect 21997 34493 22009 34496
rect 22043 34493 22055 34527
rect 21997 34487 22055 34493
rect 22094 34484 22100 34536
rect 22152 34484 22158 34536
rect 22204 34533 22232 34564
rect 22278 34552 22284 34604
rect 22336 34552 22342 34604
rect 22649 34595 22707 34601
rect 22649 34561 22661 34595
rect 22695 34561 22707 34595
rect 22649 34555 22707 34561
rect 22189 34527 22247 34533
rect 22189 34493 22201 34527
rect 22235 34524 22247 34527
rect 22462 34524 22468 34536
rect 22235 34496 22468 34524
rect 22235 34493 22247 34496
rect 22189 34487 22247 34493
rect 22462 34484 22468 34496
rect 22520 34484 22526 34536
rect 22664 34456 22692 34555
rect 22830 34552 22836 34604
rect 22888 34552 22894 34604
rect 24854 34552 24860 34604
rect 24912 34552 24918 34604
rect 25222 34552 25228 34604
rect 25280 34552 25286 34604
rect 25593 34595 25651 34601
rect 25593 34561 25605 34595
rect 25639 34592 25651 34595
rect 26053 34595 26111 34601
rect 26053 34592 26065 34595
rect 25639 34564 26065 34592
rect 25639 34561 25651 34564
rect 25593 34555 25651 34561
rect 26053 34561 26065 34564
rect 26099 34561 26111 34595
rect 26053 34555 26111 34561
rect 26142 34552 26148 34604
rect 26200 34552 26206 34604
rect 28552 34601 28580 34632
rect 28537 34595 28595 34601
rect 28537 34561 28549 34595
rect 28583 34561 28595 34595
rect 28537 34555 28595 34561
rect 28718 34552 28724 34604
rect 28776 34552 28782 34604
rect 29104 34601 29132 34632
rect 29840 34632 30196 34660
rect 28905 34595 28963 34601
rect 28905 34561 28917 34595
rect 28951 34561 28963 34595
rect 28905 34555 28963 34561
rect 29089 34595 29147 34601
rect 29089 34561 29101 34595
rect 29135 34592 29147 34595
rect 29178 34592 29184 34604
rect 29135 34564 29184 34592
rect 29135 34561 29147 34564
rect 29089 34555 29147 34561
rect 23109 34527 23167 34533
rect 23109 34493 23121 34527
rect 23155 34524 23167 34527
rect 23842 34524 23848 34536
rect 23155 34496 23848 34524
rect 23155 34493 23167 34496
rect 23109 34487 23167 34493
rect 23842 34484 23848 34496
rect 23900 34484 23906 34536
rect 25130 34484 25136 34536
rect 25188 34484 25194 34536
rect 28442 34484 28448 34536
rect 28500 34484 28506 34536
rect 28626 34484 28632 34536
rect 28684 34484 28690 34536
rect 21876 34428 22692 34456
rect 21876 34416 21882 34428
rect 23014 34416 23020 34468
rect 23072 34416 23078 34468
rect 27890 34416 27896 34468
rect 27948 34456 27954 34468
rect 28920 34456 28948 34555
rect 29178 34552 29184 34564
rect 29236 34552 29242 34604
rect 29270 34552 29276 34604
rect 29328 34592 29334 34604
rect 29840 34601 29868 34632
rect 30190 34620 30196 34632
rect 30248 34660 30254 34672
rect 30745 34663 30803 34669
rect 30248 34632 30420 34660
rect 30248 34620 30254 34632
rect 29641 34595 29699 34601
rect 29641 34592 29653 34595
rect 29328 34564 29653 34592
rect 29328 34552 29334 34564
rect 29641 34561 29653 34564
rect 29687 34561 29699 34595
rect 29641 34555 29699 34561
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 28994 34484 29000 34536
rect 29052 34524 29058 34536
rect 29549 34527 29607 34533
rect 29549 34524 29561 34527
rect 29052 34496 29561 34524
rect 29052 34484 29058 34496
rect 29549 34493 29561 34496
rect 29595 34493 29607 34527
rect 29549 34487 29607 34493
rect 27948 34428 28948 34456
rect 27948 34416 27954 34428
rect 22094 34388 22100 34400
rect 20579 34360 22100 34388
rect 20579 34357 20591 34360
rect 20533 34351 20591 34357
rect 22094 34348 22100 34360
rect 22152 34388 22158 34400
rect 22830 34388 22836 34400
rect 22152 34360 22836 34388
rect 22152 34348 22158 34360
rect 22830 34348 22836 34360
rect 22888 34348 22894 34400
rect 28994 34348 29000 34400
rect 29052 34348 29058 34400
rect 29656 34388 29684 34555
rect 30098 34552 30104 34604
rect 30156 34552 30162 34604
rect 30282 34552 30288 34604
rect 30340 34552 30346 34604
rect 30392 34601 30420 34632
rect 30745 34629 30757 34663
rect 30791 34660 30803 34663
rect 30944 34660 30972 34700
rect 30791 34632 30972 34660
rect 31220 34660 31248 34700
rect 31662 34688 31668 34740
rect 31720 34688 31726 34740
rect 31754 34660 31760 34672
rect 31220 34632 31760 34660
rect 30791 34629 30803 34632
rect 30745 34623 30803 34629
rect 31754 34620 31760 34632
rect 31812 34620 31818 34672
rect 31849 34663 31907 34669
rect 31849 34629 31861 34663
rect 31895 34660 31907 34663
rect 32125 34663 32183 34669
rect 32125 34660 32137 34663
rect 31895 34632 32137 34660
rect 31895 34629 31907 34632
rect 31849 34623 31907 34629
rect 32125 34629 32137 34632
rect 32171 34629 32183 34663
rect 32125 34623 32183 34629
rect 30377 34595 30435 34601
rect 30377 34561 30389 34595
rect 30423 34561 30435 34595
rect 30377 34555 30435 34561
rect 30469 34595 30527 34601
rect 30469 34561 30481 34595
rect 30515 34592 30527 34595
rect 30650 34592 30656 34604
rect 30515 34564 30656 34592
rect 30515 34561 30527 34564
rect 30469 34555 30527 34561
rect 30650 34552 30656 34564
rect 30708 34552 30714 34604
rect 31018 34552 31024 34604
rect 31076 34552 31082 34604
rect 31481 34595 31539 34601
rect 31481 34561 31493 34595
rect 31527 34561 31539 34595
rect 31481 34555 31539 34561
rect 31573 34595 31631 34601
rect 31573 34561 31585 34595
rect 31619 34561 31631 34595
rect 32030 34592 32036 34604
rect 31573 34555 31631 34561
rect 31726 34564 32036 34592
rect 29733 34527 29791 34533
rect 29733 34493 29745 34527
rect 29779 34524 29791 34527
rect 29914 34524 29920 34536
rect 29779 34496 29920 34524
rect 29779 34493 29791 34496
rect 29733 34487 29791 34493
rect 29914 34484 29920 34496
rect 29972 34484 29978 34536
rect 30009 34527 30067 34533
rect 30009 34493 30021 34527
rect 30055 34524 30067 34527
rect 31113 34527 31171 34533
rect 31113 34524 31125 34527
rect 30055 34496 30420 34524
rect 30055 34493 30067 34496
rect 30009 34487 30067 34493
rect 30392 34456 30420 34496
rect 30576 34496 31125 34524
rect 30466 34456 30472 34468
rect 30392 34428 30472 34456
rect 30466 34416 30472 34428
rect 30524 34416 30530 34468
rect 30576 34388 30604 34496
rect 31113 34493 31125 34496
rect 31159 34493 31171 34527
rect 31113 34487 31171 34493
rect 30650 34416 30656 34468
rect 30708 34456 30714 34468
rect 31496 34456 31524 34555
rect 31588 34524 31616 34555
rect 31726 34524 31754 34564
rect 32030 34552 32036 34564
rect 32088 34592 32094 34604
rect 32309 34595 32367 34601
rect 32309 34592 32321 34595
rect 32088 34564 32321 34592
rect 32088 34552 32094 34564
rect 32309 34561 32321 34564
rect 32355 34561 32367 34595
rect 32309 34555 32367 34561
rect 32398 34552 32404 34604
rect 32456 34552 32462 34604
rect 34057 34595 34115 34601
rect 34057 34592 34069 34595
rect 32968 34564 34069 34592
rect 31938 34524 31944 34536
rect 31588 34496 31754 34524
rect 31864 34496 31944 34524
rect 31864 34465 31892 34496
rect 31938 34484 31944 34496
rect 31996 34484 32002 34536
rect 32122 34484 32128 34536
rect 32180 34484 32186 34536
rect 32766 34484 32772 34536
rect 32824 34524 32830 34536
rect 32968 34533 32996 34564
rect 34057 34561 34069 34564
rect 34103 34561 34115 34595
rect 34057 34555 34115 34561
rect 32953 34527 33011 34533
rect 32953 34524 32965 34527
rect 32824 34496 32965 34524
rect 32824 34484 32830 34496
rect 32953 34493 32965 34496
rect 32999 34493 33011 34527
rect 32953 34487 33011 34493
rect 33134 34484 33140 34536
rect 33192 34524 33198 34536
rect 33229 34527 33287 34533
rect 33229 34524 33241 34527
rect 33192 34496 33241 34524
rect 33192 34484 33198 34496
rect 33229 34493 33241 34496
rect 33275 34493 33287 34527
rect 33229 34487 33287 34493
rect 30708 34428 31524 34456
rect 31849 34459 31907 34465
rect 30708 34416 30714 34428
rect 31849 34425 31861 34459
rect 31895 34425 31907 34459
rect 31849 34419 31907 34425
rect 29656 34360 30604 34388
rect 31202 34348 31208 34400
rect 31260 34348 31266 34400
rect 38470 34348 38476 34400
rect 38528 34348 38534 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 5169 34187 5227 34193
rect 5169 34153 5181 34187
rect 5215 34184 5227 34187
rect 5215 34156 5580 34184
rect 5215 34153 5227 34156
rect 5169 34147 5227 34153
rect 5353 34119 5411 34125
rect 5353 34085 5365 34119
rect 5399 34085 5411 34119
rect 5552 34116 5580 34156
rect 5626 34144 5632 34196
rect 5684 34144 5690 34196
rect 6825 34187 6883 34193
rect 6825 34153 6837 34187
rect 6871 34184 6883 34187
rect 7374 34184 7380 34196
rect 6871 34156 7380 34184
rect 6871 34153 6883 34156
rect 6825 34147 6883 34153
rect 7374 34144 7380 34156
rect 7432 34144 7438 34196
rect 13078 34144 13084 34196
rect 13136 34144 13142 34196
rect 13357 34187 13415 34193
rect 13357 34153 13369 34187
rect 13403 34184 13415 34187
rect 13446 34184 13452 34196
rect 13403 34156 13452 34184
rect 13403 34153 13415 34156
rect 13357 34147 13415 34153
rect 13446 34144 13452 34156
rect 13504 34144 13510 34196
rect 13541 34187 13599 34193
rect 13541 34153 13553 34187
rect 13587 34184 13599 34187
rect 13630 34184 13636 34196
rect 13587 34156 13636 34184
rect 13587 34153 13599 34156
rect 13541 34147 13599 34153
rect 13630 34144 13636 34156
rect 13688 34144 13694 34196
rect 15286 34144 15292 34196
rect 15344 34144 15350 34196
rect 18322 34144 18328 34196
rect 18380 34184 18386 34196
rect 18509 34187 18567 34193
rect 18509 34184 18521 34187
rect 18380 34156 18521 34184
rect 18380 34144 18386 34156
rect 18509 34153 18521 34156
rect 18555 34153 18567 34187
rect 18509 34147 18567 34153
rect 29178 34144 29184 34196
rect 29236 34144 29242 34196
rect 30650 34144 30656 34196
rect 30708 34184 30714 34196
rect 30837 34187 30895 34193
rect 30837 34184 30849 34187
rect 30708 34156 30849 34184
rect 30708 34144 30714 34156
rect 30837 34153 30849 34156
rect 30883 34153 30895 34187
rect 30837 34147 30895 34153
rect 6086 34116 6092 34128
rect 5552 34088 6092 34116
rect 5353 34079 5411 34085
rect 3513 34051 3571 34057
rect 3513 34048 3525 34051
rect 3344 34020 3525 34048
rect 3145 33983 3203 33989
rect 3145 33949 3157 33983
rect 3191 33980 3203 33983
rect 3234 33980 3240 33992
rect 3191 33952 3240 33980
rect 3191 33949 3203 33952
rect 3145 33943 3203 33949
rect 3234 33940 3240 33952
rect 3292 33940 3298 33992
rect 3344 33989 3372 34020
rect 3513 34017 3525 34020
rect 3559 34017 3571 34051
rect 3513 34011 3571 34017
rect 5074 34008 5080 34060
rect 5132 34008 5138 34060
rect 5368 34048 5396 34079
rect 6086 34076 6092 34088
rect 6144 34076 6150 34128
rect 5368 34020 6776 34048
rect 3329 33983 3387 33989
rect 3329 33949 3341 33983
rect 3375 33949 3387 33983
rect 3329 33943 3387 33949
rect 3418 33940 3424 33992
rect 3476 33940 3482 33992
rect 3605 33983 3663 33989
rect 3605 33949 3617 33983
rect 3651 33980 3663 33983
rect 3973 33983 4031 33989
rect 3973 33980 3985 33983
rect 3651 33952 3985 33980
rect 3651 33949 3663 33952
rect 3605 33943 3663 33949
rect 3973 33949 3985 33952
rect 4019 33949 4031 33983
rect 3973 33943 4031 33949
rect 4522 33940 4528 33992
rect 4580 33980 4586 33992
rect 4709 33983 4767 33989
rect 4709 33980 4721 33983
rect 4580 33952 4721 33980
rect 4580 33940 4586 33952
rect 4709 33949 4721 33952
rect 4755 33949 4767 33983
rect 4709 33943 4767 33949
rect 5169 33983 5227 33989
rect 5169 33949 5181 33983
rect 5215 33980 5227 33983
rect 5350 33980 5356 33992
rect 5215 33952 5356 33980
rect 5215 33949 5227 33952
rect 5169 33943 5227 33949
rect 5350 33940 5356 33952
rect 5408 33940 5414 33992
rect 6748 33989 6776 34020
rect 10318 34008 10324 34060
rect 10376 34048 10382 34060
rect 10689 34051 10747 34057
rect 10689 34048 10701 34051
rect 10376 34020 10701 34048
rect 10376 34008 10382 34020
rect 10689 34017 10701 34020
rect 10735 34017 10747 34051
rect 10689 34011 10747 34017
rect 10965 34051 11023 34057
rect 10965 34017 10977 34051
rect 11011 34048 11023 34051
rect 11054 34048 11060 34060
rect 11011 34020 11060 34048
rect 11011 34017 11023 34020
rect 10965 34011 11023 34017
rect 11054 34008 11060 34020
rect 11112 34048 11118 34060
rect 11333 34051 11391 34057
rect 11333 34048 11345 34051
rect 11112 34020 11345 34048
rect 11112 34008 11118 34020
rect 11333 34017 11345 34020
rect 11379 34048 11391 34051
rect 12158 34048 12164 34060
rect 11379 34020 12164 34048
rect 11379 34017 11391 34020
rect 11333 34011 11391 34017
rect 12158 34008 12164 34020
rect 12216 34008 12222 34060
rect 13648 34048 13676 34144
rect 30469 34119 30527 34125
rect 30469 34116 30481 34119
rect 29840 34088 30481 34116
rect 13648 34020 15148 34048
rect 6733 33983 6791 33989
rect 6733 33949 6745 33983
rect 6779 33949 6791 33983
rect 6733 33943 6791 33949
rect 6914 33940 6920 33992
rect 6972 33940 6978 33992
rect 13538 33980 13544 33992
rect 12742 33952 13544 33980
rect 13538 33940 13544 33952
rect 13596 33940 13602 33992
rect 15010 33940 15016 33992
rect 15068 33940 15074 33992
rect 15120 33989 15148 34020
rect 15746 34008 15752 34060
rect 15804 34048 15810 34060
rect 15933 34051 15991 34057
rect 15933 34048 15945 34051
rect 15804 34020 15945 34048
rect 15804 34008 15810 34020
rect 15933 34017 15945 34020
rect 15979 34017 15991 34051
rect 15933 34011 15991 34017
rect 16206 34008 16212 34060
rect 16264 34008 16270 34060
rect 17402 34008 17408 34060
rect 17460 34048 17466 34060
rect 17773 34051 17831 34057
rect 17773 34048 17785 34051
rect 17460 34020 17785 34048
rect 17460 34008 17466 34020
rect 17773 34017 17785 34020
rect 17819 34017 17831 34051
rect 17773 34011 17831 34017
rect 19242 34008 19248 34060
rect 19300 34008 19306 34060
rect 21726 34008 21732 34060
rect 21784 34008 21790 34060
rect 21913 34051 21971 34057
rect 21913 34017 21925 34051
rect 21959 34048 21971 34051
rect 22186 34048 22192 34060
rect 21959 34020 22192 34048
rect 21959 34017 21971 34020
rect 21913 34011 21971 34017
rect 22186 34008 22192 34020
rect 22244 34048 22250 34060
rect 23198 34048 23204 34060
rect 22244 34020 23204 34048
rect 22244 34008 22250 34020
rect 23198 34008 23204 34020
rect 23256 34048 23262 34060
rect 24854 34048 24860 34060
rect 23256 34020 24860 34048
rect 23256 34008 23262 34020
rect 24854 34008 24860 34020
rect 24912 34008 24918 34060
rect 25409 34051 25467 34057
rect 25409 34017 25421 34051
rect 25455 34048 25467 34051
rect 25498 34048 25504 34060
rect 25455 34020 25504 34048
rect 25455 34017 25467 34020
rect 25409 34011 25467 34017
rect 25498 34008 25504 34020
rect 25556 34008 25562 34060
rect 27430 34008 27436 34060
rect 27488 34008 27494 34060
rect 29840 34057 29868 34088
rect 30469 34085 30481 34088
rect 30515 34085 30527 34119
rect 30469 34079 30527 34085
rect 29825 34051 29883 34057
rect 29825 34017 29837 34051
rect 29871 34017 29883 34051
rect 29825 34011 29883 34017
rect 30374 34008 30380 34060
rect 30432 34048 30438 34060
rect 30432 34020 30788 34048
rect 30432 34008 30438 34020
rect 15105 33983 15163 33989
rect 15105 33949 15117 33983
rect 15151 33949 15163 33983
rect 15105 33943 15163 33949
rect 17862 33940 17868 33992
rect 17920 33980 17926 33992
rect 18785 33983 18843 33989
rect 18785 33980 18797 33983
rect 17920 33952 18797 33980
rect 17920 33940 17926 33952
rect 18785 33949 18797 33952
rect 18831 33949 18843 33983
rect 18785 33943 18843 33949
rect 30466 33940 30472 33992
rect 30524 33940 30530 33992
rect 30760 33989 30788 34020
rect 31754 34008 31760 34060
rect 31812 34048 31818 34060
rect 32309 34051 32367 34057
rect 32309 34048 32321 34051
rect 31812 34020 32321 34048
rect 31812 34008 31818 34020
rect 32309 34017 32321 34020
rect 32355 34017 32367 34051
rect 32309 34011 32367 34017
rect 32585 34051 32643 34057
rect 32585 34017 32597 34051
rect 32631 34048 32643 34051
rect 33134 34048 33140 34060
rect 32631 34020 33140 34048
rect 32631 34017 32643 34020
rect 32585 34011 32643 34017
rect 33134 34008 33140 34020
rect 33192 34048 33198 34060
rect 33192 34020 33272 34048
rect 33192 34008 33198 34020
rect 33244 33989 33272 34020
rect 30745 33983 30803 33989
rect 30745 33949 30757 33983
rect 30791 33949 30803 33983
rect 30745 33943 30803 33949
rect 33229 33983 33287 33989
rect 33229 33949 33241 33983
rect 33275 33949 33287 33983
rect 33229 33943 33287 33949
rect 5813 33915 5871 33921
rect 5813 33881 5825 33915
rect 5859 33912 5871 33915
rect 6086 33912 6092 33924
rect 5859 33884 6092 33912
rect 5859 33881 5871 33884
rect 5813 33875 5871 33881
rect 6086 33872 6092 33884
rect 6144 33872 6150 33924
rect 8754 33872 8760 33924
rect 8812 33912 8818 33924
rect 8812 33884 9522 33912
rect 8812 33872 8818 33884
rect 11606 33872 11612 33924
rect 11664 33872 11670 33924
rect 13078 33872 13084 33924
rect 13136 33912 13142 33924
rect 13173 33915 13231 33921
rect 13173 33912 13185 33915
rect 13136 33884 13185 33912
rect 13136 33872 13142 33884
rect 13173 33881 13185 33884
rect 13219 33881 13231 33915
rect 13173 33875 13231 33881
rect 13389 33915 13447 33921
rect 13389 33881 13401 33915
rect 13435 33912 13447 33915
rect 13906 33912 13912 33924
rect 13435 33884 13912 33912
rect 13435 33881 13447 33884
rect 13389 33875 13447 33881
rect 13906 33872 13912 33884
rect 13964 33872 13970 33924
rect 17586 33912 17592 33924
rect 17434 33884 17592 33912
rect 17586 33872 17592 33884
rect 17644 33872 17650 33924
rect 18417 33915 18475 33921
rect 18417 33881 18429 33915
rect 18463 33912 18475 33915
rect 18509 33915 18567 33921
rect 18509 33912 18521 33915
rect 18463 33884 18521 33912
rect 18463 33881 18475 33884
rect 18417 33875 18475 33881
rect 18509 33881 18521 33884
rect 18555 33881 18567 33915
rect 18509 33875 18567 33881
rect 19518 33872 19524 33924
rect 19576 33872 19582 33924
rect 19978 33872 19984 33924
rect 20036 33872 20042 33924
rect 22189 33915 22247 33921
rect 22189 33881 22201 33915
rect 22235 33912 22247 33915
rect 22278 33912 22284 33924
rect 22235 33884 22284 33912
rect 22235 33881 22247 33884
rect 22189 33875 22247 33881
rect 22278 33872 22284 33884
rect 22336 33872 22342 33924
rect 22388 33884 22678 33912
rect 2498 33804 2504 33856
rect 2556 33844 2562 33856
rect 3237 33847 3295 33853
rect 3237 33844 3249 33847
rect 2556 33816 3249 33844
rect 2556 33804 2562 33816
rect 3237 33813 3249 33816
rect 3283 33813 3295 33847
rect 3237 33807 3295 33813
rect 5442 33804 5448 33856
rect 5500 33804 5506 33856
rect 5613 33847 5671 33853
rect 5613 33813 5625 33847
rect 5659 33844 5671 33847
rect 5718 33844 5724 33856
rect 5659 33816 5724 33844
rect 5659 33813 5671 33816
rect 5613 33807 5671 33813
rect 5718 33804 5724 33816
rect 5776 33804 5782 33856
rect 7006 33804 7012 33856
rect 7064 33844 7070 33856
rect 7101 33847 7159 33853
rect 7101 33844 7113 33847
rect 7064 33816 7113 33844
rect 7064 33804 7070 33816
rect 7101 33813 7113 33816
rect 7147 33844 7159 33847
rect 8018 33844 8024 33856
rect 7147 33816 8024 33844
rect 7147 33813 7159 33816
rect 7101 33807 7159 33813
rect 8018 33804 8024 33816
rect 8076 33804 8082 33856
rect 9214 33804 9220 33856
rect 9272 33804 9278 33856
rect 17034 33804 17040 33856
rect 17092 33844 17098 33856
rect 17681 33847 17739 33853
rect 17681 33844 17693 33847
rect 17092 33816 17693 33844
rect 17092 33804 17098 33816
rect 17681 33813 17693 33816
rect 17727 33844 17739 33847
rect 18693 33847 18751 33853
rect 18693 33844 18705 33847
rect 17727 33816 18705 33844
rect 17727 33813 17739 33816
rect 17681 33807 17739 33813
rect 18693 33813 18705 33816
rect 18739 33813 18751 33847
rect 18693 33807 18751 33813
rect 20346 33804 20352 33856
rect 20404 33844 20410 33856
rect 20993 33847 21051 33853
rect 20993 33844 21005 33847
rect 20404 33816 21005 33844
rect 20404 33804 20410 33816
rect 20993 33813 21005 33816
rect 21039 33813 21051 33847
rect 20993 33807 21051 33813
rect 21174 33804 21180 33856
rect 21232 33804 21238 33856
rect 21358 33804 21364 33856
rect 21416 33844 21422 33856
rect 21910 33844 21916 33856
rect 21416 33816 21916 33844
rect 21416 33804 21422 33816
rect 21910 33804 21916 33816
rect 21968 33844 21974 33856
rect 22388 33844 22416 33884
rect 27706 33872 27712 33924
rect 27764 33872 27770 33924
rect 27982 33872 27988 33924
rect 28040 33912 28046 33924
rect 28040 33884 28198 33912
rect 28040 33872 28046 33884
rect 29822 33872 29828 33924
rect 29880 33912 29886 33924
rect 29880 33884 31142 33912
rect 29880 33872 29886 33884
rect 21968 33816 22416 33844
rect 21968 33804 21974 33816
rect 23658 33804 23664 33856
rect 23716 33804 23722 33856
rect 24765 33847 24823 33853
rect 24765 33813 24777 33847
rect 24811 33844 24823 33847
rect 25038 33844 25044 33856
rect 24811 33816 25044 33844
rect 24811 33813 24823 33816
rect 24765 33807 24823 33813
rect 25038 33804 25044 33816
rect 25096 33804 25102 33856
rect 25222 33804 25228 33856
rect 25280 33844 25286 33856
rect 28074 33844 28080 33856
rect 25280 33816 28080 33844
rect 25280 33804 25286 33816
rect 28074 33804 28080 33816
rect 28132 33804 28138 33856
rect 30374 33804 30380 33856
rect 30432 33804 30438 33856
rect 30650 33804 30656 33856
rect 30708 33804 30714 33856
rect 31036 33844 31064 33884
rect 34790 33844 34796 33856
rect 31036 33816 34796 33844
rect 34790 33804 34796 33816
rect 34848 33804 34854 33856
rect 1104 33754 38824 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 38824 33754
rect 1104 33680 38824 33702
rect 3418 33600 3424 33652
rect 3476 33640 3482 33652
rect 6625 33643 6683 33649
rect 3476 33612 4384 33640
rect 3476 33600 3482 33612
rect 2498 33532 2504 33584
rect 2556 33532 2562 33584
rect 3786 33572 3792 33584
rect 3726 33544 3792 33572
rect 3786 33532 3792 33544
rect 3844 33532 3850 33584
rect 4356 33513 4384 33612
rect 6625 33609 6637 33643
rect 6671 33640 6683 33643
rect 7098 33640 7104 33652
rect 6671 33612 7104 33640
rect 6671 33609 6683 33612
rect 6625 33603 6683 33609
rect 7098 33600 7104 33612
rect 7156 33600 7162 33652
rect 10226 33600 10232 33652
rect 10284 33640 10290 33652
rect 11241 33643 11299 33649
rect 11241 33640 11253 33643
rect 10284 33612 11253 33640
rect 10284 33600 10290 33612
rect 11241 33609 11253 33612
rect 11287 33609 11299 33643
rect 21174 33640 21180 33652
rect 11241 33603 11299 33609
rect 20180 33612 21180 33640
rect 6825 33575 6883 33581
rect 6825 33541 6837 33575
rect 6871 33572 6883 33575
rect 7006 33572 7012 33584
rect 6871 33544 7012 33572
rect 6871 33541 6883 33544
rect 6825 33535 6883 33541
rect 7006 33532 7012 33544
rect 7064 33532 7070 33584
rect 9217 33575 9275 33581
rect 9217 33541 9229 33575
rect 9263 33572 9275 33575
rect 9674 33572 9680 33584
rect 9263 33544 9680 33572
rect 9263 33541 9275 33544
rect 9217 33535 9275 33541
rect 9674 33532 9680 33544
rect 9732 33532 9738 33584
rect 9766 33532 9772 33584
rect 9824 33572 9830 33584
rect 10410 33572 10416 33584
rect 9824 33544 10416 33572
rect 9824 33532 9830 33544
rect 10410 33532 10416 33544
rect 10468 33572 10474 33584
rect 10841 33575 10899 33581
rect 10841 33572 10853 33575
rect 10468 33544 10853 33572
rect 10468 33532 10474 33544
rect 10841 33541 10853 33544
rect 10887 33572 10899 33575
rect 10887 33541 10916 33572
rect 10841 33535 10916 33541
rect 4341 33507 4399 33513
rect 4341 33473 4353 33507
rect 4387 33473 4399 33507
rect 4341 33467 4399 33473
rect 4614 33464 4620 33516
rect 4672 33464 4678 33516
rect 4706 33464 4712 33516
rect 4764 33464 4770 33516
rect 4893 33507 4951 33513
rect 4893 33473 4905 33507
rect 4939 33504 4951 33507
rect 5169 33507 5227 33513
rect 5169 33504 5181 33507
rect 4939 33476 5181 33504
rect 4939 33473 4951 33476
rect 4893 33467 4951 33473
rect 5169 33473 5181 33476
rect 5215 33473 5227 33507
rect 5169 33467 5227 33473
rect 7101 33507 7159 33513
rect 7101 33473 7113 33507
rect 7147 33473 7159 33507
rect 7101 33467 7159 33473
rect 2222 33396 2228 33448
rect 2280 33396 2286 33448
rect 3973 33439 4031 33445
rect 3973 33405 3985 33439
rect 4019 33436 4031 33439
rect 4522 33436 4528 33448
rect 4019 33408 4528 33436
rect 4019 33405 4031 33408
rect 3973 33399 4031 33405
rect 4522 33396 4528 33408
rect 4580 33396 4586 33448
rect 5626 33396 5632 33448
rect 5684 33436 5690 33448
rect 5721 33439 5779 33445
rect 5721 33436 5733 33439
rect 5684 33408 5733 33436
rect 5684 33396 5690 33408
rect 5721 33405 5733 33408
rect 5767 33405 5779 33439
rect 7116 33436 7144 33467
rect 7282 33464 7288 33516
rect 7340 33464 7346 33516
rect 8110 33464 8116 33516
rect 8168 33464 8174 33516
rect 10888 33504 10916 33535
rect 11054 33532 11060 33584
rect 11112 33532 11118 33584
rect 20180 33581 20208 33612
rect 21174 33600 21180 33612
rect 21232 33600 21238 33652
rect 21637 33643 21695 33649
rect 21637 33609 21649 33643
rect 21683 33640 21695 33643
rect 22189 33643 22247 33649
rect 22189 33640 22201 33643
rect 21683 33612 22201 33640
rect 21683 33609 21695 33612
rect 21637 33603 21695 33609
rect 22189 33609 22201 33612
rect 22235 33640 22247 33643
rect 22462 33640 22468 33652
rect 22235 33612 22468 33640
rect 22235 33609 22247 33612
rect 22189 33603 22247 33609
rect 22462 33600 22468 33612
rect 22520 33600 22526 33652
rect 23658 33640 23664 33652
rect 23124 33612 23664 33640
rect 20165 33575 20223 33581
rect 20165 33541 20177 33575
rect 20211 33541 20223 33575
rect 20165 33535 20223 33541
rect 21818 33532 21824 33584
rect 21876 33572 21882 33584
rect 23124 33572 23152 33612
rect 23658 33600 23664 33612
rect 23716 33640 23722 33652
rect 23716 33612 23796 33640
rect 23716 33600 23722 33612
rect 21876 33544 23152 33572
rect 21876 33532 21882 33544
rect 10962 33504 10968 33516
rect 10888 33476 10968 33504
rect 10962 33464 10968 33476
rect 11020 33504 11026 33516
rect 11149 33507 11207 33513
rect 11149 33504 11161 33507
rect 11020 33476 11161 33504
rect 11020 33464 11026 33476
rect 11149 33473 11161 33476
rect 11195 33473 11207 33507
rect 11149 33467 11207 33473
rect 11333 33507 11391 33513
rect 11333 33473 11345 33507
rect 11379 33473 11391 33507
rect 11333 33467 11391 33473
rect 7466 33436 7472 33448
rect 7116 33408 7472 33436
rect 5721 33399 5779 33405
rect 7466 33396 7472 33408
rect 7524 33396 7530 33448
rect 7745 33439 7803 33445
rect 7745 33405 7757 33439
rect 7791 33436 7803 33439
rect 8846 33436 8852 33448
rect 7791 33408 8852 33436
rect 7791 33405 7803 33408
rect 7745 33399 7803 33405
rect 8846 33396 8852 33408
rect 8904 33396 8910 33448
rect 9214 33396 9220 33448
rect 9272 33436 9278 33448
rect 9272 33408 9444 33436
rect 9272 33396 9278 33408
rect 9416 33368 9444 33408
rect 9490 33396 9496 33448
rect 9548 33396 9554 33448
rect 10045 33439 10103 33445
rect 10045 33405 10057 33439
rect 10091 33405 10103 33439
rect 10045 33399 10103 33405
rect 10597 33439 10655 33445
rect 10597 33405 10609 33439
rect 10643 33436 10655 33439
rect 11348 33436 11376 33467
rect 15562 33464 15568 33516
rect 15620 33464 15626 33516
rect 18690 33464 18696 33516
rect 18748 33504 18754 33516
rect 18877 33507 18935 33513
rect 18877 33504 18889 33507
rect 18748 33476 18889 33504
rect 18748 33464 18754 33476
rect 18877 33473 18889 33476
rect 18923 33473 18935 33507
rect 18877 33467 18935 33473
rect 21266 33464 21272 33516
rect 21324 33464 21330 33516
rect 21928 33504 21956 33544
rect 23198 33532 23204 33584
rect 23256 33532 23262 33584
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21928 33476 22017 33504
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 22281 33507 22339 33513
rect 22281 33473 22293 33507
rect 22327 33473 22339 33507
rect 22281 33467 22339 33473
rect 22373 33507 22431 33513
rect 22373 33473 22385 33507
rect 22419 33473 22431 33507
rect 22373 33467 22431 33473
rect 10643 33408 11376 33436
rect 15749 33439 15807 33445
rect 10643 33405 10655 33408
rect 10597 33399 10655 33405
rect 15749 33405 15761 33439
rect 15795 33436 15807 33439
rect 16298 33436 16304 33448
rect 15795 33408 16304 33436
rect 15795 33405 15807 33408
rect 15749 33399 15807 33405
rect 10060 33368 10088 33399
rect 16298 33396 16304 33408
rect 16356 33396 16362 33448
rect 19334 33396 19340 33448
rect 19392 33436 19398 33448
rect 19613 33439 19671 33445
rect 19613 33436 19625 33439
rect 19392 33408 19625 33436
rect 19392 33396 19398 33408
rect 19613 33405 19625 33408
rect 19659 33436 19671 33439
rect 19889 33439 19947 33445
rect 19889 33436 19901 33439
rect 19659 33408 19901 33436
rect 19659 33405 19671 33408
rect 19613 33399 19671 33405
rect 19889 33405 19901 33408
rect 19935 33405 19947 33439
rect 19889 33399 19947 33405
rect 22296 33368 22324 33467
rect 22388 33436 22416 33467
rect 22462 33464 22468 33516
rect 22520 33504 22526 33516
rect 23014 33504 23020 33516
rect 22520 33476 23020 33504
rect 22520 33464 22526 33476
rect 23014 33464 23020 33476
rect 23072 33504 23078 33516
rect 23385 33507 23443 33513
rect 23385 33504 23397 33507
rect 23072 33476 23397 33504
rect 23072 33464 23078 33476
rect 23385 33473 23397 33476
rect 23431 33473 23443 33507
rect 23385 33467 23443 33473
rect 23474 33464 23480 33516
rect 23532 33464 23538 33516
rect 23661 33507 23719 33513
rect 23661 33473 23673 33507
rect 23707 33504 23719 33507
rect 23768 33504 23796 33612
rect 23934 33600 23940 33652
rect 23992 33640 23998 33652
rect 27525 33643 27583 33649
rect 23992 33612 24992 33640
rect 23992 33600 23998 33612
rect 24964 33572 24992 33612
rect 27525 33609 27537 33643
rect 27571 33640 27583 33643
rect 27706 33640 27712 33652
rect 27571 33612 27712 33640
rect 27571 33609 27583 33612
rect 27525 33603 27583 33609
rect 27706 33600 27712 33612
rect 27764 33600 27770 33652
rect 28353 33643 28411 33649
rect 28353 33609 28365 33643
rect 28399 33640 28411 33643
rect 28442 33640 28448 33652
rect 28399 33612 28448 33640
rect 28399 33609 28411 33612
rect 28353 33603 28411 33609
rect 28442 33600 28448 33612
rect 28500 33600 28506 33652
rect 29270 33600 29276 33652
rect 29328 33600 29334 33652
rect 30374 33600 30380 33652
rect 30432 33600 30438 33652
rect 28994 33572 29000 33584
rect 24964 33544 25622 33572
rect 28000 33544 29000 33572
rect 23707 33476 23796 33504
rect 23707 33473 23719 33476
rect 23661 33467 23719 33473
rect 24854 33464 24860 33516
rect 24912 33464 24918 33516
rect 27154 33464 27160 33516
rect 27212 33504 27218 33516
rect 27249 33507 27307 33513
rect 27249 33504 27261 33507
rect 27212 33476 27261 33504
rect 27212 33464 27218 33476
rect 27249 33473 27261 33476
rect 27295 33473 27307 33507
rect 27249 33467 27307 33473
rect 27338 33464 27344 33516
rect 27396 33504 27402 33516
rect 27433 33507 27491 33513
rect 27433 33504 27445 33507
rect 27396 33476 27445 33504
rect 27396 33464 27402 33476
rect 27433 33473 27445 33476
rect 27479 33473 27491 33507
rect 27433 33467 27491 33473
rect 27801 33507 27859 33513
rect 27801 33473 27813 33507
rect 27847 33473 27859 33507
rect 27801 33467 27859 33473
rect 23753 33439 23811 33445
rect 23753 33436 23765 33439
rect 22388 33408 23765 33436
rect 23753 33405 23765 33408
rect 23799 33405 23811 33439
rect 23753 33399 23811 33405
rect 25133 33439 25191 33445
rect 25133 33405 25145 33439
rect 25179 33436 25191 33439
rect 27816 33436 27844 33467
rect 27890 33464 27896 33516
rect 27948 33464 27954 33516
rect 28000 33513 28028 33544
rect 28994 33532 29000 33544
rect 29052 33532 29058 33584
rect 29730 33532 29736 33584
rect 29788 33532 29794 33584
rect 30392 33572 30420 33600
rect 30745 33575 30803 33581
rect 30745 33572 30757 33575
rect 30392 33544 30757 33572
rect 30745 33541 30757 33544
rect 30791 33541 30803 33575
rect 34790 33572 34796 33584
rect 34730 33544 34796 33572
rect 30745 33535 30803 33541
rect 34790 33532 34796 33544
rect 34848 33572 34854 33584
rect 35526 33572 35532 33584
rect 34848 33544 35532 33572
rect 34848 33532 34854 33544
rect 35526 33532 35532 33544
rect 35584 33532 35590 33584
rect 27985 33507 28043 33513
rect 27985 33473 27997 33507
rect 28031 33473 28043 33507
rect 27985 33467 28043 33473
rect 28074 33464 28080 33516
rect 28132 33504 28138 33516
rect 28169 33507 28227 33513
rect 28169 33504 28181 33507
rect 28132 33476 28181 33504
rect 28132 33464 28138 33476
rect 28169 33473 28181 33476
rect 28215 33473 28227 33507
rect 28169 33467 28227 33473
rect 28258 33464 28264 33516
rect 28316 33464 28322 33516
rect 28445 33507 28503 33513
rect 28445 33473 28457 33507
rect 28491 33504 28503 33507
rect 28718 33504 28724 33516
rect 28491 33476 28724 33504
rect 28491 33473 28503 33476
rect 28445 33467 28503 33473
rect 28718 33464 28724 33476
rect 28776 33464 28782 33516
rect 29178 33464 29184 33516
rect 29236 33464 29242 33516
rect 33134 33464 33140 33516
rect 33192 33504 33198 33516
rect 33229 33507 33287 33513
rect 33229 33504 33241 33507
rect 33192 33476 33241 33504
rect 33192 33464 33198 33476
rect 33229 33473 33241 33476
rect 33275 33473 33287 33507
rect 33229 33467 33287 33473
rect 28537 33439 28595 33445
rect 28537 33436 28549 33439
rect 25179 33408 26280 33436
rect 27816 33408 28549 33436
rect 25179 33405 25191 33408
rect 25133 33399 25191 33405
rect 22830 33368 22836 33380
rect 4172 33340 5764 33368
rect 9416 33340 10916 33368
rect 22296 33340 22836 33368
rect 3234 33260 3240 33312
rect 3292 33300 3298 33312
rect 4172 33309 4200 33340
rect 5736 33312 5764 33340
rect 4157 33303 4215 33309
rect 4157 33300 4169 33303
rect 3292 33272 4169 33300
rect 3292 33260 3298 33272
rect 4157 33269 4169 33272
rect 4203 33269 4215 33303
rect 4157 33263 4215 33269
rect 4890 33260 4896 33312
rect 4948 33260 4954 33312
rect 5718 33260 5724 33312
rect 5776 33260 5782 33312
rect 5994 33260 6000 33312
rect 6052 33300 6058 33312
rect 6457 33303 6515 33309
rect 6457 33300 6469 33303
rect 6052 33272 6469 33300
rect 6052 33260 6058 33272
rect 6457 33269 6469 33272
rect 6503 33269 6515 33303
rect 6457 33263 6515 33269
rect 6641 33303 6699 33309
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 6917 33303 6975 33309
rect 6917 33300 6929 33303
rect 6687 33272 6929 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 6917 33269 6929 33272
rect 6963 33269 6975 33303
rect 6917 33263 6975 33269
rect 8570 33260 8576 33312
rect 8628 33300 8634 33312
rect 10888 33309 10916 33340
rect 22830 33328 22836 33340
rect 22888 33368 22894 33380
rect 23474 33368 23480 33380
rect 22888 33340 23480 33368
rect 22888 33328 22894 33340
rect 23474 33328 23480 33340
rect 23532 33328 23538 33380
rect 10689 33303 10747 33309
rect 10689 33300 10701 33303
rect 8628 33272 10701 33300
rect 8628 33260 8634 33272
rect 10689 33269 10701 33272
rect 10735 33269 10747 33303
rect 10689 33263 10747 33269
rect 10873 33303 10931 33309
rect 10873 33269 10885 33303
rect 10919 33269 10931 33303
rect 10873 33263 10931 33269
rect 15378 33260 15384 33312
rect 15436 33260 15442 33312
rect 18690 33260 18696 33312
rect 18748 33260 18754 33312
rect 21821 33303 21879 33309
rect 21821 33269 21833 33303
rect 21867 33300 21879 33303
rect 22002 33300 22008 33312
rect 21867 33272 22008 33300
rect 21867 33269 21879 33272
rect 21821 33263 21879 33269
rect 22002 33260 22008 33272
rect 22060 33260 22066 33312
rect 23290 33260 23296 33312
rect 23348 33300 23354 33312
rect 23569 33303 23627 33309
rect 23569 33300 23581 33303
rect 23348 33272 23581 33300
rect 23348 33260 23354 33272
rect 23569 33269 23581 33272
rect 23615 33269 23627 33303
rect 23768 33300 23796 33399
rect 26252 33380 26280 33408
rect 28537 33405 28549 33408
rect 28583 33405 28595 33439
rect 28537 33399 28595 33405
rect 29270 33396 29276 33448
rect 29328 33436 29334 33448
rect 29328 33408 30972 33436
rect 29328 33396 29334 33408
rect 26234 33328 26240 33380
rect 26292 33328 26298 33380
rect 29546 33368 29552 33380
rect 26528 33340 29552 33368
rect 26528 33312 26556 33340
rect 29546 33328 29552 33340
rect 29604 33328 29610 33380
rect 30944 33368 30972 33408
rect 31018 33396 31024 33448
rect 31076 33396 31082 33448
rect 31665 33439 31723 33445
rect 31665 33405 31677 33439
rect 31711 33405 31723 33439
rect 31665 33399 31723 33405
rect 31680 33368 31708 33399
rect 30944 33340 31708 33368
rect 26510 33300 26516 33312
rect 23768 33272 26516 33300
rect 23569 33263 23627 33269
rect 26510 33260 26516 33272
rect 26568 33260 26574 33312
rect 26602 33260 26608 33312
rect 26660 33260 26666 33312
rect 27062 33260 27068 33312
rect 27120 33260 27126 33312
rect 27982 33260 27988 33312
rect 28040 33300 28046 33312
rect 28442 33300 28448 33312
rect 28040 33272 28448 33300
rect 28040 33260 28046 33272
rect 28442 33260 28448 33272
rect 28500 33260 28506 33312
rect 30742 33260 30748 33312
rect 30800 33300 30806 33312
rect 31113 33303 31171 33309
rect 31113 33300 31125 33303
rect 30800 33272 31125 33300
rect 30800 33260 30806 33272
rect 31113 33269 31125 33272
rect 31159 33269 31171 33303
rect 33244 33300 33272 33467
rect 33502 33396 33508 33448
rect 33560 33396 33566 33448
rect 33594 33396 33600 33448
rect 33652 33436 33658 33448
rect 34238 33436 34244 33448
rect 33652 33408 34244 33436
rect 33652 33396 33658 33408
rect 34238 33396 34244 33408
rect 34296 33436 34302 33448
rect 34977 33439 35035 33445
rect 34977 33436 34989 33439
rect 34296 33408 34989 33436
rect 34296 33396 34302 33408
rect 34977 33405 34989 33408
rect 35023 33436 35035 33439
rect 35621 33439 35679 33445
rect 35621 33436 35633 33439
rect 35023 33408 35633 33436
rect 35023 33405 35035 33408
rect 34977 33399 35035 33405
rect 35621 33405 35633 33408
rect 35667 33405 35679 33439
rect 35621 33399 35679 33405
rect 34514 33328 34520 33380
rect 34572 33368 34578 33380
rect 35069 33371 35127 33377
rect 35069 33368 35081 33371
rect 34572 33340 35081 33368
rect 34572 33328 34578 33340
rect 35069 33337 35081 33340
rect 35115 33337 35127 33371
rect 35069 33331 35127 33337
rect 38470 33328 38476 33380
rect 38528 33328 38534 33380
rect 34790 33300 34796 33312
rect 33244 33272 34796 33300
rect 31113 33263 31171 33269
rect 34790 33260 34796 33272
rect 34848 33260 34854 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 4890 33096 4896 33108
rect 3804 33068 4896 33096
rect 3418 32852 3424 32904
rect 3476 32852 3482 32904
rect 3605 32895 3663 32901
rect 3605 32861 3617 32895
rect 3651 32892 3663 32895
rect 3804 32892 3832 33068
rect 4890 33056 4896 33068
rect 4948 33056 4954 33108
rect 9674 33056 9680 33108
rect 9732 33056 9738 33108
rect 10597 33099 10655 33105
rect 10597 33065 10609 33099
rect 10643 33096 10655 33099
rect 10778 33096 10784 33108
rect 10643 33068 10784 33096
rect 10643 33065 10655 33068
rect 10597 33059 10655 33065
rect 10778 33056 10784 33068
rect 10836 33056 10842 33108
rect 10962 33056 10968 33108
rect 11020 33056 11026 33108
rect 11149 33099 11207 33105
rect 11149 33065 11161 33099
rect 11195 33096 11207 33099
rect 11790 33096 11796 33108
rect 11195 33068 11796 33096
rect 11195 33065 11207 33068
rect 11149 33059 11207 33065
rect 11790 33056 11796 33068
rect 11848 33056 11854 33108
rect 17034 33056 17040 33108
rect 17092 33056 17098 33108
rect 18138 33056 18144 33108
rect 18196 33056 18202 33108
rect 19518 33056 19524 33108
rect 19576 33096 19582 33108
rect 19889 33099 19947 33105
rect 19889 33096 19901 33099
rect 19576 33068 19901 33096
rect 19576 33056 19582 33068
rect 19889 33065 19901 33068
rect 19935 33065 19947 33099
rect 19889 33059 19947 33065
rect 22005 33099 22063 33105
rect 22005 33065 22017 33099
rect 22051 33065 22063 33099
rect 22005 33059 22063 33065
rect 22189 33099 22247 33105
rect 22189 33065 22201 33099
rect 22235 33096 22247 33099
rect 22278 33096 22284 33108
rect 22235 33068 22284 33096
rect 22235 33065 22247 33068
rect 22189 33059 22247 33065
rect 11054 33028 11060 33040
rect 8956 33000 11060 33028
rect 3878 32920 3884 32972
rect 3936 32960 3942 32972
rect 5721 32963 5779 32969
rect 5721 32960 5733 32963
rect 3936 32932 5733 32960
rect 3936 32920 3942 32932
rect 5721 32929 5733 32932
rect 5767 32929 5779 32963
rect 5721 32923 5779 32929
rect 5994 32920 6000 32972
rect 6052 32920 6058 32972
rect 7282 32920 7288 32972
rect 7340 32960 7346 32972
rect 7340 32932 8616 32960
rect 7340 32920 7346 32932
rect 7760 32901 7788 32932
rect 8588 32904 8616 32932
rect 8846 32920 8852 32972
rect 8904 32960 8910 32972
rect 8956 32969 8984 33000
rect 8941 32963 8999 32969
rect 8941 32960 8953 32963
rect 8904 32932 8953 32960
rect 8904 32920 8910 32932
rect 8941 32929 8953 32932
rect 8987 32929 8999 32963
rect 8941 32923 8999 32929
rect 9585 32963 9643 32969
rect 9585 32929 9597 32963
rect 9631 32960 9643 32963
rect 10137 32963 10195 32969
rect 10137 32960 10149 32963
rect 9631 32932 10149 32960
rect 9631 32929 9643 32932
rect 9585 32923 9643 32929
rect 10137 32929 10149 32932
rect 10183 32929 10195 32963
rect 10137 32923 10195 32929
rect 3651 32864 3832 32892
rect 7745 32895 7803 32901
rect 3651 32861 3663 32864
rect 3605 32855 3663 32861
rect 7745 32861 7757 32895
rect 7791 32861 7803 32895
rect 7745 32855 7803 32861
rect 7837 32895 7895 32901
rect 7837 32861 7849 32895
rect 7883 32861 7895 32895
rect 7837 32855 7895 32861
rect 3513 32827 3571 32833
rect 3513 32793 3525 32827
rect 3559 32824 3571 32827
rect 4157 32827 4215 32833
rect 4157 32824 4169 32827
rect 3559 32796 4169 32824
rect 3559 32793 3571 32796
rect 3513 32787 3571 32793
rect 4157 32793 4169 32796
rect 4203 32793 4215 32827
rect 4157 32787 4215 32793
rect 4448 32796 4646 32824
rect 3694 32716 3700 32768
rect 3752 32756 3758 32768
rect 3970 32756 3976 32768
rect 3752 32728 3976 32756
rect 3752 32716 3758 32728
rect 3970 32716 3976 32728
rect 4028 32756 4034 32768
rect 4448 32756 4476 32796
rect 7006 32784 7012 32836
rect 7064 32784 7070 32836
rect 7852 32824 7880 32855
rect 8018 32852 8024 32904
rect 8076 32892 8082 32904
rect 8389 32895 8447 32901
rect 8389 32892 8401 32895
rect 8076 32864 8401 32892
rect 8076 32852 8082 32864
rect 8389 32861 8401 32864
rect 8435 32861 8447 32895
rect 8389 32855 8447 32861
rect 7484 32796 7880 32824
rect 7484 32768 7512 32796
rect 4028 32728 4476 32756
rect 4028 32716 4034 32728
rect 5626 32716 5632 32768
rect 5684 32716 5690 32768
rect 7466 32716 7472 32768
rect 7524 32716 7530 32768
rect 7558 32716 7564 32768
rect 7616 32716 7622 32768
rect 8404 32756 8432 32855
rect 8570 32852 8576 32904
rect 8628 32852 8634 32904
rect 9861 32895 9919 32901
rect 9861 32861 9873 32895
rect 9907 32861 9919 32895
rect 9861 32855 9919 32861
rect 8481 32827 8539 32833
rect 8481 32793 8493 32827
rect 8527 32824 8539 32827
rect 9876 32824 9904 32855
rect 9950 32852 9956 32904
rect 10008 32892 10014 32904
rect 10888 32901 10916 33000
rect 11054 32988 11060 33000
rect 11112 32988 11118 33040
rect 15197 33031 15255 33037
rect 15197 32997 15209 33031
rect 15243 33028 15255 33031
rect 15562 33028 15568 33040
rect 15243 33000 15568 33028
rect 15243 32997 15255 33000
rect 15197 32991 15255 32997
rect 15562 32988 15568 33000
rect 15620 33028 15626 33040
rect 15930 33028 15936 33040
rect 15620 33000 15936 33028
rect 15620 32988 15626 33000
rect 15930 32988 15936 33000
rect 15988 33028 15994 33040
rect 16669 33031 16727 33037
rect 16669 33028 16681 33031
rect 15988 33000 16681 33028
rect 15988 32988 15994 33000
rect 16669 32997 16681 33000
rect 16715 33028 16727 33031
rect 17957 33031 18015 33037
rect 17957 33028 17969 33031
rect 16715 33000 17969 33028
rect 16715 32997 16727 33000
rect 16669 32991 16727 32997
rect 17957 32997 17969 33000
rect 18003 32997 18015 33031
rect 17957 32991 18015 32997
rect 20073 33031 20131 33037
rect 20073 32997 20085 33031
rect 20119 33028 20131 33031
rect 20438 33028 20444 33040
rect 20119 33000 20444 33028
rect 20119 32997 20131 33000
rect 20073 32991 20131 32997
rect 20438 32988 20444 33000
rect 20496 33028 20502 33040
rect 22020 33028 22048 33059
rect 22278 33056 22284 33068
rect 22336 33056 22342 33108
rect 24397 33099 24455 33105
rect 24397 33065 24409 33099
rect 24443 33096 24455 33099
rect 25498 33096 25504 33108
rect 24443 33068 25504 33096
rect 24443 33065 24455 33068
rect 24397 33059 24455 33065
rect 25498 33056 25504 33068
rect 25556 33056 25562 33108
rect 26234 33056 26240 33108
rect 26292 33056 26298 33108
rect 27890 33056 27896 33108
rect 27948 33096 27954 33108
rect 27985 33099 28043 33105
rect 27985 33096 27997 33099
rect 27948 33068 27997 33096
rect 27948 33056 27954 33068
rect 27985 33065 27997 33068
rect 28031 33096 28043 33099
rect 28626 33096 28632 33108
rect 28031 33068 28632 33096
rect 28031 33065 28043 33068
rect 27985 33059 28043 33065
rect 28626 33056 28632 33068
rect 28684 33056 28690 33108
rect 30650 33056 30656 33108
rect 30708 33056 30714 33108
rect 31662 33056 31668 33108
rect 31720 33096 31726 33108
rect 32766 33096 32772 33108
rect 31720 33068 32772 33096
rect 31720 33056 31726 33068
rect 32766 33056 32772 33068
rect 32824 33056 32830 33108
rect 33502 33056 33508 33108
rect 33560 33096 33566 33108
rect 33597 33099 33655 33105
rect 33597 33096 33609 33099
rect 33560 33068 33609 33096
rect 33560 33056 33566 33068
rect 33597 33065 33609 33068
rect 33643 33065 33655 33099
rect 35526 33096 35532 33108
rect 33597 33059 33655 33065
rect 33704 33068 35532 33096
rect 23290 33028 23296 33040
rect 20496 33000 21864 33028
rect 22020 33000 23296 33028
rect 20496 32988 20502 33000
rect 18690 32960 18696 32972
rect 12406 32932 18696 32960
rect 10045 32895 10103 32901
rect 10045 32892 10057 32895
rect 10008 32864 10057 32892
rect 10008 32852 10014 32864
rect 10045 32861 10057 32864
rect 10091 32892 10103 32895
rect 10689 32895 10747 32901
rect 10689 32892 10701 32895
rect 10091 32864 10701 32892
rect 10091 32861 10103 32864
rect 10045 32855 10103 32861
rect 10689 32861 10701 32864
rect 10735 32861 10747 32895
rect 10689 32855 10747 32861
rect 10873 32895 10931 32901
rect 10873 32861 10885 32895
rect 10919 32861 10931 32895
rect 10873 32855 10931 32861
rect 11054 32852 11060 32904
rect 11112 32892 11118 32904
rect 11425 32895 11483 32901
rect 11425 32892 11437 32895
rect 11112 32864 11437 32892
rect 11112 32852 11118 32864
rect 11425 32861 11437 32864
rect 11471 32892 11483 32895
rect 11609 32895 11667 32901
rect 11609 32892 11621 32895
rect 11471 32864 11621 32892
rect 11471 32861 11483 32864
rect 11425 32855 11483 32861
rect 11609 32861 11621 32864
rect 11655 32892 11667 32895
rect 12406 32892 12434 32932
rect 18690 32920 18696 32932
rect 18748 32920 18754 32972
rect 20346 32920 20352 32972
rect 20404 32920 20410 32972
rect 11655 32864 12434 32892
rect 11655 32861 11667 32864
rect 11609 32855 11667 32861
rect 14182 32852 14188 32904
rect 14240 32892 14246 32904
rect 15013 32895 15071 32901
rect 15013 32892 15025 32895
rect 14240 32864 15025 32892
rect 14240 32852 14246 32864
rect 15013 32861 15025 32864
rect 15059 32861 15071 32895
rect 15013 32855 15071 32861
rect 15289 32895 15347 32901
rect 15289 32861 15301 32895
rect 15335 32892 15347 32895
rect 15749 32895 15807 32901
rect 15749 32892 15761 32895
rect 15335 32864 15761 32892
rect 15335 32861 15347 32864
rect 15289 32855 15347 32861
rect 15749 32861 15761 32864
rect 15795 32861 15807 32895
rect 15749 32855 15807 32861
rect 16298 32852 16304 32904
rect 16356 32852 16362 32904
rect 17494 32852 17500 32904
rect 17552 32852 17558 32904
rect 17589 32895 17647 32901
rect 17589 32861 17601 32895
rect 17635 32861 17647 32895
rect 17589 32855 17647 32861
rect 8527 32796 9904 32824
rect 10229 32827 10287 32833
rect 8527 32793 8539 32796
rect 8481 32787 8539 32793
rect 10229 32793 10241 32827
rect 10275 32793 10287 32827
rect 10229 32787 10287 32793
rect 10413 32827 10471 32833
rect 10413 32793 10425 32827
rect 10459 32824 10471 32827
rect 10781 32827 10839 32833
rect 10781 32824 10793 32827
rect 10459 32796 10793 32824
rect 10459 32793 10471 32796
rect 10413 32787 10471 32793
rect 10781 32793 10793 32796
rect 10827 32793 10839 32827
rect 10781 32787 10839 32793
rect 10244 32756 10272 32787
rect 11330 32784 11336 32836
rect 11388 32784 11394 32836
rect 12158 32784 12164 32836
rect 12216 32824 12222 32836
rect 12437 32827 12495 32833
rect 12437 32824 12449 32827
rect 12216 32796 12449 32824
rect 12216 32784 12222 32796
rect 12437 32793 12449 32796
rect 12483 32824 12495 32827
rect 13078 32824 13084 32836
rect 12483 32796 13084 32824
rect 12483 32793 12495 32796
rect 12437 32787 12495 32793
rect 13078 32784 13084 32796
rect 13136 32824 13142 32836
rect 13538 32824 13544 32836
rect 13136 32796 13544 32824
rect 13136 32784 13142 32796
rect 13538 32784 13544 32796
rect 13596 32784 13602 32836
rect 13630 32784 13636 32836
rect 13688 32824 13694 32836
rect 14918 32824 14924 32836
rect 13688 32796 14924 32824
rect 13688 32784 13694 32796
rect 14918 32784 14924 32796
rect 14976 32784 14982 32836
rect 17037 32827 17095 32833
rect 17037 32793 17049 32827
rect 17083 32824 17095 32827
rect 17083 32796 17356 32824
rect 17083 32793 17095 32796
rect 17037 32787 17095 32793
rect 11146 32765 11152 32768
rect 8404 32728 10272 32756
rect 11133 32759 11152 32765
rect 11133 32725 11145 32759
rect 11133 32719 11152 32725
rect 11146 32716 11152 32719
rect 11204 32716 11210 32768
rect 14642 32716 14648 32768
rect 14700 32756 14706 32768
rect 14829 32759 14887 32765
rect 14829 32756 14841 32759
rect 14700 32728 14841 32756
rect 14700 32716 14706 32728
rect 14829 32725 14841 32728
rect 14875 32725 14887 32759
rect 14829 32719 14887 32725
rect 16942 32716 16948 32768
rect 17000 32756 17006 32768
rect 17328 32765 17356 32796
rect 17221 32759 17279 32765
rect 17221 32756 17233 32759
rect 17000 32728 17233 32756
rect 17000 32716 17006 32728
rect 17221 32725 17233 32728
rect 17267 32725 17279 32759
rect 17221 32719 17279 32725
rect 17313 32759 17371 32765
rect 17313 32725 17325 32759
rect 17359 32725 17371 32759
rect 17604 32756 17632 32855
rect 17678 32852 17684 32904
rect 17736 32852 17742 32904
rect 17773 32895 17831 32901
rect 17773 32861 17785 32895
rect 17819 32892 17831 32895
rect 18138 32892 18144 32904
rect 17819 32864 18144 32892
rect 17819 32861 17831 32864
rect 17773 32855 17831 32861
rect 18138 32852 18144 32864
rect 18196 32852 18202 32904
rect 19334 32852 19340 32904
rect 19392 32852 19398 32904
rect 21836 32833 21864 33000
rect 23290 32988 23296 33000
rect 23348 32988 23354 33040
rect 27430 33028 27436 33040
rect 26160 33000 27436 33028
rect 26160 32969 26188 33000
rect 27430 32988 27436 33000
rect 27488 32988 27494 33040
rect 28350 33028 28356 33040
rect 27632 33000 28356 33028
rect 26145 32963 26203 32969
rect 26145 32929 26157 32963
rect 26191 32929 26203 32963
rect 26145 32923 26203 32929
rect 26602 32920 26608 32972
rect 26660 32960 26666 32972
rect 26881 32963 26939 32969
rect 26881 32960 26893 32963
rect 26660 32932 26893 32960
rect 26660 32920 26666 32932
rect 26881 32929 26893 32932
rect 26927 32960 26939 32963
rect 26927 32932 27384 32960
rect 26927 32929 26939 32932
rect 26881 32923 26939 32929
rect 22186 32852 22192 32904
rect 22244 32892 22250 32904
rect 22373 32895 22431 32901
rect 22373 32892 22385 32895
rect 22244 32864 22385 32892
rect 22244 32852 22250 32864
rect 22373 32861 22385 32864
rect 22419 32861 22431 32895
rect 22373 32855 22431 32861
rect 27065 32895 27123 32901
rect 27065 32861 27077 32895
rect 27111 32892 27123 32895
rect 27154 32892 27160 32904
rect 27111 32864 27160 32892
rect 27111 32861 27123 32864
rect 27065 32855 27123 32861
rect 27154 32852 27160 32864
rect 27212 32852 27218 32904
rect 27246 32852 27252 32904
rect 27304 32852 27310 32904
rect 27356 32894 27384 32932
rect 27433 32895 27491 32901
rect 27433 32894 27445 32895
rect 27356 32866 27445 32894
rect 27433 32861 27445 32866
rect 27479 32892 27491 32895
rect 27632 32892 27660 33000
rect 28350 32988 28356 33000
rect 28408 33028 28414 33040
rect 28534 33028 28540 33040
rect 28408 33000 28540 33028
rect 28408 32988 28414 33000
rect 28534 32988 28540 33000
rect 28592 32988 28598 33040
rect 33704 33028 33732 33068
rect 35526 33056 35532 33068
rect 35584 33056 35590 33108
rect 34330 33028 34336 33040
rect 33152 33000 33732 33028
rect 33980 33000 34336 33028
rect 27798 32920 27804 32972
rect 27856 32960 27862 32972
rect 30837 32963 30895 32969
rect 30837 32960 30849 32963
rect 27856 32932 29040 32960
rect 27856 32920 27862 32932
rect 27479 32864 27660 32892
rect 27709 32895 27767 32901
rect 27479 32861 27491 32864
rect 27433 32855 27491 32861
rect 27709 32861 27721 32895
rect 27755 32892 27767 32895
rect 28718 32892 28724 32904
rect 27755 32864 28724 32892
rect 27755 32861 27767 32864
rect 27709 32855 27767 32861
rect 28718 32852 28724 32864
rect 28776 32852 28782 32904
rect 29012 32901 29040 32932
rect 29564 32932 30849 32960
rect 29564 32904 29592 32932
rect 30837 32929 30849 32932
rect 30883 32929 30895 32963
rect 30837 32923 30895 32929
rect 28997 32895 29055 32901
rect 28997 32861 29009 32895
rect 29043 32861 29055 32895
rect 28997 32855 29055 32861
rect 18325 32827 18383 32833
rect 18325 32824 18337 32827
rect 18064 32796 18337 32824
rect 17770 32756 17776 32768
rect 17604 32728 17776 32756
rect 17313 32719 17371 32725
rect 17770 32716 17776 32728
rect 17828 32756 17834 32768
rect 18064 32756 18092 32796
rect 18325 32793 18337 32796
rect 18371 32793 18383 32827
rect 18325 32787 18383 32793
rect 21821 32827 21879 32833
rect 21821 32793 21833 32827
rect 21867 32793 21879 32827
rect 21821 32787 21879 32793
rect 23934 32784 23940 32836
rect 23992 32824 23998 32836
rect 24210 32824 24216 32836
rect 23992 32796 24216 32824
rect 23992 32784 23998 32796
rect 24210 32784 24216 32796
rect 24268 32824 24274 32836
rect 24268 32796 24702 32824
rect 24268 32784 24274 32796
rect 25590 32784 25596 32836
rect 25648 32824 25654 32836
rect 25869 32827 25927 32833
rect 25869 32824 25881 32827
rect 25648 32796 25881 32824
rect 25648 32784 25654 32796
rect 25869 32793 25881 32796
rect 25915 32793 25927 32827
rect 25869 32787 25927 32793
rect 25958 32784 25964 32836
rect 26016 32824 26022 32836
rect 26605 32827 26663 32833
rect 26605 32824 26617 32827
rect 26016 32796 26617 32824
rect 26016 32784 26022 32796
rect 26605 32793 26617 32796
rect 26651 32824 26663 32827
rect 27617 32827 27675 32833
rect 26651 32796 27200 32824
rect 26651 32793 26663 32796
rect 26605 32787 26663 32793
rect 17828 32728 18092 32756
rect 18125 32759 18183 32765
rect 17828 32716 17834 32728
rect 18125 32725 18137 32759
rect 18171 32756 18183 32759
rect 18230 32756 18236 32768
rect 18171 32728 18236 32756
rect 18171 32725 18183 32728
rect 18125 32719 18183 32725
rect 18230 32716 18236 32728
rect 18288 32716 18294 32768
rect 22002 32716 22008 32768
rect 22060 32765 22066 32768
rect 22060 32759 22079 32765
rect 22067 32725 22079 32759
rect 22060 32719 22079 32725
rect 22060 32716 22066 32719
rect 26694 32716 26700 32768
rect 26752 32716 26758 32768
rect 27172 32765 27200 32796
rect 27617 32793 27629 32827
rect 27663 32824 27675 32827
rect 28258 32824 28264 32836
rect 27663 32796 28264 32824
rect 27663 32793 27675 32796
rect 27617 32787 27675 32793
rect 28258 32784 28264 32796
rect 28316 32784 28322 32836
rect 29012 32824 29040 32855
rect 29546 32852 29552 32904
rect 29604 32852 29610 32904
rect 30742 32852 30748 32904
rect 30800 32852 30806 32904
rect 30852 32892 30880 32923
rect 31018 32920 31024 32972
rect 31076 32960 31082 32972
rect 31757 32963 31815 32969
rect 31757 32960 31769 32963
rect 31076 32932 31769 32960
rect 31076 32920 31082 32932
rect 31757 32929 31769 32932
rect 31803 32929 31815 32963
rect 31757 32923 31815 32929
rect 31662 32892 31668 32904
rect 30852 32864 31668 32892
rect 31662 32852 31668 32864
rect 31720 32852 31726 32904
rect 33152 32878 33180 33000
rect 33318 32920 33324 32972
rect 33376 32960 33382 32972
rect 33980 32969 34008 33000
rect 34330 32988 34336 33000
rect 34388 32988 34394 33040
rect 34517 33031 34575 33037
rect 34517 32997 34529 33031
rect 34563 33028 34575 33031
rect 34563 33000 35020 33028
rect 34563 32997 34575 33000
rect 34517 32991 34575 32997
rect 33965 32963 34023 32969
rect 33965 32960 33977 32963
rect 33376 32932 33977 32960
rect 33376 32920 33382 32932
rect 33965 32929 33977 32932
rect 34011 32929 34023 32963
rect 33965 32923 34023 32929
rect 34149 32963 34207 32969
rect 34149 32929 34161 32963
rect 34195 32960 34207 32963
rect 34195 32932 34376 32960
rect 34195 32929 34207 32932
rect 34149 32923 34207 32929
rect 33870 32852 33876 32904
rect 33928 32892 33934 32904
rect 34164 32892 34192 32923
rect 33928 32864 34192 32892
rect 33928 32852 33934 32864
rect 34238 32852 34244 32904
rect 34296 32852 34302 32904
rect 34348 32901 34376 32932
rect 34790 32920 34796 32972
rect 34848 32960 34854 32972
rect 34885 32963 34943 32969
rect 34885 32960 34897 32963
rect 34848 32932 34897 32960
rect 34848 32920 34854 32932
rect 34885 32929 34897 32932
rect 34931 32929 34943 32963
rect 34992 32960 35020 33000
rect 35161 32963 35219 32969
rect 35161 32960 35173 32963
rect 34992 32932 35173 32960
rect 34885 32923 34943 32929
rect 35161 32929 35173 32932
rect 35207 32929 35219 32963
rect 35161 32923 35219 32929
rect 35526 32920 35532 32972
rect 35584 32960 35590 32972
rect 35584 32932 36216 32960
rect 35584 32920 35590 32932
rect 34333 32895 34391 32901
rect 34333 32861 34345 32895
rect 34379 32861 34391 32895
rect 34333 32855 34391 32861
rect 34517 32895 34575 32901
rect 34517 32861 34529 32895
rect 34563 32892 34575 32895
rect 34606 32892 34612 32904
rect 34563 32864 34612 32892
rect 34563 32861 34575 32864
rect 34517 32855 34575 32861
rect 34606 32852 34612 32864
rect 34664 32852 34670 32904
rect 36188 32836 36216 32932
rect 30006 32824 30012 32836
rect 29012 32796 30012 32824
rect 30006 32784 30012 32796
rect 30064 32824 30070 32836
rect 30285 32827 30343 32833
rect 30285 32824 30297 32827
rect 30064 32796 30297 32824
rect 30064 32784 30070 32796
rect 30285 32793 30297 32796
rect 30331 32824 30343 32827
rect 31018 32824 31024 32836
rect 30331 32796 31024 32824
rect 30331 32793 30343 32796
rect 30285 32787 30343 32793
rect 31018 32784 31024 32796
rect 31076 32784 31082 32836
rect 32033 32827 32091 32833
rect 32033 32793 32045 32827
rect 32079 32824 32091 32827
rect 32122 32824 32128 32836
rect 32079 32796 32128 32824
rect 32079 32793 32091 32796
rect 32033 32787 32091 32793
rect 32122 32784 32128 32796
rect 32180 32784 32186 32836
rect 33597 32827 33655 32833
rect 33597 32793 33609 32827
rect 33643 32824 33655 32827
rect 33965 32827 34023 32833
rect 33965 32824 33977 32827
rect 33643 32796 33977 32824
rect 33643 32793 33655 32796
rect 33597 32787 33655 32793
rect 33965 32793 33977 32796
rect 34011 32793 34023 32827
rect 33965 32787 34023 32793
rect 36170 32784 36176 32836
rect 36228 32784 36234 32836
rect 27157 32759 27215 32765
rect 27157 32725 27169 32759
rect 27203 32756 27215 32759
rect 27801 32759 27859 32765
rect 27801 32756 27813 32759
rect 27203 32728 27813 32756
rect 27203 32725 27215 32728
rect 27157 32719 27215 32725
rect 27801 32725 27813 32728
rect 27847 32756 27859 32759
rect 27982 32756 27988 32768
rect 27847 32728 27988 32756
rect 27847 32725 27859 32728
rect 27801 32719 27859 32725
rect 27982 32716 27988 32728
rect 28040 32716 28046 32768
rect 28166 32716 28172 32768
rect 28224 32716 28230 32768
rect 33502 32716 33508 32768
rect 33560 32716 33566 32768
rect 33781 32759 33839 32765
rect 33781 32725 33793 32759
rect 33827 32756 33839 32759
rect 34514 32756 34520 32768
rect 33827 32728 34520 32756
rect 33827 32725 33839 32728
rect 33781 32719 33839 32725
rect 34514 32716 34520 32728
rect 34572 32716 34578 32768
rect 36633 32759 36691 32765
rect 36633 32725 36645 32759
rect 36679 32756 36691 32759
rect 36722 32756 36728 32768
rect 36679 32728 36728 32756
rect 36679 32725 36691 32728
rect 36633 32719 36691 32725
rect 36722 32716 36728 32728
rect 36780 32716 36786 32768
rect 1104 32666 38824 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 38824 32666
rect 1104 32592 38824 32614
rect 3970 32512 3976 32564
rect 4028 32561 4034 32564
rect 4028 32555 4057 32561
rect 4045 32552 4057 32555
rect 4522 32552 4528 32564
rect 4045 32524 4528 32552
rect 4045 32521 4057 32524
rect 4028 32515 4057 32521
rect 4028 32512 4034 32515
rect 4522 32512 4528 32524
rect 4580 32512 4586 32564
rect 4706 32512 4712 32564
rect 4764 32552 4770 32564
rect 4893 32555 4951 32561
rect 4893 32552 4905 32555
rect 4764 32524 4905 32552
rect 4764 32512 4770 32524
rect 4893 32521 4905 32524
rect 4939 32521 4951 32555
rect 4893 32515 4951 32521
rect 6914 32512 6920 32564
rect 6972 32512 6978 32564
rect 7098 32512 7104 32564
rect 7156 32512 7162 32564
rect 11790 32512 11796 32564
rect 11848 32512 11854 32564
rect 12618 32512 12624 32564
rect 12676 32552 12682 32564
rect 12676 32524 12940 32552
rect 12676 32512 12682 32524
rect 3789 32487 3847 32493
rect 3789 32453 3801 32487
rect 3835 32484 3847 32487
rect 7466 32484 7472 32496
rect 3835 32456 4384 32484
rect 3835 32453 3847 32456
rect 3789 32447 3847 32453
rect 4356 32357 4384 32456
rect 6564 32456 7472 32484
rect 6564 32425 6592 32456
rect 7466 32444 7472 32456
rect 7524 32444 7530 32496
rect 9766 32444 9772 32496
rect 9824 32484 9830 32496
rect 12912 32484 12940 32524
rect 14182 32512 14188 32564
rect 14240 32512 14246 32564
rect 15654 32552 15660 32564
rect 14476 32524 15660 32552
rect 13630 32484 13636 32496
rect 9824 32456 10350 32484
rect 12834 32456 13636 32484
rect 9824 32444 9830 32456
rect 13630 32444 13636 32456
rect 13688 32444 13694 32496
rect 14476 32484 14504 32524
rect 15654 32512 15660 32524
rect 15712 32512 15718 32564
rect 16117 32555 16175 32561
rect 16117 32521 16129 32555
rect 16163 32552 16175 32555
rect 16298 32552 16304 32564
rect 16163 32524 16304 32552
rect 16163 32521 16175 32524
rect 16117 32515 16175 32521
rect 16298 32512 16304 32524
rect 16356 32512 16362 32564
rect 19334 32552 19340 32564
rect 16684 32524 19340 32552
rect 13924 32456 14504 32484
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32385 6607 32419
rect 6549 32379 6607 32385
rect 6638 32376 6644 32428
rect 6696 32376 6702 32428
rect 6733 32419 6791 32425
rect 6733 32385 6745 32419
rect 6779 32416 6791 32419
rect 6914 32416 6920 32428
rect 6779 32388 6920 32416
rect 6779 32385 6791 32388
rect 6733 32379 6791 32385
rect 6914 32376 6920 32388
rect 6972 32376 6978 32428
rect 7193 32419 7251 32425
rect 7193 32385 7205 32419
rect 7239 32416 7251 32419
rect 7558 32416 7564 32428
rect 7239 32388 7564 32416
rect 7239 32385 7251 32388
rect 7193 32379 7251 32385
rect 7558 32376 7564 32388
rect 7616 32376 7622 32428
rect 9490 32376 9496 32428
rect 9548 32416 9554 32428
rect 9585 32419 9643 32425
rect 9585 32416 9597 32419
rect 9548 32388 9597 32416
rect 9548 32376 9554 32388
rect 9585 32385 9597 32388
rect 9631 32385 9643 32419
rect 9585 32379 9643 32385
rect 13538 32376 13544 32428
rect 13596 32416 13602 32428
rect 13924 32416 13952 32456
rect 13596 32388 13952 32416
rect 13596 32376 13602 32388
rect 14090 32376 14096 32428
rect 14148 32376 14154 32428
rect 14384 32425 14412 32456
rect 14642 32444 14648 32496
rect 14700 32444 14706 32496
rect 14918 32444 14924 32496
rect 14976 32484 14982 32496
rect 14976 32456 15134 32484
rect 14976 32444 14982 32456
rect 16684 32425 16712 32524
rect 19334 32512 19340 32524
rect 19392 32512 19398 32564
rect 23750 32512 23756 32564
rect 23808 32552 23814 32564
rect 24147 32555 24205 32561
rect 24147 32552 24159 32555
rect 23808 32524 24159 32552
rect 23808 32512 23814 32524
rect 24147 32521 24159 32524
rect 24193 32552 24205 32555
rect 24302 32552 24308 32564
rect 24193 32524 24308 32552
rect 24193 32521 24205 32524
rect 24147 32515 24205 32521
rect 24302 32512 24308 32524
rect 24360 32552 24366 32564
rect 24670 32552 24676 32564
rect 24360 32524 24676 32552
rect 24360 32512 24366 32524
rect 24670 32512 24676 32524
rect 24728 32552 24734 32564
rect 24728 32524 25544 32552
rect 24728 32512 24734 32524
rect 16942 32444 16948 32496
rect 17000 32444 17006 32496
rect 18506 32444 18512 32496
rect 18564 32444 18570 32496
rect 18725 32487 18783 32493
rect 18725 32453 18737 32487
rect 18771 32484 18783 32487
rect 18874 32484 18880 32496
rect 18771 32456 18880 32484
rect 18771 32453 18783 32456
rect 18725 32447 18783 32453
rect 18874 32444 18880 32456
rect 18932 32444 18938 32496
rect 21910 32444 21916 32496
rect 21968 32484 21974 32496
rect 21968 32456 22862 32484
rect 21968 32444 21974 32456
rect 23658 32444 23664 32496
rect 23716 32484 23722 32496
rect 23937 32487 23995 32493
rect 23937 32484 23949 32487
rect 23716 32456 23949 32484
rect 23716 32444 23722 32456
rect 23937 32453 23949 32456
rect 23983 32453 23995 32487
rect 25130 32484 25136 32496
rect 23937 32447 23995 32453
rect 24596 32456 25136 32484
rect 14277 32419 14335 32425
rect 14277 32385 14289 32419
rect 14323 32385 14335 32419
rect 14277 32379 14335 32385
rect 14369 32419 14427 32425
rect 14369 32385 14381 32419
rect 14415 32385 14427 32419
rect 14369 32379 14427 32385
rect 16669 32419 16727 32425
rect 16669 32385 16681 32419
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 4341 32351 4399 32357
rect 4341 32317 4353 32351
rect 4387 32348 4399 32351
rect 4614 32348 4620 32360
rect 4387 32320 4620 32348
rect 4387 32317 4399 32320
rect 4341 32311 4399 32317
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 4798 32308 4804 32360
rect 4856 32348 4862 32360
rect 4985 32351 5043 32357
rect 4985 32348 4997 32351
rect 4856 32320 4997 32348
rect 4856 32308 4862 32320
rect 4985 32317 4997 32320
rect 5031 32317 5043 32351
rect 5626 32348 5632 32360
rect 4985 32311 5043 32317
rect 5184 32320 5632 32348
rect 3418 32240 3424 32292
rect 3476 32280 3482 32292
rect 4157 32283 4215 32289
rect 4157 32280 4169 32283
rect 3476 32252 4169 32280
rect 3476 32240 3482 32252
rect 4157 32249 4169 32252
rect 4203 32249 4215 32283
rect 4157 32243 4215 32249
rect 3973 32215 4031 32221
rect 3973 32181 3985 32215
rect 4019 32212 4031 32215
rect 5184 32212 5212 32320
rect 5626 32308 5632 32320
rect 5684 32308 5690 32360
rect 9861 32351 9919 32357
rect 9861 32317 9873 32351
rect 9907 32348 9919 32351
rect 10226 32348 10232 32360
rect 9907 32320 10232 32348
rect 9907 32317 9919 32320
rect 9861 32311 9919 32317
rect 10226 32308 10232 32320
rect 10284 32308 10290 32360
rect 12526 32308 12532 32360
rect 12584 32348 12590 32360
rect 13265 32351 13323 32357
rect 13265 32348 13277 32351
rect 12584 32320 13277 32348
rect 12584 32308 12590 32320
rect 13265 32317 13277 32320
rect 13311 32317 13323 32351
rect 14292 32348 14320 32379
rect 15378 32348 15384 32360
rect 14292 32320 15384 32348
rect 13265 32311 13323 32317
rect 15378 32308 15384 32320
rect 15436 32308 15442 32360
rect 16390 32308 16396 32360
rect 16448 32348 16454 32360
rect 16485 32351 16543 32357
rect 16485 32348 16497 32351
rect 16448 32320 16497 32348
rect 16448 32308 16454 32320
rect 16485 32317 16497 32320
rect 16531 32348 16543 32351
rect 18064 32348 18092 32402
rect 18230 32376 18236 32428
rect 18288 32416 18294 32428
rect 18969 32419 19027 32425
rect 18969 32416 18981 32419
rect 18288 32388 18981 32416
rect 18288 32376 18294 32388
rect 18969 32385 18981 32388
rect 19015 32385 19027 32419
rect 18969 32379 19027 32385
rect 19150 32376 19156 32428
rect 19208 32376 19214 32428
rect 22094 32376 22100 32428
rect 22152 32376 22158 32428
rect 24596 32425 24624 32456
rect 25130 32444 25136 32456
rect 25188 32444 25194 32496
rect 25516 32484 25544 32524
rect 25590 32512 25596 32564
rect 25648 32512 25654 32564
rect 25777 32555 25835 32561
rect 25777 32521 25789 32555
rect 25823 32552 25835 32555
rect 26694 32552 26700 32564
rect 25823 32524 26700 32552
rect 25823 32521 25835 32524
rect 25777 32515 25835 32521
rect 26694 32512 26700 32524
rect 26752 32512 26758 32564
rect 27890 32512 27896 32564
rect 27948 32512 27954 32564
rect 28261 32555 28319 32561
rect 28261 32521 28273 32555
rect 28307 32552 28319 32555
rect 28718 32552 28724 32564
rect 28307 32524 28724 32552
rect 28307 32521 28319 32524
rect 28261 32515 28319 32521
rect 28718 32512 28724 32524
rect 28776 32512 28782 32564
rect 32122 32512 32128 32564
rect 32180 32512 32186 32564
rect 32293 32555 32351 32561
rect 32293 32552 32305 32555
rect 32232 32524 32305 32552
rect 27908 32484 27936 32512
rect 28074 32484 28080 32496
rect 25516 32456 25728 32484
rect 24581 32419 24639 32425
rect 24581 32416 24593 32419
rect 24136 32388 24593 32416
rect 16531 32320 18092 32348
rect 16531 32317 16543 32320
rect 16485 32311 16543 32317
rect 22370 32308 22376 32360
rect 22428 32308 22434 32360
rect 23842 32308 23848 32360
rect 23900 32348 23906 32360
rect 24136 32348 24164 32388
rect 24581 32385 24593 32388
rect 24627 32385 24639 32419
rect 24581 32379 24639 32385
rect 24670 32376 24676 32428
rect 24728 32376 24734 32428
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32385 25007 32419
rect 24949 32379 25007 32385
rect 24964 32348 24992 32379
rect 25038 32376 25044 32428
rect 25096 32416 25102 32428
rect 25096 32388 25141 32416
rect 25096 32376 25102 32388
rect 25222 32376 25228 32428
rect 25280 32376 25286 32428
rect 25314 32376 25320 32428
rect 25372 32376 25378 32428
rect 25700 32425 25728 32456
rect 27540 32456 28080 32484
rect 25455 32419 25513 32425
rect 25455 32385 25467 32419
rect 25501 32416 25513 32419
rect 25685 32419 25743 32425
rect 25501 32388 25636 32416
rect 25501 32385 25513 32388
rect 25455 32379 25513 32385
rect 23900 32320 24164 32348
rect 23900 32308 23906 32320
rect 5261 32283 5319 32289
rect 5261 32249 5273 32283
rect 5307 32280 5319 32283
rect 6270 32280 6276 32292
rect 5307 32252 6276 32280
rect 5307 32249 5319 32252
rect 5261 32243 5319 32249
rect 6270 32240 6276 32252
rect 6328 32240 6334 32292
rect 19337 32283 19395 32289
rect 19337 32280 19349 32283
rect 18708 32252 19349 32280
rect 4019 32184 5212 32212
rect 4019 32181 4031 32184
rect 3973 32175 4031 32181
rect 5350 32172 5356 32224
rect 5408 32212 5414 32224
rect 5445 32215 5503 32221
rect 5445 32212 5457 32215
rect 5408 32184 5457 32212
rect 5408 32172 5414 32184
rect 5445 32181 5457 32184
rect 5491 32181 5503 32215
rect 5445 32175 5503 32181
rect 11330 32172 11336 32224
rect 11388 32172 11394 32224
rect 17494 32172 17500 32224
rect 17552 32212 17558 32224
rect 17954 32212 17960 32224
rect 17552 32184 17960 32212
rect 17552 32172 17558 32184
rect 17954 32172 17960 32184
rect 18012 32172 18018 32224
rect 18138 32172 18144 32224
rect 18196 32212 18202 32224
rect 18708 32221 18736 32252
rect 19337 32249 19349 32252
rect 19383 32249 19395 32283
rect 19337 32243 19395 32249
rect 18417 32215 18475 32221
rect 18417 32212 18429 32215
rect 18196 32184 18429 32212
rect 18196 32172 18202 32184
rect 18417 32181 18429 32184
rect 18463 32181 18475 32215
rect 18417 32175 18475 32181
rect 18693 32215 18751 32221
rect 18693 32181 18705 32215
rect 18739 32181 18751 32215
rect 18693 32175 18751 32181
rect 18877 32215 18935 32221
rect 18877 32181 18889 32215
rect 18923 32212 18935 32215
rect 20714 32212 20720 32224
rect 18923 32184 20720 32212
rect 18923 32181 18935 32184
rect 18877 32175 18935 32181
rect 20714 32172 20720 32184
rect 20772 32172 20778 32224
rect 24136 32221 24164 32320
rect 24320 32320 24992 32348
rect 25608 32348 25636 32388
rect 25685 32385 25697 32419
rect 25731 32385 25743 32419
rect 25685 32379 25743 32385
rect 25869 32419 25927 32425
rect 25869 32385 25881 32419
rect 25915 32416 25927 32419
rect 25958 32416 25964 32428
rect 25915 32388 25964 32416
rect 25915 32385 25927 32388
rect 25869 32379 25927 32385
rect 25884 32348 25912 32379
rect 25958 32376 25964 32388
rect 26016 32376 26022 32428
rect 26418 32376 26424 32428
rect 26476 32416 26482 32428
rect 27062 32416 27068 32428
rect 26476 32388 27068 32416
rect 26476 32376 26482 32388
rect 27062 32376 27068 32388
rect 27120 32416 27126 32428
rect 27540 32425 27568 32456
rect 28074 32444 28080 32456
rect 28132 32444 28138 32496
rect 29270 32444 29276 32496
rect 29328 32444 29334 32496
rect 32232 32484 32260 32524
rect 32293 32521 32305 32524
rect 32339 32552 32351 32555
rect 33505 32555 33563 32561
rect 33505 32552 33517 32555
rect 32339 32524 33517 32552
rect 32339 32521 32351 32524
rect 32293 32515 32351 32521
rect 33505 32521 33517 32524
rect 33551 32521 33563 32555
rect 33870 32552 33876 32564
rect 33505 32515 33563 32521
rect 33796 32524 33876 32552
rect 33796 32493 33824 32524
rect 33870 32512 33876 32524
rect 33928 32512 33934 32564
rect 34606 32512 34612 32564
rect 34664 32512 34670 32564
rect 31496 32456 32260 32484
rect 32493 32487 32551 32493
rect 27157 32419 27215 32425
rect 27157 32416 27169 32419
rect 27120 32388 27169 32416
rect 27120 32376 27126 32388
rect 27157 32385 27169 32388
rect 27203 32385 27215 32419
rect 27157 32379 27215 32385
rect 27525 32419 27583 32425
rect 27525 32385 27537 32419
rect 27571 32385 27583 32419
rect 27525 32379 27583 32385
rect 27709 32419 27767 32425
rect 27709 32385 27721 32419
rect 27755 32385 27767 32419
rect 27709 32379 27767 32385
rect 25608 32320 25912 32348
rect 27724 32348 27752 32379
rect 27798 32376 27804 32428
rect 27856 32376 27862 32428
rect 27893 32419 27951 32425
rect 27893 32385 27905 32419
rect 27939 32416 27951 32419
rect 28166 32416 28172 32428
rect 27939 32388 28172 32416
rect 27939 32385 27951 32388
rect 27893 32379 27951 32385
rect 28166 32376 28172 32388
rect 28224 32376 28230 32428
rect 30006 32376 30012 32428
rect 30064 32416 30070 32428
rect 30282 32416 30288 32428
rect 30064 32388 30288 32416
rect 30064 32376 30070 32388
rect 30282 32376 30288 32388
rect 30340 32376 30346 32428
rect 31386 32376 31392 32428
rect 31444 32376 31450 32428
rect 31496 32425 31524 32456
rect 32493 32453 32505 32487
rect 32539 32453 32551 32487
rect 33781 32487 33839 32493
rect 32493 32447 32551 32453
rect 33060 32456 33732 32484
rect 31481 32419 31539 32425
rect 31481 32385 31493 32419
rect 31527 32385 31539 32419
rect 31481 32379 31539 32385
rect 31754 32376 31760 32428
rect 31812 32376 31818 32428
rect 28074 32348 28080 32360
rect 27724 32320 28080 32348
rect 24320 32289 24348 32320
rect 28074 32308 28080 32320
rect 28132 32308 28138 32360
rect 29733 32351 29791 32357
rect 29733 32348 29745 32351
rect 28184 32320 29745 32348
rect 24305 32283 24363 32289
rect 24305 32249 24317 32283
rect 24351 32249 24363 32283
rect 24305 32243 24363 32249
rect 26694 32240 26700 32292
rect 26752 32280 26758 32292
rect 28184 32289 28212 32320
rect 29733 32317 29745 32320
rect 29779 32317 29791 32351
rect 29733 32311 29791 32317
rect 30558 32308 30564 32360
rect 30616 32348 30622 32360
rect 31021 32351 31079 32357
rect 31021 32348 31033 32351
rect 30616 32320 31033 32348
rect 30616 32308 30622 32320
rect 31021 32317 31033 32320
rect 31067 32348 31079 32351
rect 31573 32351 31631 32357
rect 31573 32348 31585 32351
rect 31067 32320 31585 32348
rect 31067 32317 31079 32320
rect 31021 32311 31079 32317
rect 31573 32317 31585 32320
rect 31619 32317 31631 32351
rect 31573 32311 31631 32317
rect 28169 32283 28227 32289
rect 26752 32252 27476 32280
rect 26752 32240 26758 32252
rect 24121 32215 24179 32221
rect 24121 32181 24133 32215
rect 24167 32181 24179 32215
rect 24121 32175 24179 32181
rect 24486 32172 24492 32224
rect 24544 32212 24550 32224
rect 24673 32215 24731 32221
rect 24673 32212 24685 32215
rect 24544 32184 24685 32212
rect 24544 32172 24550 32184
rect 24673 32181 24685 32184
rect 24719 32181 24731 32215
rect 24673 32175 24731 32181
rect 27338 32172 27344 32224
rect 27396 32172 27402 32224
rect 27448 32212 27476 32252
rect 28169 32249 28181 32283
rect 28215 32249 28227 32283
rect 32508 32280 32536 32447
rect 33060 32425 33088 32456
rect 33045 32419 33103 32425
rect 33045 32385 33057 32419
rect 33091 32385 33103 32419
rect 33045 32379 33103 32385
rect 33321 32419 33379 32425
rect 33321 32385 33333 32419
rect 33367 32416 33379 32419
rect 33502 32416 33508 32428
rect 33367 32388 33508 32416
rect 33367 32385 33379 32388
rect 33321 32379 33379 32385
rect 33502 32376 33508 32388
rect 33560 32376 33566 32428
rect 33594 32376 33600 32428
rect 33652 32376 33658 32428
rect 33704 32416 33732 32456
rect 33781 32453 33793 32487
rect 33827 32453 33839 32487
rect 33781 32447 33839 32453
rect 33870 32416 33876 32428
rect 33704 32388 33876 32416
rect 33870 32376 33876 32388
rect 33928 32416 33934 32428
rect 34057 32419 34115 32425
rect 34057 32416 34069 32419
rect 33928 32388 34069 32416
rect 33928 32376 33934 32388
rect 34057 32385 34069 32388
rect 34103 32385 34115 32419
rect 34057 32379 34115 32385
rect 34241 32419 34299 32425
rect 34241 32385 34253 32419
rect 34287 32416 34299 32419
rect 34333 32419 34391 32425
rect 34333 32416 34345 32419
rect 34287 32388 34345 32416
rect 34287 32385 34299 32388
rect 34241 32379 34299 32385
rect 34333 32385 34345 32388
rect 34379 32416 34391 32419
rect 36722 32416 36728 32428
rect 34379 32388 36728 32416
rect 34379 32385 34391 32388
rect 34333 32379 34391 32385
rect 33134 32308 33140 32360
rect 33192 32308 33198 32360
rect 33229 32351 33287 32357
rect 33229 32317 33241 32351
rect 33275 32348 33287 32351
rect 33275 32320 33456 32348
rect 33275 32317 33287 32320
rect 33229 32311 33287 32317
rect 33318 32280 33324 32292
rect 32508 32252 33324 32280
rect 28169 32243 28227 32249
rect 33318 32240 33324 32252
rect 33376 32240 33382 32292
rect 33428 32224 33456 32320
rect 34072 32280 34100 32379
rect 34425 32283 34483 32289
rect 34425 32280 34437 32283
rect 34072 32252 34437 32280
rect 34425 32249 34437 32252
rect 34471 32249 34483 32283
rect 34425 32243 34483 32249
rect 28258 32212 28264 32224
rect 27448 32184 28264 32212
rect 28258 32172 28264 32184
rect 28316 32172 28322 32224
rect 30650 32172 30656 32224
rect 30708 32212 30714 32224
rect 31205 32215 31263 32221
rect 31205 32212 31217 32215
rect 30708 32184 31217 32212
rect 30708 32172 30714 32184
rect 31205 32181 31217 32184
rect 31251 32181 31263 32215
rect 31205 32175 31263 32181
rect 32309 32215 32367 32221
rect 32309 32181 32321 32215
rect 32355 32212 32367 32215
rect 32861 32215 32919 32221
rect 32861 32212 32873 32215
rect 32355 32184 32873 32212
rect 32355 32181 32367 32184
rect 32309 32175 32367 32181
rect 32861 32181 32873 32184
rect 32907 32181 32919 32215
rect 32861 32175 32919 32181
rect 33410 32172 33416 32224
rect 33468 32212 33474 32224
rect 34532 32212 34560 32388
rect 36722 32376 36728 32388
rect 36780 32376 36786 32428
rect 34606 32308 34612 32360
rect 34664 32308 34670 32360
rect 33468 32184 34560 32212
rect 33468 32172 33474 32184
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 2222 32008 2228 32020
rect 1872 31980 2228 32008
rect 1872 31881 1900 31980
rect 2222 31968 2228 31980
rect 2280 31968 2286 32020
rect 2498 31968 2504 32020
rect 2556 32008 2562 32020
rect 4709 32011 4767 32017
rect 4709 32008 4721 32011
rect 2556 31980 4721 32008
rect 2556 31968 2562 31980
rect 4709 31977 4721 31980
rect 4755 31977 4767 32011
rect 4709 31971 4767 31977
rect 6181 32011 6239 32017
rect 6181 31977 6193 32011
rect 6227 32008 6239 32011
rect 6638 32008 6644 32020
rect 6227 31980 6644 32008
rect 6227 31977 6239 31980
rect 6181 31971 6239 31977
rect 6638 31968 6644 31980
rect 6696 31968 6702 32020
rect 10226 31968 10232 32020
rect 10284 31968 10290 32020
rect 10502 31968 10508 32020
rect 10560 32008 10566 32020
rect 10870 32008 10876 32020
rect 10560 31980 10876 32008
rect 10560 31968 10566 31980
rect 10870 31968 10876 31980
rect 10928 32008 10934 32020
rect 10928 31980 12434 32008
rect 10928 31968 10934 31980
rect 3605 31943 3663 31949
rect 3605 31909 3617 31943
rect 3651 31940 3663 31943
rect 4614 31940 4620 31952
rect 3651 31912 4620 31940
rect 3651 31909 3663 31912
rect 3605 31903 3663 31909
rect 1857 31875 1915 31881
rect 1857 31841 1869 31875
rect 1903 31841 1915 31875
rect 1857 31835 1915 31841
rect 2133 31875 2191 31881
rect 2133 31841 2145 31875
rect 2179 31872 2191 31875
rect 2498 31872 2504 31884
rect 2179 31844 2504 31872
rect 2179 31841 2191 31844
rect 2133 31835 2191 31841
rect 2498 31832 2504 31844
rect 2556 31832 2562 31884
rect 3988 31881 4016 31912
rect 4614 31900 4620 31912
rect 4672 31940 4678 31952
rect 4672 31912 5580 31940
rect 4672 31900 4678 31912
rect 5552 31881 5580 31912
rect 6270 31900 6276 31952
rect 6328 31900 6334 31952
rect 10321 31943 10379 31949
rect 10321 31909 10333 31943
rect 10367 31940 10379 31943
rect 10597 31943 10655 31949
rect 10597 31940 10609 31943
rect 10367 31912 10609 31940
rect 10367 31909 10379 31912
rect 10321 31903 10379 31909
rect 10597 31909 10609 31912
rect 10643 31909 10655 31943
rect 11146 31940 11152 31952
rect 10597 31903 10655 31909
rect 10888 31912 11152 31940
rect 3973 31875 4031 31881
rect 3973 31841 3985 31875
rect 4019 31841 4031 31875
rect 4985 31875 5043 31881
rect 4985 31872 4997 31875
rect 3973 31835 4031 31841
rect 4172 31844 4997 31872
rect 3786 31804 3792 31816
rect 3266 31776 3792 31804
rect 3786 31764 3792 31776
rect 3844 31764 3850 31816
rect 4172 31804 4200 31844
rect 4985 31841 4997 31844
rect 5031 31841 5043 31875
rect 4985 31835 5043 31841
rect 5537 31875 5595 31881
rect 5537 31841 5549 31875
rect 5583 31841 5595 31875
rect 5537 31835 5595 31841
rect 6022 31875 6080 31881
rect 6022 31841 6034 31875
rect 6068 31872 6080 31875
rect 6546 31872 6552 31884
rect 6068 31844 6552 31872
rect 6068 31841 6080 31844
rect 6022 31835 6080 31841
rect 6546 31832 6552 31844
rect 6604 31832 6610 31884
rect 6641 31875 6699 31881
rect 6641 31841 6653 31875
rect 6687 31872 6699 31875
rect 6914 31872 6920 31884
rect 6687 31844 6920 31872
rect 6687 31841 6699 31844
rect 6641 31835 6699 31841
rect 6914 31832 6920 31844
rect 6972 31872 6978 31884
rect 7282 31872 7288 31884
rect 6972 31844 7288 31872
rect 6972 31832 6978 31844
rect 7282 31832 7288 31844
rect 7340 31832 7346 31884
rect 10137 31875 10195 31881
rect 10137 31841 10149 31875
rect 10183 31872 10195 31875
rect 10502 31872 10508 31884
rect 10183 31844 10508 31872
rect 10183 31841 10195 31844
rect 10137 31835 10195 31841
rect 10502 31832 10508 31844
rect 10560 31832 10566 31884
rect 4080 31776 4200 31804
rect 4617 31807 4675 31813
rect 4080 31748 4108 31776
rect 4617 31773 4629 31807
rect 4663 31804 4675 31807
rect 5077 31807 5135 31813
rect 5077 31804 5089 31807
rect 4663 31776 5089 31804
rect 4663 31773 4675 31776
rect 4617 31767 4675 31773
rect 5077 31773 5089 31776
rect 5123 31773 5135 31807
rect 6457 31807 6515 31813
rect 6457 31804 6469 31807
rect 6435 31776 6469 31804
rect 5077 31767 5135 31773
rect 6457 31773 6469 31776
rect 6503 31773 6515 31807
rect 6457 31767 6515 31773
rect 4062 31696 4068 31748
rect 4120 31696 4126 31748
rect 6472 31736 6500 31767
rect 6730 31764 6736 31816
rect 6788 31764 6794 31816
rect 7101 31807 7159 31813
rect 7101 31804 7113 31807
rect 7079 31776 7113 31804
rect 7101 31773 7113 31776
rect 7147 31804 7159 31807
rect 7558 31804 7564 31816
rect 7147 31776 7564 31804
rect 7147 31773 7159 31776
rect 7101 31767 7159 31773
rect 7116 31736 7144 31767
rect 7558 31764 7564 31776
rect 7616 31764 7622 31816
rect 7742 31764 7748 31816
rect 7800 31804 7806 31816
rect 8113 31807 8171 31813
rect 8113 31804 8125 31807
rect 7800 31776 8125 31804
rect 7800 31764 7806 31776
rect 8113 31773 8125 31776
rect 8159 31773 8171 31807
rect 8113 31767 8171 31773
rect 10410 31764 10416 31816
rect 10468 31764 10474 31816
rect 10888 31813 10916 31912
rect 11146 31900 11152 31912
rect 11204 31900 11210 31952
rect 12406 31940 12434 31980
rect 12526 31968 12532 32020
rect 12584 31968 12590 32020
rect 14829 32011 14887 32017
rect 14829 31977 14841 32011
rect 14875 32008 14887 32011
rect 15378 32008 15384 32020
rect 14875 31980 15384 32008
rect 14875 31977 14887 31980
rect 14829 31971 14887 31977
rect 15378 31968 15384 31980
rect 15436 31968 15442 32020
rect 15933 32011 15991 32017
rect 15933 32008 15945 32011
rect 15580 31980 15945 32008
rect 12406 31912 12664 31940
rect 11330 31832 11336 31884
rect 11388 31872 11394 31884
rect 11517 31875 11575 31881
rect 11517 31872 11529 31875
rect 11388 31844 11529 31872
rect 11388 31832 11394 31844
rect 11517 31841 11529 31844
rect 11563 31841 11575 31875
rect 11517 31835 11575 31841
rect 10873 31807 10931 31813
rect 10873 31773 10885 31807
rect 10919 31773 10931 31807
rect 10873 31767 10931 31773
rect 12253 31807 12311 31813
rect 12253 31773 12265 31807
rect 12299 31773 12311 31807
rect 12253 31767 12311 31773
rect 7190 31736 7196 31748
rect 6472 31708 7196 31736
rect 7190 31696 7196 31708
rect 7248 31696 7254 31748
rect 7282 31696 7288 31748
rect 7340 31696 7346 31748
rect 7469 31739 7527 31745
rect 7469 31705 7481 31739
rect 7515 31736 7527 31739
rect 7650 31736 7656 31748
rect 7515 31708 7656 31736
rect 7515 31705 7527 31708
rect 7469 31699 7527 31705
rect 7650 31696 7656 31708
rect 7708 31696 7714 31748
rect 10597 31739 10655 31745
rect 10597 31705 10609 31739
rect 10643 31736 10655 31739
rect 10686 31736 10692 31748
rect 10643 31708 10692 31736
rect 10643 31705 10655 31708
rect 10597 31699 10655 31705
rect 10686 31696 10692 31708
rect 10744 31696 10750 31748
rect 10962 31696 10968 31748
rect 11020 31696 11026 31748
rect 11790 31736 11796 31748
rect 11532 31708 11796 31736
rect 5810 31628 5816 31680
rect 5868 31628 5874 31680
rect 5905 31671 5963 31677
rect 5905 31637 5917 31671
rect 5951 31668 5963 31671
rect 6730 31668 6736 31680
rect 5951 31640 6736 31668
rect 5951 31637 5963 31640
rect 5905 31631 5963 31637
rect 6730 31628 6736 31640
rect 6788 31628 6794 31680
rect 7558 31628 7564 31680
rect 7616 31628 7622 31680
rect 10781 31671 10839 31677
rect 10781 31637 10793 31671
rect 10827 31668 10839 31671
rect 11532 31668 11560 31708
rect 11790 31696 11796 31708
rect 11848 31736 11854 31748
rect 12268 31736 12296 31767
rect 12434 31764 12440 31816
rect 12492 31764 12498 31816
rect 12636 31813 12664 31912
rect 15286 31872 15292 31884
rect 14660 31844 15292 31872
rect 14660 31813 14688 31844
rect 15286 31832 15292 31844
rect 15344 31832 15350 31884
rect 12621 31807 12679 31813
rect 12621 31773 12633 31807
rect 12667 31773 12679 31807
rect 12621 31767 12679 31773
rect 14645 31807 14703 31813
rect 14645 31773 14657 31807
rect 14691 31773 14703 31807
rect 14645 31767 14703 31773
rect 14921 31807 14979 31813
rect 14921 31773 14933 31807
rect 14967 31804 14979 31807
rect 15013 31807 15071 31813
rect 15013 31804 15025 31807
rect 14967 31776 15025 31804
rect 14967 31773 14979 31776
rect 14921 31767 14979 31773
rect 15013 31773 15025 31776
rect 15059 31773 15071 31807
rect 15013 31767 15071 31773
rect 15194 31764 15200 31816
rect 15252 31804 15258 31816
rect 15580 31813 15608 31980
rect 15933 31977 15945 31980
rect 15979 31977 15991 32011
rect 15933 31971 15991 31977
rect 17034 31968 17040 32020
rect 17092 32008 17098 32020
rect 18506 32008 18512 32020
rect 17092 31980 18512 32008
rect 17092 31968 17098 31980
rect 18506 31968 18512 31980
rect 18564 32008 18570 32020
rect 18601 32011 18659 32017
rect 18601 32008 18613 32011
rect 18564 31980 18613 32008
rect 18564 31968 18570 31980
rect 18601 31977 18613 31980
rect 18647 31977 18659 32011
rect 18601 31971 18659 31977
rect 18874 31968 18880 32020
rect 18932 32008 18938 32020
rect 18969 32011 19027 32017
rect 18969 32008 18981 32011
rect 18932 31980 18981 32008
rect 18932 31968 18938 31980
rect 18969 31977 18981 31980
rect 19015 31977 19027 32011
rect 18969 31971 19027 31977
rect 25314 31968 25320 32020
rect 25372 32008 25378 32020
rect 25590 32008 25596 32020
rect 25372 31980 25596 32008
rect 25372 31968 25378 31980
rect 25590 31968 25596 31980
rect 25648 32008 25654 32020
rect 25961 32011 26019 32017
rect 25961 32008 25973 32011
rect 25648 31980 25973 32008
rect 25648 31968 25654 31980
rect 25961 31977 25973 31980
rect 26007 31977 26019 32011
rect 27065 32011 27123 32017
rect 25961 31971 26019 31977
rect 26436 31980 26832 32008
rect 17129 31943 17187 31949
rect 17129 31909 17141 31943
rect 17175 31940 17187 31943
rect 17678 31940 17684 31952
rect 17175 31912 17684 31940
rect 17175 31909 17187 31912
rect 17129 31903 17187 31909
rect 17678 31900 17684 31912
rect 17736 31900 17742 31952
rect 17770 31900 17776 31952
rect 17828 31940 17834 31952
rect 17828 31912 18184 31940
rect 17828 31900 17834 31912
rect 17494 31832 17500 31884
rect 17552 31872 17558 31884
rect 17865 31875 17923 31881
rect 17865 31872 17877 31875
rect 17552 31844 17877 31872
rect 17552 31832 17558 31844
rect 17865 31841 17877 31844
rect 17911 31841 17923 31875
rect 18156 31872 18184 31912
rect 18230 31900 18236 31952
rect 18288 31900 18294 31952
rect 18785 31943 18843 31949
rect 18785 31909 18797 31943
rect 18831 31940 18843 31943
rect 22557 31943 22615 31949
rect 18831 31912 19748 31940
rect 18831 31909 18843 31912
rect 18785 31903 18843 31909
rect 19150 31872 19156 31884
rect 18156 31844 19156 31872
rect 17865 31835 17923 31841
rect 15565 31807 15623 31813
rect 15565 31804 15577 31807
rect 15252 31776 15577 31804
rect 15252 31764 15258 31776
rect 15565 31773 15577 31776
rect 15611 31773 15623 31807
rect 17589 31807 17647 31813
rect 15565 31767 15623 31773
rect 16546 31776 17172 31804
rect 11848 31708 12296 31736
rect 15749 31739 15807 31745
rect 11848 31696 11854 31708
rect 15749 31705 15761 31739
rect 15795 31705 15807 31739
rect 15749 31699 15807 31705
rect 10827 31640 11560 31668
rect 10827 31637 10839 31640
rect 10781 31631 10839 31637
rect 11698 31628 11704 31680
rect 11756 31628 11762 31680
rect 14366 31628 14372 31680
rect 14424 31668 14430 31680
rect 14461 31671 14519 31677
rect 14461 31668 14473 31671
rect 14424 31640 14473 31668
rect 14424 31628 14430 31640
rect 14461 31637 14473 31640
rect 14507 31637 14519 31671
rect 15764 31668 15792 31699
rect 15930 31696 15936 31748
rect 15988 31745 15994 31748
rect 15988 31739 16007 31745
rect 15995 31705 16007 31739
rect 16298 31736 16304 31748
rect 15988 31699 16007 31705
rect 16040 31708 16304 31736
rect 15988 31696 15994 31699
rect 16040 31668 16068 31708
rect 16298 31696 16304 31708
rect 16356 31736 16362 31748
rect 16546 31736 16574 31776
rect 17144 31745 17172 31776
rect 17589 31773 17601 31807
rect 17635 31804 17647 31807
rect 18138 31804 18144 31816
rect 17635 31776 18144 31804
rect 17635 31773 17647 31776
rect 17589 31767 17647 31773
rect 18138 31764 18144 31776
rect 18196 31764 18202 31816
rect 18230 31764 18236 31816
rect 18288 31804 18294 31816
rect 19076 31813 19104 31844
rect 19150 31832 19156 31844
rect 19208 31872 19214 31884
rect 19245 31875 19303 31881
rect 19245 31872 19257 31875
rect 19208 31844 19257 31872
rect 19208 31832 19214 31844
rect 19245 31841 19257 31844
rect 19291 31841 19303 31875
rect 19720 31872 19748 31912
rect 22557 31909 22569 31943
rect 22603 31909 22615 31943
rect 22557 31903 22615 31909
rect 20070 31872 20076 31884
rect 19720 31844 20076 31872
rect 19245 31835 19303 31841
rect 20070 31832 20076 31844
rect 20128 31832 20134 31884
rect 20714 31832 20720 31884
rect 20772 31832 20778 31884
rect 22572 31872 22600 31903
rect 24762 31900 24768 31952
rect 24820 31940 24826 31952
rect 26436 31940 26464 31980
rect 24820 31912 26464 31940
rect 24820 31900 24826 31912
rect 23293 31875 23351 31881
rect 23293 31872 23305 31875
rect 22572 31844 23305 31872
rect 23293 31841 23305 31844
rect 23339 31872 23351 31875
rect 23658 31872 23664 31884
rect 23339 31844 23664 31872
rect 23339 31841 23351 31844
rect 23293 31835 23351 31841
rect 23658 31832 23664 31844
rect 23716 31832 23722 31884
rect 26602 31832 26608 31884
rect 26660 31832 26666 31884
rect 18877 31807 18935 31813
rect 18877 31804 18889 31807
rect 18288 31776 18889 31804
rect 18288 31764 18294 31776
rect 18877 31773 18889 31776
rect 18923 31773 18935 31807
rect 18877 31767 18935 31773
rect 19061 31807 19119 31813
rect 19061 31773 19073 31807
rect 19107 31773 19119 31807
rect 19061 31767 19119 31773
rect 20990 31764 20996 31816
rect 21048 31804 21054 31816
rect 21177 31807 21235 31813
rect 21177 31804 21189 31807
rect 21048 31776 21189 31804
rect 21048 31764 21054 31776
rect 21177 31773 21189 31776
rect 21223 31804 21235 31807
rect 21223 31776 22140 31804
rect 21223 31773 21235 31776
rect 21177 31767 21235 31773
rect 22112 31748 22140 31776
rect 23566 31764 23572 31816
rect 23624 31804 23630 31816
rect 23937 31807 23995 31813
rect 23937 31804 23949 31807
rect 23624 31776 23949 31804
rect 23624 31764 23630 31776
rect 23937 31773 23949 31776
rect 23983 31773 23995 31807
rect 23937 31767 23995 31773
rect 24946 31764 24952 31816
rect 25004 31764 25010 31816
rect 25038 31764 25044 31816
rect 25096 31804 25102 31816
rect 25317 31807 25375 31813
rect 25317 31804 25329 31807
rect 25096 31776 25329 31804
rect 25096 31764 25102 31776
rect 25317 31773 25329 31776
rect 25363 31773 25375 31807
rect 25317 31767 25375 31773
rect 26513 31807 26571 31813
rect 26513 31773 26525 31807
rect 26559 31804 26571 31807
rect 26620 31804 26648 31832
rect 26559 31776 26648 31804
rect 26559 31773 26571 31776
rect 26513 31767 26571 31773
rect 26694 31764 26700 31816
rect 26752 31764 26758 31816
rect 26804 31813 26832 31980
rect 27065 31977 27077 32011
rect 27111 32008 27123 32011
rect 27798 32008 27804 32020
rect 27111 31980 27804 32008
rect 27111 31977 27123 31980
rect 27065 31971 27123 31977
rect 27798 31968 27804 31980
rect 27856 31968 27862 32020
rect 28074 31968 28080 32020
rect 28132 32008 28138 32020
rect 28537 32011 28595 32017
rect 28537 32008 28549 32011
rect 28132 31980 28549 32008
rect 28132 31968 28138 31980
rect 28537 31977 28549 31980
rect 28583 31977 28595 32011
rect 28537 31971 28595 31977
rect 31386 31968 31392 32020
rect 31444 32008 31450 32020
rect 33137 32011 33195 32017
rect 33137 32008 33149 32011
rect 31444 31980 33149 32008
rect 31444 31968 31450 31980
rect 33137 31977 33149 31980
rect 33183 31977 33195 32011
rect 33137 31971 33195 31977
rect 33226 31968 33232 32020
rect 33284 32008 33290 32020
rect 33594 32008 33600 32020
rect 33284 31980 33600 32008
rect 33284 31968 33290 31980
rect 33594 31968 33600 31980
rect 33652 31968 33658 32020
rect 27157 31943 27215 31949
rect 27157 31909 27169 31943
rect 27203 31940 27215 31943
rect 27614 31940 27620 31952
rect 27203 31912 27620 31940
rect 27203 31909 27215 31912
rect 27157 31903 27215 31909
rect 27614 31900 27620 31912
rect 27672 31900 27678 31952
rect 27338 31832 27344 31884
rect 27396 31832 27402 31884
rect 27893 31875 27951 31881
rect 27893 31872 27905 31875
rect 27632 31844 27905 31872
rect 26789 31807 26847 31813
rect 26789 31773 26801 31807
rect 26835 31804 26847 31807
rect 27356 31804 27384 31832
rect 27632 31813 27660 31844
rect 27893 31841 27905 31844
rect 27939 31841 27951 31875
rect 27893 31835 27951 31841
rect 27982 31832 27988 31884
rect 28040 31872 28046 31884
rect 28040 31844 28396 31872
rect 28040 31832 28046 31844
rect 27433 31807 27491 31813
rect 27433 31804 27445 31807
rect 26835 31776 27445 31804
rect 26835 31773 26847 31776
rect 26789 31767 26847 31773
rect 27433 31773 27445 31776
rect 27479 31773 27491 31807
rect 27433 31767 27491 31773
rect 27525 31807 27583 31813
rect 27525 31773 27537 31807
rect 27571 31773 27583 31807
rect 27632 31807 27696 31813
rect 27632 31776 27650 31807
rect 27525 31767 27583 31773
rect 27638 31773 27650 31776
rect 27684 31773 27696 31807
rect 27798 31804 27804 31816
rect 27638 31767 27696 31773
rect 27724 31776 27804 31804
rect 17129 31739 17187 31745
rect 17129 31736 17141 31739
rect 16356 31708 16574 31736
rect 17107 31708 17141 31736
rect 16356 31696 16362 31708
rect 17129 31705 17141 31708
rect 17175 31705 17187 31739
rect 17129 31699 17187 31705
rect 17678 31696 17684 31748
rect 17736 31696 17742 31748
rect 19978 31696 19984 31748
rect 20036 31696 20042 31748
rect 21444 31739 21502 31745
rect 21444 31705 21456 31739
rect 21490 31736 21502 31739
rect 22002 31736 22008 31748
rect 21490 31708 22008 31736
rect 21490 31705 21502 31708
rect 21444 31699 21502 31705
rect 22002 31696 22008 31708
rect 22060 31696 22066 31748
rect 22094 31696 22100 31748
rect 22152 31736 22158 31748
rect 22554 31736 22560 31748
rect 22152 31708 22560 31736
rect 22152 31696 22158 31708
rect 22554 31696 22560 31708
rect 22612 31696 22618 31748
rect 26605 31739 26663 31745
rect 26605 31705 26617 31739
rect 26651 31736 26663 31739
rect 27065 31739 27123 31745
rect 27065 31736 27077 31739
rect 26651 31708 27077 31736
rect 26651 31705 26663 31708
rect 26605 31699 26663 31705
rect 27065 31705 27077 31708
rect 27111 31736 27123 31739
rect 27540 31736 27568 31767
rect 27111 31708 27568 31736
rect 27111 31705 27123 31708
rect 27065 31699 27123 31705
rect 15764 31640 16068 31668
rect 14461 31631 14519 31637
rect 16114 31628 16120 31680
rect 16172 31628 16178 31680
rect 18598 31628 18604 31680
rect 18656 31628 18662 31680
rect 22186 31628 22192 31680
rect 22244 31668 22250 31680
rect 22649 31671 22707 31677
rect 22649 31668 22661 31671
rect 22244 31640 22661 31668
rect 22244 31628 22250 31640
rect 22649 31637 22661 31640
rect 22695 31637 22707 31671
rect 22649 31631 22707 31637
rect 22830 31628 22836 31680
rect 22888 31668 22894 31680
rect 23385 31671 23443 31677
rect 23385 31668 23397 31671
rect 22888 31640 23397 31668
rect 22888 31628 22894 31640
rect 23385 31637 23397 31640
rect 23431 31637 23443 31671
rect 23385 31631 23443 31637
rect 24394 31628 24400 31680
rect 24452 31628 24458 31680
rect 26881 31671 26939 31677
rect 26881 31637 26893 31671
rect 26927 31668 26939 31671
rect 27724 31668 27752 31776
rect 27798 31764 27804 31776
rect 27856 31764 27862 31816
rect 28077 31807 28135 31813
rect 28077 31773 28089 31807
rect 28123 31804 28135 31807
rect 28258 31804 28264 31816
rect 28123 31776 28264 31804
rect 28123 31773 28135 31776
rect 28077 31767 28135 31773
rect 28258 31764 28264 31776
rect 28316 31764 28322 31816
rect 28368 31813 28396 31844
rect 30282 31832 30288 31884
rect 30340 31872 30346 31884
rect 30377 31875 30435 31881
rect 30377 31872 30389 31875
rect 30340 31844 30389 31872
rect 30340 31832 30346 31844
rect 30377 31841 30389 31844
rect 30423 31841 30435 31875
rect 30377 31835 30435 31841
rect 30650 31832 30656 31884
rect 30708 31832 30714 31884
rect 31846 31872 31852 31884
rect 31772 31844 31852 31872
rect 28353 31807 28411 31813
rect 28353 31773 28365 31807
rect 28399 31773 28411 31807
rect 28353 31767 28411 31773
rect 28626 31764 28632 31816
rect 28684 31764 28690 31816
rect 31772 31790 31800 31844
rect 31846 31832 31852 31844
rect 31904 31832 31910 31884
rect 32125 31875 32183 31881
rect 32125 31841 32137 31875
rect 32171 31841 32183 31875
rect 32125 31835 32183 31841
rect 32140 31804 32168 31835
rect 32401 31807 32459 31813
rect 32401 31804 32413 31807
rect 32140 31776 32413 31804
rect 32401 31773 32413 31776
rect 32447 31804 32459 31807
rect 32766 31804 32772 31816
rect 32447 31776 32772 31804
rect 32447 31773 32459 31776
rect 32401 31767 32459 31773
rect 32766 31764 32772 31776
rect 32824 31764 32830 31816
rect 32953 31807 33011 31813
rect 32953 31773 32965 31807
rect 32999 31804 33011 31807
rect 33045 31807 33103 31813
rect 33045 31804 33057 31807
rect 32999 31776 33057 31804
rect 32999 31773 33011 31776
rect 32953 31767 33011 31773
rect 33045 31773 33057 31776
rect 33091 31773 33103 31807
rect 33045 31767 33103 31773
rect 34698 31764 34704 31816
rect 34756 31804 34762 31816
rect 35529 31807 35587 31813
rect 35529 31804 35541 31807
rect 34756 31776 35541 31804
rect 34756 31764 34762 31776
rect 35529 31773 35541 31776
rect 35575 31773 35587 31807
rect 35529 31767 35587 31773
rect 36173 31807 36231 31813
rect 36173 31773 36185 31807
rect 36219 31804 36231 31807
rect 36630 31804 36636 31816
rect 36219 31776 36636 31804
rect 36219 31773 36231 31776
rect 36173 31767 36231 31773
rect 36630 31764 36636 31776
rect 36688 31764 36694 31816
rect 38470 31764 38476 31816
rect 38528 31764 38534 31816
rect 26927 31640 27752 31668
rect 28261 31671 28319 31677
rect 26927 31637 26939 31640
rect 26881 31631 26939 31637
rect 28261 31637 28273 31671
rect 28307 31668 28319 31671
rect 28350 31668 28356 31680
rect 28307 31640 28356 31668
rect 28307 31637 28319 31640
rect 28261 31631 28319 31637
rect 28350 31628 28356 31640
rect 28408 31628 28414 31680
rect 1104 31578 38824 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 38824 31578
rect 1104 31504 38824 31526
rect 3786 31424 3792 31476
rect 3844 31464 3850 31476
rect 3844 31436 4936 31464
rect 3844 31424 3850 31436
rect 4908 31396 4936 31436
rect 6730 31424 6736 31476
rect 6788 31424 6794 31476
rect 6822 31424 6828 31476
rect 6880 31464 6886 31476
rect 7742 31464 7748 31476
rect 6880 31436 7748 31464
rect 6880 31424 6886 31436
rect 7742 31424 7748 31436
rect 7800 31424 7806 31476
rect 12069 31467 12127 31473
rect 12069 31433 12081 31467
rect 12115 31464 12127 31467
rect 12434 31464 12440 31476
rect 12115 31436 12440 31464
rect 12115 31433 12127 31436
rect 12069 31427 12127 31433
rect 12434 31424 12440 31436
rect 12492 31424 12498 31476
rect 14090 31424 14096 31476
rect 14148 31464 14154 31476
rect 14829 31467 14887 31473
rect 14148 31436 14780 31464
rect 14148 31424 14154 31436
rect 5718 31396 5724 31408
rect 4830 31368 5724 31396
rect 5718 31356 5724 31368
rect 5776 31356 5782 31408
rect 6549 31399 6607 31405
rect 6549 31365 6561 31399
rect 6595 31396 6607 31399
rect 7190 31396 7196 31408
rect 6595 31368 7196 31396
rect 6595 31365 6607 31368
rect 6549 31359 6607 31365
rect 7190 31356 7196 31368
rect 7248 31356 7254 31408
rect 12618 31356 12624 31408
rect 12676 31396 12682 31408
rect 13354 31396 13360 31408
rect 12676 31368 13360 31396
rect 12676 31356 12682 31368
rect 13354 31356 13360 31368
rect 13412 31396 13418 31408
rect 14752 31396 14780 31436
rect 14829 31433 14841 31467
rect 14875 31464 14887 31467
rect 15194 31464 15200 31476
rect 14875 31436 15200 31464
rect 14875 31433 14887 31436
rect 14829 31427 14887 31433
rect 15194 31424 15200 31436
rect 15252 31424 15258 31476
rect 15286 31424 15292 31476
rect 15344 31424 15350 31476
rect 16206 31464 16212 31476
rect 15856 31436 16212 31464
rect 15856 31396 15884 31436
rect 16206 31424 16212 31436
rect 16264 31424 16270 31476
rect 17034 31424 17040 31476
rect 17092 31424 17098 31476
rect 18141 31467 18199 31473
rect 18141 31433 18153 31467
rect 18187 31464 18199 31467
rect 18230 31464 18236 31476
rect 18187 31436 18236 31464
rect 18187 31433 18199 31436
rect 18141 31427 18199 31433
rect 18230 31424 18236 31436
rect 18288 31424 18294 31476
rect 18598 31424 18604 31476
rect 18656 31424 18662 31476
rect 19978 31424 19984 31476
rect 20036 31424 20042 31476
rect 22002 31424 22008 31476
rect 22060 31464 22066 31476
rect 22465 31467 22523 31473
rect 22465 31464 22477 31467
rect 22060 31436 22477 31464
rect 22060 31424 22066 31436
rect 22465 31433 22477 31436
rect 22511 31433 22523 31467
rect 24305 31467 24363 31473
rect 22465 31427 22523 31433
rect 22572 31436 22968 31464
rect 16114 31396 16120 31408
rect 13412 31368 13846 31396
rect 14752 31368 15884 31396
rect 15948 31368 16120 31396
rect 13412 31356 13418 31368
rect 2222 31288 2228 31340
rect 2280 31328 2286 31340
rect 3329 31331 3387 31337
rect 3329 31328 3341 31331
rect 2280 31300 3341 31328
rect 2280 31288 2286 31300
rect 3329 31297 3341 31300
rect 3375 31297 3387 31331
rect 5810 31328 5816 31340
rect 3329 31291 3387 31297
rect 5092 31300 5816 31328
rect 3602 31220 3608 31272
rect 3660 31220 3666 31272
rect 5092 31269 5120 31300
rect 5810 31288 5816 31300
rect 5868 31288 5874 31340
rect 6638 31288 6644 31340
rect 6696 31328 6702 31340
rect 6822 31328 6828 31340
rect 6696 31300 6828 31328
rect 6696 31288 6702 31300
rect 6822 31288 6828 31300
rect 6880 31288 6886 31340
rect 7285 31331 7343 31337
rect 7285 31297 7297 31331
rect 7331 31328 7343 31331
rect 7558 31328 7564 31340
rect 7331 31300 7564 31328
rect 7331 31297 7343 31300
rect 7285 31291 7343 31297
rect 7558 31288 7564 31300
rect 7616 31288 7622 31340
rect 8110 31288 8116 31340
rect 8168 31288 8174 31340
rect 10965 31331 11023 31337
rect 10965 31297 10977 31331
rect 11011 31297 11023 31331
rect 10965 31291 11023 31297
rect 5077 31263 5135 31269
rect 5077 31229 5089 31263
rect 5123 31229 5135 31263
rect 5077 31223 5135 31229
rect 7374 31220 7380 31272
rect 7432 31220 7438 31272
rect 9217 31263 9275 31269
rect 9217 31260 9229 31263
rect 7668 31232 9229 31260
rect 4614 31152 4620 31204
rect 4672 31192 4678 31204
rect 5169 31195 5227 31201
rect 5169 31192 5181 31195
rect 4672 31164 5181 31192
rect 4672 31152 4678 31164
rect 5169 31161 5181 31164
rect 5215 31161 5227 31195
rect 5169 31155 5227 31161
rect 6917 31195 6975 31201
rect 6917 31161 6929 31195
rect 6963 31192 6975 31195
rect 7282 31192 7288 31204
rect 6963 31164 7288 31192
rect 6963 31161 6975 31164
rect 6917 31155 6975 31161
rect 7282 31152 7288 31164
rect 7340 31152 7346 31204
rect 7668 31201 7696 31232
rect 9217 31229 9229 31232
rect 9263 31229 9275 31263
rect 9217 31223 9275 31229
rect 9490 31220 9496 31272
rect 9548 31220 9554 31272
rect 10410 31220 10416 31272
rect 10468 31260 10474 31272
rect 10689 31263 10747 31269
rect 10689 31260 10701 31263
rect 10468 31232 10701 31260
rect 10468 31220 10474 31232
rect 10689 31229 10701 31232
rect 10735 31229 10747 31263
rect 10980 31260 11008 31291
rect 11698 31288 11704 31340
rect 11756 31288 11762 31340
rect 12342 31288 12348 31340
rect 12400 31328 12406 31340
rect 13078 31328 13084 31340
rect 12400 31300 13084 31328
rect 12400 31288 12406 31300
rect 13078 31288 13084 31300
rect 13136 31288 13142 31340
rect 15197 31331 15255 31337
rect 15197 31297 15209 31331
rect 15243 31297 15255 31331
rect 15197 31291 15255 31297
rect 15381 31331 15439 31337
rect 15381 31297 15393 31331
rect 15427 31328 15439 31331
rect 15948 31328 15976 31368
rect 16114 31356 16120 31368
rect 16172 31396 16178 31408
rect 17373 31399 17431 31405
rect 17373 31396 17385 31399
rect 16172 31368 17385 31396
rect 16172 31356 16178 31368
rect 15427 31300 15976 31328
rect 16025 31331 16083 31337
rect 15427 31297 15439 31300
rect 15381 31291 15439 31297
rect 16025 31297 16037 31331
rect 16071 31297 16083 31331
rect 16025 31291 16083 31297
rect 11146 31260 11152 31272
rect 10980 31232 11152 31260
rect 10689 31223 10747 31229
rect 11146 31220 11152 31232
rect 11204 31260 11210 31272
rect 11790 31260 11796 31272
rect 11204 31232 11796 31260
rect 11204 31220 11210 31232
rect 11790 31220 11796 31232
rect 11848 31220 11854 31272
rect 13357 31263 13415 31269
rect 13357 31229 13369 31263
rect 13403 31260 13415 31263
rect 14366 31260 14372 31272
rect 13403 31232 14372 31260
rect 13403 31229 13415 31232
rect 13357 31223 13415 31229
rect 14366 31220 14372 31232
rect 14424 31220 14430 31272
rect 15212 31260 15240 31291
rect 16040 31260 16068 31291
rect 16206 31288 16212 31340
rect 16264 31288 16270 31340
rect 16316 31337 16344 31368
rect 17373 31365 17385 31368
rect 17419 31365 17431 31399
rect 17373 31359 17431 31365
rect 17589 31399 17647 31405
rect 17589 31365 17601 31399
rect 17635 31396 17647 31399
rect 17678 31396 17684 31408
rect 17635 31368 17684 31396
rect 17635 31365 17647 31368
rect 17589 31359 17647 31365
rect 17678 31356 17684 31368
rect 17736 31356 17742 31408
rect 19996 31396 20024 31424
rect 19734 31368 20024 31396
rect 20070 31356 20076 31408
rect 20128 31396 20134 31408
rect 20165 31399 20223 31405
rect 20165 31396 20177 31399
rect 20128 31368 20177 31396
rect 20128 31356 20134 31368
rect 20165 31365 20177 31368
rect 20211 31365 20223 31399
rect 22572 31396 22600 31436
rect 20165 31359 20223 31365
rect 22480 31368 22600 31396
rect 16301 31331 16359 31337
rect 16301 31297 16313 31331
rect 16347 31297 16359 31331
rect 16301 31291 16359 31297
rect 16942 31288 16948 31340
rect 17000 31288 17006 31340
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 16114 31260 16120 31272
rect 15212 31232 16120 31260
rect 7653 31195 7711 31201
rect 7653 31161 7665 31195
rect 7699 31161 7711 31195
rect 7653 31155 7711 31161
rect 4798 31084 4804 31136
rect 4856 31124 4862 31136
rect 5442 31124 5448 31136
rect 4856 31096 5448 31124
rect 4856 31084 4862 31096
rect 5442 31084 5448 31096
rect 5500 31124 5506 31136
rect 6365 31127 6423 31133
rect 6365 31124 6377 31127
rect 5500 31096 6377 31124
rect 5500 31084 5506 31096
rect 6365 31093 6377 31096
rect 6411 31093 6423 31127
rect 6365 31087 6423 31093
rect 10134 31084 10140 31136
rect 10192 31124 10198 31136
rect 10781 31127 10839 31133
rect 10781 31124 10793 31127
rect 10192 31096 10793 31124
rect 10192 31084 10198 31096
rect 10781 31093 10793 31096
rect 10827 31093 10839 31127
rect 10781 31087 10839 31093
rect 10873 31127 10931 31133
rect 10873 31093 10885 31127
rect 10919 31124 10931 31127
rect 11238 31124 11244 31136
rect 10919 31096 11244 31124
rect 10919 31093 10931 31096
rect 10873 31087 10931 31093
rect 11238 31084 11244 31096
rect 11296 31084 11302 31136
rect 13906 31084 13912 31136
rect 13964 31124 13970 31136
rect 15212 31124 15240 31232
rect 16114 31220 16120 31232
rect 16172 31220 16178 31272
rect 16390 31220 16396 31272
rect 16448 31260 16454 31272
rect 17144 31260 17172 31291
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18138 31328 18144 31340
rect 18012 31300 18144 31328
rect 18012 31288 18018 31300
rect 18138 31288 18144 31300
rect 18196 31328 18202 31340
rect 18233 31331 18291 31337
rect 18233 31328 18245 31331
rect 18196 31300 18245 31328
rect 18196 31288 18202 31300
rect 18233 31297 18245 31300
rect 18279 31297 18291 31331
rect 18233 31291 18291 31297
rect 18417 31331 18475 31337
rect 18417 31297 18429 31331
rect 18463 31297 18475 31331
rect 18417 31291 18475 31297
rect 20441 31331 20499 31337
rect 20441 31297 20453 31331
rect 20487 31328 20499 31331
rect 20990 31328 20996 31340
rect 20487 31300 20996 31328
rect 20487 31297 20499 31300
rect 20441 31291 20499 31297
rect 16448 31232 17172 31260
rect 16448 31220 16454 31232
rect 17586 31220 17592 31272
rect 17644 31260 17650 31272
rect 17773 31263 17831 31269
rect 17773 31260 17785 31263
rect 17644 31232 17785 31260
rect 17644 31220 17650 31232
rect 17773 31229 17785 31232
rect 17819 31260 17831 31263
rect 18432 31260 18460 31291
rect 20990 31288 20996 31300
rect 21048 31288 21054 31340
rect 21818 31288 21824 31340
rect 21876 31288 21882 31340
rect 21910 31288 21916 31340
rect 21968 31328 21974 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21968 31300 22017 31328
rect 21968 31288 21974 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 22097 31331 22155 31337
rect 22097 31297 22109 31331
rect 22143 31297 22155 31331
rect 22097 31291 22155 31297
rect 18693 31263 18751 31269
rect 18693 31260 18705 31263
rect 17819 31232 18705 31260
rect 17819 31229 17831 31232
rect 17773 31223 17831 31229
rect 18693 31229 18705 31232
rect 18739 31229 18751 31263
rect 18693 31223 18751 31229
rect 21634 31152 21640 31204
rect 21692 31192 21698 31204
rect 22020 31192 22048 31291
rect 22112 31260 22140 31291
rect 22186 31288 22192 31340
rect 22244 31288 22250 31340
rect 22278 31260 22284 31272
rect 22112 31232 22284 31260
rect 22278 31220 22284 31232
rect 22336 31220 22342 31272
rect 22480 31192 22508 31368
rect 22830 31356 22836 31408
rect 22888 31356 22894 31408
rect 22940 31396 22968 31436
rect 24305 31433 24317 31467
rect 24351 31464 24363 31467
rect 24946 31464 24952 31476
rect 24351 31436 24952 31464
rect 24351 31433 24363 31436
rect 24305 31427 24363 31433
rect 24946 31424 24952 31436
rect 25004 31424 25010 31476
rect 25038 31424 25044 31476
rect 25096 31424 25102 31476
rect 28258 31424 28264 31476
rect 28316 31464 28322 31476
rect 29089 31467 29147 31473
rect 29089 31464 29101 31467
rect 28316 31436 29101 31464
rect 28316 31424 28322 31436
rect 29089 31433 29101 31436
rect 29135 31433 29147 31467
rect 29089 31427 29147 31433
rect 36630 31424 36636 31476
rect 36688 31424 36694 31476
rect 26234 31396 26240 31408
rect 22940 31368 23322 31396
rect 26082 31368 26240 31396
rect 26234 31356 26240 31368
rect 26292 31396 26298 31408
rect 26292 31368 26924 31396
rect 26292 31356 26298 31368
rect 22554 31288 22560 31340
rect 22612 31288 22618 31340
rect 24486 31288 24492 31340
rect 24544 31288 24550 31340
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 24596 31260 24624 31291
rect 26418 31260 26424 31272
rect 24596 31232 26424 31260
rect 26418 31220 26424 31232
rect 26476 31220 26482 31272
rect 26513 31263 26571 31269
rect 26513 31229 26525 31263
rect 26559 31260 26571 31263
rect 26559 31232 26740 31260
rect 26559 31229 26571 31232
rect 26513 31223 26571 31229
rect 21692 31164 22508 31192
rect 26712 31192 26740 31232
rect 26786 31220 26792 31272
rect 26844 31220 26850 31272
rect 26896 31260 26924 31368
rect 27614 31356 27620 31408
rect 27672 31356 27678 31408
rect 28350 31356 28356 31408
rect 28408 31356 28414 31408
rect 34606 31356 34612 31408
rect 34664 31396 34670 31408
rect 35161 31399 35219 31405
rect 35161 31396 35173 31399
rect 34664 31368 35173 31396
rect 34664 31356 34670 31368
rect 35161 31365 35173 31368
rect 35207 31365 35219 31399
rect 35161 31359 35219 31365
rect 36170 31356 36176 31408
rect 36228 31356 36234 31408
rect 27338 31288 27344 31340
rect 27396 31288 27402 31340
rect 32766 31288 32772 31340
rect 32824 31288 32830 31340
rect 32953 31331 33011 31337
rect 32953 31297 32965 31331
rect 32999 31328 33011 31331
rect 33134 31328 33140 31340
rect 32999 31300 33140 31328
rect 32999 31297 33011 31300
rect 32953 31291 33011 31297
rect 33134 31288 33140 31300
rect 33192 31328 33198 31340
rect 33502 31328 33508 31340
rect 33192 31300 33508 31328
rect 33192 31288 33198 31300
rect 33502 31288 33508 31300
rect 33560 31288 33566 31340
rect 28350 31260 28356 31272
rect 26896 31232 28356 31260
rect 28350 31220 28356 31232
rect 28408 31220 28414 31272
rect 31754 31220 31760 31272
rect 31812 31260 31818 31272
rect 33965 31263 34023 31269
rect 33965 31260 33977 31263
rect 31812 31232 33977 31260
rect 31812 31220 31818 31232
rect 33965 31229 33977 31232
rect 34011 31229 34023 31263
rect 33965 31223 34023 31229
rect 34241 31263 34299 31269
rect 34241 31229 34253 31263
rect 34287 31260 34299 31263
rect 34422 31260 34428 31272
rect 34287 31232 34428 31260
rect 34287 31229 34299 31232
rect 34241 31223 34299 31229
rect 34422 31220 34428 31232
rect 34480 31220 34486 31272
rect 34885 31263 34943 31269
rect 34885 31229 34897 31263
rect 34931 31229 34943 31263
rect 34885 31223 34943 31229
rect 26970 31192 26976 31204
rect 26712 31164 26976 31192
rect 21692 31152 21698 31164
rect 26970 31152 26976 31164
rect 27028 31152 27034 31204
rect 13964 31096 15240 31124
rect 13964 31084 13970 31096
rect 15746 31084 15752 31136
rect 15804 31124 15810 31136
rect 16025 31127 16083 31133
rect 16025 31124 16037 31127
rect 15804 31096 16037 31124
rect 15804 31084 15810 31096
rect 16025 31093 16037 31096
rect 16071 31093 16083 31127
rect 16025 31087 16083 31093
rect 16666 31084 16672 31136
rect 16724 31124 16730 31136
rect 17221 31127 17279 31133
rect 17221 31124 17233 31127
rect 16724 31096 17233 31124
rect 16724 31084 16730 31096
rect 17221 31093 17233 31096
rect 17267 31093 17279 31127
rect 17221 31087 17279 31093
rect 17402 31084 17408 31136
rect 17460 31084 17466 31136
rect 24765 31127 24823 31133
rect 24765 31093 24777 31127
rect 24811 31124 24823 31127
rect 24854 31124 24860 31136
rect 24811 31096 24860 31124
rect 24811 31093 24823 31096
rect 24765 31087 24823 31093
rect 24854 31084 24860 31096
rect 24912 31084 24918 31136
rect 29914 31084 29920 31136
rect 29972 31084 29978 31136
rect 30466 31084 30472 31136
rect 30524 31084 30530 31136
rect 32582 31084 32588 31136
rect 32640 31084 32646 31136
rect 32953 31127 33011 31133
rect 32953 31093 32965 31127
rect 32999 31124 33011 31127
rect 33134 31124 33140 31136
rect 32999 31096 33140 31124
rect 32999 31093 33011 31096
rect 32953 31087 33011 31093
rect 33134 31084 33140 31096
rect 33192 31124 33198 31136
rect 33410 31124 33416 31136
rect 33192 31096 33416 31124
rect 33192 31084 33198 31096
rect 33410 31084 33416 31096
rect 33468 31084 33474 31136
rect 34900 31124 34928 31223
rect 35342 31124 35348 31136
rect 34900 31096 35348 31124
rect 35342 31084 35348 31096
rect 35400 31084 35406 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 3602 30880 3608 30932
rect 3660 30920 3666 30932
rect 3881 30923 3939 30929
rect 3881 30920 3893 30923
rect 3660 30892 3893 30920
rect 3660 30880 3666 30892
rect 3881 30889 3893 30892
rect 3927 30889 3939 30923
rect 3881 30883 3939 30889
rect 6730 30880 6736 30932
rect 6788 30880 6794 30932
rect 7285 30923 7343 30929
rect 7285 30889 7297 30923
rect 7331 30920 7343 30923
rect 7374 30920 7380 30932
rect 7331 30892 7380 30920
rect 7331 30889 7343 30892
rect 7285 30883 7343 30889
rect 7374 30880 7380 30892
rect 7432 30880 7438 30932
rect 11790 30880 11796 30932
rect 11848 30920 11854 30932
rect 12437 30923 12495 30929
rect 12437 30920 12449 30923
rect 11848 30892 12449 30920
rect 11848 30880 11854 30892
rect 12437 30889 12449 30892
rect 12483 30889 12495 30923
rect 14090 30920 14096 30932
rect 12437 30883 12495 30889
rect 13372 30892 14096 30920
rect 4798 30812 4804 30864
rect 4856 30812 4862 30864
rect 4816 30784 4844 30812
rect 4448 30756 4844 30784
rect 5261 30787 5319 30793
rect 3881 30719 3939 30725
rect 3881 30685 3893 30719
rect 3927 30685 3939 30719
rect 3881 30679 3939 30685
rect 3896 30648 3924 30679
rect 4062 30676 4068 30728
rect 4120 30676 4126 30728
rect 4448 30725 4476 30756
rect 5261 30753 5273 30787
rect 5307 30784 5319 30787
rect 5350 30784 5356 30796
rect 5307 30756 5356 30784
rect 5307 30753 5319 30756
rect 5261 30747 5319 30753
rect 5350 30744 5356 30756
rect 5408 30744 5414 30796
rect 7392 30784 7420 30880
rect 7469 30787 7527 30793
rect 7469 30784 7481 30787
rect 7392 30756 7481 30784
rect 7469 30753 7481 30756
rect 7515 30753 7527 30787
rect 7469 30747 7527 30753
rect 9490 30744 9496 30796
rect 9548 30784 9554 30796
rect 9861 30787 9919 30793
rect 9861 30784 9873 30787
rect 9548 30756 9873 30784
rect 9548 30744 9554 30756
rect 9861 30753 9873 30756
rect 9907 30784 9919 30787
rect 11146 30784 11152 30796
rect 9907 30756 11152 30784
rect 9907 30753 9919 30756
rect 9861 30747 9919 30753
rect 11146 30744 11152 30756
rect 11204 30744 11210 30796
rect 11609 30787 11667 30793
rect 11609 30753 11621 30787
rect 11655 30784 11667 30787
rect 12253 30787 12311 30793
rect 12253 30784 12265 30787
rect 11655 30756 12265 30784
rect 11655 30753 11667 30756
rect 11609 30747 11667 30753
rect 12253 30753 12265 30756
rect 12299 30784 12311 30787
rect 12805 30787 12863 30793
rect 12805 30784 12817 30787
rect 12299 30756 12817 30784
rect 12299 30753 12311 30756
rect 12253 30747 12311 30753
rect 12805 30753 12817 30756
rect 12851 30753 12863 30787
rect 12805 30747 12863 30753
rect 4433 30719 4491 30725
rect 4433 30685 4445 30719
rect 4479 30685 4491 30719
rect 4433 30679 4491 30685
rect 4614 30676 4620 30728
rect 4672 30676 4678 30728
rect 4798 30676 4804 30728
rect 4856 30716 4862 30728
rect 4985 30719 5043 30725
rect 4985 30716 4997 30719
rect 4856 30688 4997 30716
rect 4856 30676 4862 30688
rect 4985 30685 4997 30688
rect 5031 30685 5043 30719
rect 4985 30679 5043 30685
rect 7190 30676 7196 30728
rect 7248 30676 7254 30728
rect 7374 30676 7380 30728
rect 7432 30676 7438 30728
rect 7650 30676 7656 30728
rect 7708 30676 7714 30728
rect 12618 30676 12624 30728
rect 12676 30676 12682 30728
rect 13372 30725 13400 30892
rect 14090 30880 14096 30892
rect 14148 30880 14154 30932
rect 15933 30923 15991 30929
rect 15933 30889 15945 30923
rect 15979 30920 15991 30923
rect 16022 30920 16028 30932
rect 15979 30892 16028 30920
rect 15979 30889 15991 30892
rect 15933 30883 15991 30889
rect 16022 30880 16028 30892
rect 16080 30880 16086 30932
rect 16114 30880 16120 30932
rect 16172 30880 16178 30932
rect 16298 30880 16304 30932
rect 16356 30920 16362 30932
rect 16942 30920 16948 30932
rect 16356 30892 16948 30920
rect 16356 30880 16362 30892
rect 16942 30880 16948 30892
rect 17000 30880 17006 30932
rect 23566 30880 23572 30932
rect 23624 30880 23630 30932
rect 26970 30880 26976 30932
rect 27028 30880 27034 30932
rect 31754 30880 31760 30932
rect 31812 30920 31818 30932
rect 32217 30923 32275 30929
rect 32217 30920 32229 30923
rect 31812 30892 32229 30920
rect 31812 30880 31818 30892
rect 32217 30889 32229 30892
rect 32263 30889 32275 30923
rect 32217 30883 32275 30889
rect 33318 30880 33324 30932
rect 33376 30920 33382 30932
rect 33413 30923 33471 30929
rect 33413 30920 33425 30923
rect 33376 30892 33425 30920
rect 33376 30880 33382 30892
rect 33413 30889 33425 30892
rect 33459 30889 33471 30923
rect 33413 30883 33471 30889
rect 33781 30923 33839 30929
rect 33781 30889 33793 30923
rect 33827 30920 33839 30923
rect 33870 30920 33876 30932
rect 33827 30892 33876 30920
rect 33827 30889 33839 30892
rect 33781 30883 33839 30889
rect 33870 30880 33876 30892
rect 33928 30880 33934 30932
rect 33965 30923 34023 30929
rect 33965 30889 33977 30923
rect 34011 30920 34023 30923
rect 34238 30920 34244 30932
rect 34011 30892 34244 30920
rect 34011 30889 34023 30892
rect 33965 30883 34023 30889
rect 34238 30880 34244 30892
rect 34296 30880 34302 30932
rect 35069 30923 35127 30929
rect 35069 30889 35081 30923
rect 35115 30889 35127 30923
rect 35069 30883 35127 30889
rect 13909 30855 13967 30861
rect 13909 30821 13921 30855
rect 13955 30821 13967 30855
rect 13909 30815 13967 30821
rect 15473 30855 15531 30861
rect 15473 30821 15485 30855
rect 15519 30821 15531 30855
rect 15473 30815 15531 30821
rect 13924 30784 13952 30815
rect 14642 30784 14648 30796
rect 13924 30756 14412 30784
rect 13357 30719 13415 30725
rect 13357 30685 13369 30719
rect 13403 30685 13415 30719
rect 13357 30679 13415 30685
rect 13541 30719 13599 30725
rect 13541 30685 13553 30719
rect 13587 30716 13599 30719
rect 13630 30716 13636 30728
rect 13587 30688 13636 30716
rect 13587 30685 13599 30688
rect 13541 30679 13599 30685
rect 13630 30676 13636 30688
rect 13688 30676 13694 30728
rect 14384 30725 14412 30756
rect 14476 30756 14648 30784
rect 13725 30719 13783 30725
rect 13725 30685 13737 30719
rect 13771 30716 13783 30719
rect 14369 30719 14427 30725
rect 13771 30688 14320 30716
rect 13771 30685 13783 30688
rect 13725 30679 13783 30685
rect 4525 30651 4583 30657
rect 4525 30648 4537 30651
rect 3896 30620 4537 30648
rect 4525 30617 4537 30620
rect 4571 30617 4583 30651
rect 4525 30611 4583 30617
rect 5718 30608 5724 30660
rect 5776 30608 5782 30660
rect 10134 30608 10140 30660
rect 10192 30608 10198 30660
rect 10226 30608 10232 30660
rect 10284 30648 10290 30660
rect 13449 30651 13507 30657
rect 10284 30620 10626 30648
rect 10284 30608 10290 30620
rect 13449 30617 13461 30651
rect 13495 30648 13507 30651
rect 13495 30620 13860 30648
rect 13495 30617 13507 30620
rect 13449 30611 13507 30617
rect 7837 30583 7895 30589
rect 7837 30549 7849 30583
rect 7883 30580 7895 30583
rect 9030 30580 9036 30592
rect 7883 30552 9036 30580
rect 7883 30549 7895 30552
rect 7837 30543 7895 30549
rect 9030 30540 9036 30552
rect 9088 30540 9094 30592
rect 9766 30540 9772 30592
rect 9824 30580 9830 30592
rect 10244 30580 10272 30608
rect 9824 30552 10272 30580
rect 9824 30540 9830 30552
rect 11698 30540 11704 30592
rect 11756 30540 11762 30592
rect 13832 30580 13860 30620
rect 13906 30608 13912 30660
rect 13964 30608 13970 30660
rect 13998 30608 14004 30660
rect 14056 30648 14062 30660
rect 14185 30651 14243 30657
rect 14185 30648 14197 30651
rect 14056 30620 14197 30648
rect 14056 30608 14062 30620
rect 14185 30617 14197 30620
rect 14231 30617 14243 30651
rect 14292 30648 14320 30688
rect 14369 30685 14381 30719
rect 14415 30685 14427 30719
rect 14369 30679 14427 30685
rect 14476 30648 14504 30756
rect 14642 30744 14648 30756
rect 14700 30744 14706 30796
rect 15194 30744 15200 30796
rect 15252 30744 15258 30796
rect 15488 30784 15516 30815
rect 16206 30812 16212 30864
rect 16264 30852 16270 30864
rect 17218 30852 17224 30864
rect 16264 30824 17224 30852
rect 16264 30812 16270 30824
rect 17218 30812 17224 30824
rect 17276 30852 17282 30864
rect 17678 30852 17684 30864
rect 17276 30824 17684 30852
rect 17276 30812 17282 30824
rect 17328 30793 17356 30824
rect 17678 30812 17684 30824
rect 17736 30812 17742 30864
rect 22094 30812 22100 30864
rect 22152 30852 22158 30864
rect 22465 30855 22523 30861
rect 22465 30852 22477 30855
rect 22152 30824 22477 30852
rect 22152 30812 22158 30824
rect 22465 30821 22477 30824
rect 22511 30852 22523 30855
rect 24854 30852 24860 30864
rect 22511 30824 23980 30852
rect 22511 30821 22523 30824
rect 22465 30815 22523 30821
rect 17313 30787 17371 30793
rect 15488 30756 16804 30784
rect 14550 30676 14556 30728
rect 14608 30676 14614 30728
rect 14829 30719 14887 30725
rect 14829 30685 14841 30719
rect 14875 30716 14887 30719
rect 15010 30716 15016 30728
rect 14875 30688 15016 30716
rect 14875 30685 14887 30688
rect 14829 30679 14887 30685
rect 15010 30676 15016 30688
rect 15068 30676 15074 30728
rect 15746 30676 15752 30728
rect 15804 30676 15810 30728
rect 16025 30719 16083 30725
rect 16025 30685 16037 30719
rect 16071 30716 16083 30719
rect 16669 30719 16727 30725
rect 16669 30716 16681 30719
rect 16071 30688 16681 30716
rect 16071 30685 16083 30688
rect 16025 30679 16083 30685
rect 16669 30685 16681 30688
rect 16715 30685 16727 30719
rect 16776 30716 16804 30756
rect 17313 30753 17325 30787
rect 17359 30753 17371 30787
rect 17313 30747 17371 30753
rect 20990 30744 20996 30796
rect 21048 30784 21054 30796
rect 21085 30787 21143 30793
rect 21085 30784 21097 30787
rect 21048 30756 21097 30784
rect 21048 30744 21054 30756
rect 21085 30753 21097 30756
rect 21131 30753 21143 30787
rect 21085 30747 21143 30753
rect 17957 30719 18015 30725
rect 17957 30716 17969 30719
rect 16776 30688 17969 30716
rect 16669 30679 16727 30685
rect 17957 30685 17969 30688
rect 18003 30685 18015 30719
rect 17957 30679 18015 30685
rect 18138 30676 18144 30728
rect 18196 30676 18202 30728
rect 23750 30676 23756 30728
rect 23808 30676 23814 30728
rect 23842 30676 23848 30728
rect 23900 30676 23906 30728
rect 23952 30725 23980 30824
rect 24044 30824 24860 30852
rect 24044 30725 24072 30824
rect 24854 30812 24860 30824
rect 24912 30812 24918 30864
rect 26145 30855 26203 30861
rect 26145 30821 26157 30855
rect 26191 30852 26203 30855
rect 26191 30824 26372 30852
rect 26191 30821 26203 30824
rect 26145 30815 26203 30821
rect 24213 30787 24271 30793
rect 24213 30753 24225 30787
rect 24259 30784 24271 30787
rect 24394 30784 24400 30796
rect 24259 30756 24400 30784
rect 24259 30753 24271 30756
rect 24213 30747 24271 30753
rect 23937 30719 23995 30725
rect 23937 30685 23949 30719
rect 23983 30685 23995 30719
rect 24044 30719 24113 30725
rect 24044 30688 24067 30719
rect 23937 30679 23995 30685
rect 24055 30685 24067 30688
rect 24101 30685 24113 30719
rect 24055 30679 24113 30685
rect 14292 30620 14504 30648
rect 14185 30611 14243 30617
rect 15286 30608 15292 30660
rect 15344 30657 15350 30660
rect 15344 30651 15372 30657
rect 15360 30617 15372 30651
rect 15344 30611 15372 30617
rect 15488 30620 16252 30648
rect 15344 30608 15350 30611
rect 14090 30580 14096 30592
rect 13832 30552 14096 30580
rect 14090 30540 14096 30552
rect 14148 30540 14154 30592
rect 15105 30583 15163 30589
rect 15105 30549 15117 30583
rect 15151 30580 15163 30583
rect 15488 30580 15516 30620
rect 15151 30552 15516 30580
rect 15565 30583 15623 30589
rect 15151 30549 15163 30552
rect 15105 30543 15163 30549
rect 15565 30549 15577 30583
rect 15611 30580 15623 30583
rect 15746 30580 15752 30592
rect 15611 30552 15752 30580
rect 15611 30549 15623 30552
rect 15565 30543 15623 30549
rect 15746 30540 15752 30552
rect 15804 30540 15810 30592
rect 16224 30580 16252 30620
rect 16298 30608 16304 30660
rect 16356 30608 16362 30660
rect 16390 30608 16396 30660
rect 16448 30648 16454 30660
rect 16485 30651 16543 30657
rect 16485 30648 16497 30651
rect 16448 30620 16497 30648
rect 16448 30608 16454 30620
rect 16485 30617 16497 30620
rect 16531 30617 16543 30651
rect 16485 30611 16543 30617
rect 16574 30608 16580 30660
rect 16632 30648 16638 30660
rect 17497 30651 17555 30657
rect 17497 30648 17509 30651
rect 16632 30620 17509 30648
rect 16632 30608 16638 30620
rect 17497 30617 17509 30620
rect 17543 30617 17555 30651
rect 17497 30611 17555 30617
rect 17310 30580 17316 30592
rect 16224 30552 17316 30580
rect 17310 30540 17316 30552
rect 17368 30540 17374 30592
rect 17512 30580 17540 30611
rect 17862 30608 17868 30660
rect 17920 30608 17926 30660
rect 18325 30651 18383 30657
rect 18325 30617 18337 30651
rect 18371 30648 18383 30651
rect 18782 30648 18788 30660
rect 18371 30620 18788 30648
rect 18371 30617 18383 30620
rect 18325 30611 18383 30617
rect 18782 30608 18788 30620
rect 18840 30608 18846 30660
rect 21358 30657 21364 30660
rect 21352 30611 21364 30657
rect 21358 30608 21364 30611
rect 21416 30608 21422 30660
rect 22738 30608 22744 30660
rect 22796 30608 22802 30660
rect 18417 30583 18475 30589
rect 18417 30580 18429 30583
rect 17512 30552 18429 30580
rect 18417 30549 18429 30552
rect 18463 30549 18475 30583
rect 18417 30543 18475 30549
rect 22278 30540 22284 30592
rect 22336 30580 22342 30592
rect 22646 30580 22652 30592
rect 22336 30552 22652 30580
rect 22336 30540 22342 30552
rect 22646 30540 22652 30552
rect 22704 30580 22710 30592
rect 22833 30583 22891 30589
rect 22833 30580 22845 30583
rect 22704 30552 22845 30580
rect 22704 30540 22710 30552
rect 22833 30549 22845 30552
rect 22879 30549 22891 30583
rect 22833 30543 22891 30549
rect 23474 30540 23480 30592
rect 23532 30580 23538 30592
rect 24228 30580 24256 30747
rect 24394 30744 24400 30756
rect 24452 30744 24458 30796
rect 24872 30784 24900 30812
rect 25222 30784 25228 30796
rect 24872 30756 25228 30784
rect 25222 30744 25228 30756
rect 25280 30784 25286 30796
rect 26344 30793 26372 30824
rect 32766 30812 32772 30864
rect 32824 30812 32830 30864
rect 33888 30852 33916 30880
rect 34701 30855 34759 30861
rect 34701 30852 34713 30855
rect 33888 30824 34713 30852
rect 34701 30821 34713 30824
rect 34747 30821 34759 30855
rect 34701 30815 34759 30821
rect 26329 30787 26387 30793
rect 25280 30756 25820 30784
rect 25280 30744 25286 30756
rect 25406 30676 25412 30728
rect 25464 30676 25470 30728
rect 25590 30676 25596 30728
rect 25648 30676 25654 30728
rect 25792 30725 25820 30756
rect 26329 30753 26341 30787
rect 26375 30753 26387 30787
rect 26329 30747 26387 30753
rect 29641 30787 29699 30793
rect 29641 30753 29653 30787
rect 29687 30784 29699 30787
rect 30282 30784 30288 30796
rect 29687 30756 30288 30784
rect 29687 30753 29699 30756
rect 29641 30747 29699 30753
rect 30282 30744 30288 30756
rect 30340 30744 30346 30796
rect 31389 30787 31447 30793
rect 31389 30753 31401 30787
rect 31435 30784 31447 30787
rect 32493 30787 32551 30793
rect 32493 30784 32505 30787
rect 31435 30756 32168 30784
rect 31435 30753 31447 30756
rect 31389 30747 31447 30753
rect 25777 30719 25835 30725
rect 25777 30685 25789 30719
rect 25823 30685 25835 30719
rect 25777 30679 25835 30685
rect 25958 30676 25964 30728
rect 26016 30676 26022 30728
rect 32140 30660 32168 30756
rect 32416 30756 32505 30784
rect 32306 30676 32312 30728
rect 32364 30676 32370 30728
rect 32416 30725 32444 30756
rect 32493 30753 32505 30756
rect 32539 30753 32551 30787
rect 32784 30784 32812 30812
rect 32784 30756 32996 30784
rect 32493 30747 32551 30753
rect 32401 30719 32459 30725
rect 32401 30685 32413 30719
rect 32447 30685 32459 30719
rect 32401 30679 32459 30685
rect 32769 30719 32827 30725
rect 32769 30685 32781 30719
rect 32815 30685 32827 30719
rect 32769 30679 32827 30685
rect 24397 30651 24455 30657
rect 24397 30617 24409 30651
rect 24443 30648 24455 30651
rect 24486 30648 24492 30660
rect 24443 30620 24492 30648
rect 24443 30617 24455 30620
rect 24397 30611 24455 30617
rect 24486 30608 24492 30620
rect 24544 30608 24550 30660
rect 24578 30608 24584 30660
rect 24636 30608 24642 30660
rect 24765 30651 24823 30657
rect 24765 30617 24777 30651
rect 24811 30648 24823 30651
rect 25222 30648 25228 30660
rect 24811 30620 25228 30648
rect 24811 30617 24823 30620
rect 24765 30611 24823 30617
rect 25222 30608 25228 30620
rect 25280 30608 25286 30660
rect 25869 30651 25927 30657
rect 25869 30617 25881 30651
rect 25915 30648 25927 30651
rect 26050 30648 26056 30660
rect 25915 30620 26056 30648
rect 25915 30617 25927 30620
rect 25869 30611 25927 30617
rect 26050 30608 26056 30620
rect 26108 30608 26114 30660
rect 29914 30608 29920 30660
rect 29972 30608 29978 30660
rect 31846 30648 31852 30660
rect 31142 30620 31852 30648
rect 31846 30608 31852 30620
rect 31904 30608 31910 30660
rect 32122 30608 32128 30660
rect 32180 30608 32186 30660
rect 32784 30648 32812 30679
rect 32858 30676 32864 30728
rect 32916 30676 32922 30728
rect 32968 30725 32996 30756
rect 33502 30744 33508 30796
rect 33560 30744 33566 30796
rect 33962 30744 33968 30796
rect 34020 30784 34026 30796
rect 34333 30787 34391 30793
rect 34333 30784 34345 30787
rect 34020 30756 34345 30784
rect 34020 30744 34026 30756
rect 34333 30753 34345 30756
rect 34379 30753 34391 30787
rect 34333 30747 34391 30753
rect 34422 30744 34428 30796
rect 34480 30784 34486 30796
rect 34517 30787 34575 30793
rect 34517 30784 34529 30787
rect 34480 30756 34529 30784
rect 34480 30744 34486 30756
rect 34517 30753 34529 30756
rect 34563 30784 34575 30787
rect 35084 30784 35112 30883
rect 35986 30784 35992 30796
rect 34563 30756 35112 30784
rect 35176 30756 35992 30784
rect 34563 30753 34575 30756
rect 34517 30747 34575 30753
rect 32953 30719 33011 30725
rect 32953 30685 32965 30719
rect 32999 30685 33011 30719
rect 32953 30679 33011 30685
rect 33134 30676 33140 30728
rect 33192 30676 33198 30728
rect 33226 30676 33232 30728
rect 33284 30716 33290 30728
rect 33413 30719 33471 30725
rect 33413 30716 33425 30719
rect 33284 30688 33425 30716
rect 33284 30676 33290 30688
rect 33413 30685 33425 30688
rect 33459 30716 33471 30719
rect 33459 30688 33640 30716
rect 33459 30685 33471 30688
rect 33413 30679 33471 30685
rect 32784 30620 33272 30648
rect 23532 30552 24256 30580
rect 23532 30540 23538 30552
rect 24854 30540 24860 30592
rect 24912 30540 24918 30592
rect 33244 30589 33272 30620
rect 33229 30583 33287 30589
rect 33229 30549 33241 30583
rect 33275 30549 33287 30583
rect 33612 30580 33640 30688
rect 33686 30676 33692 30728
rect 33744 30716 33750 30728
rect 34238 30716 34244 30728
rect 33744 30688 34244 30716
rect 33744 30676 33750 30688
rect 34238 30676 34244 30688
rect 34296 30676 34302 30728
rect 34149 30651 34207 30657
rect 34149 30648 34161 30651
rect 33888 30620 34161 30648
rect 33888 30580 33916 30620
rect 34149 30617 34161 30620
rect 34195 30648 34207 30651
rect 35176 30648 35204 30756
rect 35986 30744 35992 30756
rect 36044 30744 36050 30796
rect 35342 30676 35348 30728
rect 35400 30676 35406 30728
rect 38470 30676 38476 30728
rect 38528 30676 38534 30728
rect 35621 30651 35679 30657
rect 35621 30648 35633 30651
rect 34195 30620 35204 30648
rect 35268 30620 35633 30648
rect 34195 30617 34207 30620
rect 34149 30611 34207 30617
rect 33962 30589 33968 30592
rect 33612 30552 33916 30580
rect 33944 30583 33968 30589
rect 33229 30543 33287 30549
rect 33944 30549 33956 30583
rect 33944 30543 33968 30549
rect 33962 30540 33968 30543
rect 34020 30540 34026 30592
rect 34514 30540 34520 30592
rect 34572 30540 34578 30592
rect 35066 30540 35072 30592
rect 35124 30540 35130 30592
rect 35268 30589 35296 30620
rect 35621 30617 35633 30620
rect 35667 30617 35679 30651
rect 35621 30611 35679 30617
rect 36078 30608 36084 30660
rect 36136 30608 36142 30660
rect 35253 30583 35311 30589
rect 35253 30549 35265 30583
rect 35299 30549 35311 30583
rect 35253 30543 35311 30549
rect 37093 30583 37151 30589
rect 37093 30549 37105 30583
rect 37139 30580 37151 30583
rect 37182 30580 37188 30592
rect 37139 30552 37188 30580
rect 37139 30549 37151 30552
rect 37093 30543 37151 30549
rect 37182 30540 37188 30552
rect 37240 30540 37246 30592
rect 1104 30490 38824 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 38824 30490
rect 1104 30416 38824 30438
rect 4062 30336 4068 30388
rect 4120 30336 4126 30388
rect 7374 30336 7380 30388
rect 7432 30376 7438 30388
rect 7561 30379 7619 30385
rect 7561 30376 7573 30379
rect 7432 30348 7573 30376
rect 7432 30336 7438 30348
rect 7561 30345 7573 30348
rect 7607 30345 7619 30379
rect 7561 30339 7619 30345
rect 14642 30336 14648 30388
rect 14700 30376 14706 30388
rect 14829 30379 14887 30385
rect 14829 30376 14841 30379
rect 14700 30348 14841 30376
rect 14700 30336 14706 30348
rect 14829 30345 14841 30348
rect 14875 30345 14887 30379
rect 14829 30339 14887 30345
rect 16117 30379 16175 30385
rect 16117 30345 16129 30379
rect 16163 30376 16175 30379
rect 16206 30376 16212 30388
rect 16163 30348 16212 30376
rect 16163 30345 16175 30348
rect 16117 30339 16175 30345
rect 16206 30336 16212 30348
rect 16264 30336 16270 30388
rect 17313 30379 17371 30385
rect 17313 30345 17325 30379
rect 17359 30376 17371 30379
rect 17402 30376 17408 30388
rect 17359 30348 17408 30376
rect 17359 30345 17371 30348
rect 17313 30339 17371 30345
rect 4080 30308 4108 30336
rect 5169 30311 5227 30317
rect 5169 30308 5181 30311
rect 4080 30280 5181 30308
rect 5169 30277 5181 30280
rect 5215 30277 5227 30311
rect 5169 30271 5227 30277
rect 8018 30268 8024 30320
rect 8076 30268 8082 30320
rect 9030 30268 9036 30320
rect 9088 30268 9094 30320
rect 10229 30311 10287 30317
rect 10229 30308 10241 30311
rect 9600 30280 10241 30308
rect 3786 30200 3792 30252
rect 3844 30240 3850 30252
rect 4065 30243 4123 30249
rect 4065 30240 4077 30243
rect 3844 30212 4077 30240
rect 3844 30200 3850 30212
rect 4065 30209 4077 30212
rect 4111 30209 4123 30243
rect 4065 30203 4123 30209
rect 5353 30243 5411 30249
rect 5353 30209 5365 30243
rect 5399 30240 5411 30243
rect 5442 30240 5448 30252
rect 5399 30212 5448 30240
rect 5399 30209 5411 30212
rect 5353 30203 5411 30209
rect 5442 30200 5448 30212
rect 5500 30200 5506 30252
rect 5537 30243 5595 30249
rect 5537 30209 5549 30243
rect 5583 30240 5595 30243
rect 5810 30240 5816 30252
rect 5583 30212 5816 30240
rect 5583 30209 5595 30212
rect 5537 30203 5595 30209
rect 5810 30200 5816 30212
rect 5868 30200 5874 30252
rect 6822 30200 6828 30252
rect 6880 30200 6886 30252
rect 9309 30243 9367 30249
rect 9309 30209 9321 30243
rect 9355 30240 9367 30243
rect 9490 30240 9496 30252
rect 9355 30212 9496 30240
rect 9355 30209 9367 30212
rect 9309 30203 9367 30209
rect 9490 30200 9496 30212
rect 9548 30200 9554 30252
rect 9600 30249 9628 30280
rect 10229 30277 10241 30280
rect 10275 30277 10287 30311
rect 10229 30271 10287 30277
rect 11146 30268 11152 30320
rect 11204 30308 11210 30320
rect 11204 30280 12388 30308
rect 11204 30268 11210 30280
rect 12360 30252 12388 30280
rect 13354 30268 13360 30320
rect 13412 30268 13418 30320
rect 13906 30268 13912 30320
rect 13964 30308 13970 30320
rect 14550 30308 14556 30320
rect 13964 30280 14556 30308
rect 13964 30268 13970 30280
rect 14550 30268 14556 30280
rect 14608 30308 14614 30320
rect 15565 30311 15623 30317
rect 15565 30308 15577 30311
rect 14608 30280 15577 30308
rect 14608 30268 14614 30280
rect 15565 30277 15577 30280
rect 15611 30277 15623 30311
rect 16485 30311 16543 30317
rect 15565 30271 15623 30277
rect 15764 30280 16160 30308
rect 9585 30243 9643 30249
rect 9585 30209 9597 30243
rect 9631 30209 9643 30243
rect 9585 30203 9643 30209
rect 9769 30243 9827 30249
rect 9769 30209 9781 30243
rect 9815 30240 9827 30243
rect 10410 30240 10416 30252
rect 9815 30212 10416 30240
rect 9815 30209 9827 30212
rect 9769 30203 9827 30209
rect 10410 30200 10416 30212
rect 10468 30200 10474 30252
rect 11057 30243 11115 30249
rect 11057 30209 11069 30243
rect 11103 30209 11115 30243
rect 11057 30203 11115 30209
rect 11241 30243 11299 30249
rect 11241 30209 11253 30243
rect 11287 30240 11299 30243
rect 11698 30240 11704 30252
rect 11287 30212 11704 30240
rect 11287 30209 11299 30212
rect 11241 30203 11299 30209
rect 10870 30132 10876 30184
rect 10928 30132 10934 30184
rect 11072 30172 11100 30203
rect 11698 30200 11704 30212
rect 11756 30200 11762 30252
rect 12342 30200 12348 30252
rect 12400 30200 12406 30252
rect 14090 30200 14096 30252
rect 14148 30240 14154 30252
rect 15764 30249 15792 30280
rect 14369 30243 14427 30249
rect 14369 30240 14381 30243
rect 14148 30212 14381 30240
rect 14148 30200 14154 30212
rect 14369 30209 14381 30212
rect 14415 30209 14427 30243
rect 15749 30243 15807 30249
rect 15749 30240 15761 30243
rect 14369 30203 14427 30209
rect 14568 30212 15761 30240
rect 14568 30181 14596 30212
rect 15749 30209 15761 30212
rect 15795 30209 15807 30243
rect 15749 30203 15807 30209
rect 16022 30200 16028 30252
rect 16080 30200 16086 30252
rect 12621 30175 12679 30181
rect 11072 30144 12434 30172
rect 842 30064 848 30116
rect 900 30104 906 30116
rect 1397 30107 1455 30113
rect 1397 30104 1409 30107
rect 900 30076 1409 30104
rect 900 30064 906 30076
rect 1397 30073 1409 30076
rect 1443 30073 1455 30107
rect 1397 30067 1455 30073
rect 3878 30064 3884 30116
rect 3936 30104 3942 30116
rect 7098 30104 7104 30116
rect 3936 30076 7104 30104
rect 3936 30064 3942 30076
rect 7098 30064 7104 30076
rect 7156 30064 7162 30116
rect 11057 30107 11115 30113
rect 11057 30073 11069 30107
rect 11103 30104 11115 30107
rect 11238 30104 11244 30116
rect 11103 30076 11244 30104
rect 11103 30073 11115 30076
rect 11057 30067 11115 30073
rect 11238 30064 11244 30076
rect 11296 30064 11302 30116
rect 9214 29996 9220 30048
rect 9272 30036 9278 30048
rect 9677 30039 9735 30045
rect 9677 30036 9689 30039
rect 9272 30008 9689 30036
rect 9272 29996 9278 30008
rect 9677 30005 9689 30008
rect 9723 30005 9735 30039
rect 12406 30036 12434 30144
rect 12621 30141 12633 30175
rect 12667 30172 12679 30175
rect 14185 30175 14243 30181
rect 14185 30172 14197 30175
rect 12667 30144 14197 30172
rect 12667 30141 12679 30144
rect 12621 30135 12679 30141
rect 14185 30141 14197 30144
rect 14231 30141 14243 30175
rect 14185 30135 14243 30141
rect 14553 30175 14611 30181
rect 14553 30141 14565 30175
rect 14599 30141 14611 30175
rect 14553 30135 14611 30141
rect 14642 30132 14648 30184
rect 14700 30132 14706 30184
rect 14826 30132 14832 30184
rect 14884 30172 14890 30184
rect 15286 30172 15292 30184
rect 14884 30144 15292 30172
rect 14884 30132 14890 30144
rect 15286 30132 15292 30144
rect 15344 30172 15350 30184
rect 15381 30175 15439 30181
rect 15381 30172 15393 30175
rect 15344 30144 15393 30172
rect 15344 30132 15350 30144
rect 15381 30141 15393 30144
rect 15427 30141 15439 30175
rect 15381 30135 15439 30141
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30141 15991 30175
rect 16132 30172 16160 30280
rect 16485 30277 16497 30311
rect 16531 30308 16543 30311
rect 17037 30311 17095 30317
rect 17037 30308 17049 30311
rect 16531 30280 17049 30308
rect 16531 30277 16543 30280
rect 16485 30271 16543 30277
rect 17037 30277 17049 30280
rect 17083 30277 17095 30311
rect 17037 30271 17095 30277
rect 16301 30243 16359 30249
rect 16301 30209 16313 30243
rect 16347 30240 16359 30243
rect 17328 30240 17356 30339
rect 17402 30336 17408 30348
rect 17460 30336 17466 30388
rect 17862 30336 17868 30388
rect 17920 30376 17926 30388
rect 20717 30379 20775 30385
rect 17920 30348 19656 30376
rect 17920 30336 17926 30348
rect 18432 30308 18460 30348
rect 18354 30280 18460 30308
rect 16347 30212 17356 30240
rect 19061 30243 19119 30249
rect 16347 30209 16359 30212
rect 16301 30203 16359 30209
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 19334 30240 19340 30252
rect 19107 30212 19340 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 19334 30200 19340 30212
rect 19392 30200 19398 30252
rect 19426 30200 19432 30252
rect 19484 30200 19490 30252
rect 19628 30249 19656 30348
rect 20717 30345 20729 30379
rect 20763 30345 20775 30379
rect 20717 30339 20775 30345
rect 21269 30379 21327 30385
rect 21269 30345 21281 30379
rect 21315 30376 21327 30379
rect 21358 30376 21364 30388
rect 21315 30348 21364 30376
rect 21315 30345 21327 30348
rect 21269 30339 21327 30345
rect 20732 30308 20760 30339
rect 21358 30336 21364 30348
rect 21416 30336 21422 30388
rect 31846 30376 31852 30388
rect 30024 30348 31852 30376
rect 20272 30280 21680 30308
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30240 19671 30243
rect 19978 30240 19984 30252
rect 19659 30212 19984 30240
rect 19659 30209 19671 30212
rect 19613 30203 19671 30209
rect 19978 30200 19984 30212
rect 20036 30200 20042 30252
rect 20272 30249 20300 30280
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30209 20315 30243
rect 20257 30203 20315 30209
rect 20346 30200 20352 30252
rect 20404 30200 20410 30252
rect 20901 30243 20959 30249
rect 20901 30209 20913 30243
rect 20947 30240 20959 30243
rect 21082 30240 21088 30252
rect 20947 30212 21088 30240
rect 20947 30209 20959 30212
rect 20901 30203 20959 30209
rect 21082 30200 21088 30212
rect 21140 30200 21146 30252
rect 21453 30243 21511 30249
rect 21453 30209 21465 30243
rect 21499 30209 21511 30243
rect 21453 30203 21511 30209
rect 16666 30172 16672 30184
rect 16132 30144 16672 30172
rect 15933 30135 15991 30141
rect 14093 30107 14151 30113
rect 14093 30073 14105 30107
rect 14139 30104 14151 30107
rect 15010 30104 15016 30116
rect 14139 30076 15016 30104
rect 14139 30073 14151 30076
rect 14093 30067 14151 30073
rect 15010 30064 15016 30076
rect 15068 30104 15074 30116
rect 15948 30104 15976 30135
rect 16666 30132 16672 30144
rect 16724 30132 16730 30184
rect 18785 30175 18843 30181
rect 18785 30172 18797 30175
rect 17236 30144 18797 30172
rect 17236 30113 17264 30144
rect 18785 30141 18797 30144
rect 18831 30141 18843 30175
rect 18785 30135 18843 30141
rect 15068 30076 15976 30104
rect 17221 30107 17279 30113
rect 15068 30064 15074 30076
rect 17221 30073 17233 30107
rect 17267 30073 17279 30107
rect 21468 30104 21496 30203
rect 21652 30184 21680 30280
rect 22094 30268 22100 30320
rect 22152 30268 22158 30320
rect 23293 30311 23351 30317
rect 23293 30277 23305 30311
rect 23339 30308 23351 30311
rect 24397 30311 24455 30317
rect 24397 30308 24409 30311
rect 23339 30280 24409 30308
rect 23339 30277 23351 30280
rect 23293 30271 23351 30277
rect 24397 30277 24409 30280
rect 24443 30277 24455 30311
rect 26234 30308 26240 30320
rect 25622 30280 26240 30308
rect 24397 30271 24455 30277
rect 26234 30268 26240 30280
rect 26292 30268 26298 30320
rect 29270 30268 29276 30320
rect 29328 30308 29334 30320
rect 30024 30308 30052 30348
rect 30282 30308 30288 30320
rect 29328 30280 30052 30308
rect 30116 30280 30288 30308
rect 29328 30268 29334 30280
rect 21726 30200 21732 30252
rect 21784 30240 21790 30252
rect 21821 30243 21879 30249
rect 21821 30240 21833 30243
rect 21784 30212 21833 30240
rect 21784 30200 21790 30212
rect 21821 30209 21833 30212
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 21910 30200 21916 30252
rect 21968 30240 21974 30252
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21968 30212 22017 30240
rect 21968 30200 21974 30212
rect 22005 30209 22017 30212
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 21634 30132 21640 30184
rect 21692 30132 21698 30184
rect 22094 30132 22100 30184
rect 22152 30172 22158 30184
rect 22204 30172 22232 30203
rect 23474 30200 23480 30252
rect 23532 30200 23538 30252
rect 23842 30200 23848 30252
rect 23900 30200 23906 30252
rect 24026 30200 24032 30252
rect 24084 30200 24090 30252
rect 24118 30200 24124 30252
rect 24176 30200 24182 30252
rect 29638 30200 29644 30252
rect 29696 30200 29702 30252
rect 30116 30249 30144 30280
rect 30282 30268 30288 30280
rect 30340 30268 30346 30320
rect 30377 30311 30435 30317
rect 30377 30277 30389 30311
rect 30423 30308 30435 30311
rect 30466 30308 30472 30320
rect 30423 30280 30472 30308
rect 30423 30277 30435 30280
rect 30377 30271 30435 30277
rect 30466 30268 30472 30280
rect 30524 30268 30530 30320
rect 30576 30308 30604 30348
rect 31846 30336 31852 30348
rect 31904 30336 31910 30388
rect 34238 30336 34244 30388
rect 34296 30376 34302 30388
rect 34296 30348 34652 30376
rect 34296 30336 34302 30348
rect 30834 30308 30840 30320
rect 30576 30280 30840 30308
rect 30834 30268 30840 30280
rect 30892 30268 30898 30320
rect 33318 30308 33324 30320
rect 32784 30280 33324 30308
rect 30101 30243 30159 30249
rect 30101 30209 30113 30243
rect 30147 30209 30159 30243
rect 30101 30203 30159 30209
rect 32122 30200 32128 30252
rect 32180 30240 32186 30252
rect 32493 30243 32551 30249
rect 32493 30240 32505 30243
rect 32180 30212 32505 30240
rect 32180 30200 32186 30212
rect 32493 30209 32505 30212
rect 32539 30209 32551 30243
rect 32493 30203 32551 30209
rect 32582 30200 32588 30252
rect 32640 30240 32646 30252
rect 32784 30249 32812 30280
rect 33318 30268 33324 30280
rect 33376 30268 33382 30320
rect 34514 30268 34520 30320
rect 34572 30268 34578 30320
rect 34624 30308 34652 30348
rect 35066 30336 35072 30388
rect 35124 30376 35130 30388
rect 35437 30379 35495 30385
rect 35437 30376 35449 30379
rect 35124 30348 35449 30376
rect 35124 30336 35130 30348
rect 35437 30345 35449 30348
rect 35483 30345 35495 30379
rect 35437 30339 35495 30345
rect 34624 30280 35848 30308
rect 32677 30243 32735 30249
rect 32677 30240 32689 30243
rect 32640 30212 32689 30240
rect 32640 30200 32646 30212
rect 32677 30209 32689 30212
rect 32723 30209 32735 30243
rect 32677 30203 32735 30209
rect 32769 30243 32827 30249
rect 32769 30209 32781 30243
rect 32815 30209 32827 30243
rect 32769 30203 32827 30209
rect 32950 30200 32956 30252
rect 33008 30200 33014 30252
rect 33870 30200 33876 30252
rect 33928 30240 33934 30252
rect 34241 30243 34299 30249
rect 34241 30240 34253 30243
rect 33928 30212 34253 30240
rect 33928 30200 33934 30212
rect 34241 30209 34253 30212
rect 34287 30209 34299 30243
rect 34241 30203 34299 30209
rect 34333 30243 34391 30249
rect 34333 30209 34345 30243
rect 34379 30240 34391 30243
rect 34698 30240 34704 30252
rect 34379 30212 34704 30240
rect 34379 30209 34391 30212
rect 34333 30203 34391 30209
rect 34698 30200 34704 30212
rect 34756 30200 34762 30252
rect 35253 30243 35311 30249
rect 35253 30209 35265 30243
rect 35299 30240 35311 30243
rect 35342 30240 35348 30252
rect 35299 30212 35348 30240
rect 35299 30209 35311 30212
rect 35253 30203 35311 30209
rect 35342 30200 35348 30212
rect 35400 30200 35406 30252
rect 35434 30200 35440 30252
rect 35492 30240 35498 30252
rect 35820 30249 35848 30280
rect 35713 30243 35771 30249
rect 35713 30240 35725 30243
rect 35492 30212 35725 30240
rect 35492 30200 35498 30212
rect 35713 30209 35725 30212
rect 35759 30209 35771 30243
rect 35713 30203 35771 30209
rect 35805 30243 35863 30249
rect 35805 30209 35817 30243
rect 35851 30240 35863 30243
rect 36630 30240 36636 30252
rect 35851 30212 36636 30240
rect 35851 30209 35863 30212
rect 35805 30203 35863 30209
rect 36630 30200 36636 30212
rect 36688 30200 36694 30252
rect 22152 30144 22232 30172
rect 22152 30132 22158 30144
rect 23658 30132 23664 30184
rect 23716 30132 23722 30184
rect 23753 30175 23811 30181
rect 23753 30141 23765 30175
rect 23799 30172 23811 30175
rect 24854 30172 24860 30184
rect 23799 30144 24860 30172
rect 23799 30141 23811 30144
rect 23753 30135 23811 30141
rect 24854 30132 24860 30144
rect 24912 30132 24918 30184
rect 26050 30132 26056 30184
rect 26108 30172 26114 30184
rect 26513 30175 26571 30181
rect 26513 30172 26525 30175
rect 26108 30144 26525 30172
rect 26108 30132 26114 30144
rect 26513 30141 26525 30144
rect 26559 30141 26571 30175
rect 26513 30135 26571 30141
rect 26970 30132 26976 30184
rect 27028 30132 27034 30184
rect 34422 30132 34428 30184
rect 34480 30172 34486 30184
rect 35621 30175 35679 30181
rect 35621 30172 35633 30175
rect 34480 30144 35633 30172
rect 34480 30132 34486 30144
rect 35621 30141 35633 30144
rect 35667 30141 35679 30175
rect 35621 30135 35679 30141
rect 35897 30175 35955 30181
rect 35897 30141 35909 30175
rect 35943 30172 35955 30175
rect 35986 30172 35992 30184
rect 35943 30144 35992 30172
rect 35943 30141 35955 30144
rect 35897 30135 35955 30141
rect 35986 30132 35992 30144
rect 36044 30172 36050 30184
rect 37182 30172 37188 30184
rect 36044 30144 37188 30172
rect 36044 30132 36050 30144
rect 37182 30132 37188 30144
rect 37240 30132 37246 30184
rect 22373 30107 22431 30113
rect 22373 30104 22385 30107
rect 21468 30076 22385 30104
rect 17221 30067 17279 30073
rect 22373 30073 22385 30076
rect 22419 30073 22431 30107
rect 22373 30067 22431 30073
rect 22554 30064 22560 30116
rect 22612 30104 22618 30116
rect 24118 30104 24124 30116
rect 22612 30076 24124 30104
rect 22612 30064 22618 30076
rect 24118 30064 24124 30076
rect 24176 30064 24182 30116
rect 31849 30107 31907 30113
rect 31849 30073 31861 30107
rect 31895 30104 31907 30107
rect 32306 30104 32312 30116
rect 31895 30076 32312 30104
rect 31895 30073 31907 30076
rect 31849 30067 31907 30073
rect 32306 30064 32312 30076
rect 32364 30104 32370 30116
rect 32585 30107 32643 30113
rect 32585 30104 32597 30107
rect 32364 30076 32597 30104
rect 32364 30064 32370 30076
rect 32585 30073 32597 30076
rect 32631 30073 32643 30107
rect 32585 30067 32643 30073
rect 34517 30107 34575 30113
rect 34517 30073 34529 30107
rect 34563 30104 34575 30107
rect 34606 30104 34612 30116
rect 34563 30076 34612 30104
rect 34563 30073 34575 30076
rect 34517 30067 34575 30073
rect 34606 30064 34612 30076
rect 34664 30064 34670 30116
rect 12618 30036 12624 30048
rect 12406 30008 12624 30036
rect 9677 29999 9735 30005
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 17034 29996 17040 30048
rect 17092 29996 17098 30048
rect 19150 29996 19156 30048
rect 19208 30036 19214 30048
rect 19245 30039 19303 30045
rect 19245 30036 19257 30039
rect 19208 30008 19257 30036
rect 19208 29996 19214 30008
rect 19245 30005 19257 30008
rect 19291 30005 19303 30039
rect 19245 29999 19303 30005
rect 20530 29996 20536 30048
rect 20588 29996 20594 30048
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 24578 30036 24584 30048
rect 20864 30008 24584 30036
rect 20864 29996 20870 30008
rect 24578 29996 24584 30008
rect 24636 29996 24642 30048
rect 24946 29996 24952 30048
rect 25004 30036 25010 30048
rect 25406 30036 25412 30048
rect 25004 30008 25412 30036
rect 25004 29996 25010 30008
rect 25406 29996 25412 30008
rect 25464 30036 25470 30048
rect 25869 30039 25927 30045
rect 25869 30036 25881 30039
rect 25464 30008 25881 30036
rect 25464 29996 25470 30008
rect 25869 30005 25881 30008
rect 25915 30005 25927 30039
rect 25869 29999 25927 30005
rect 25958 29996 25964 30048
rect 26016 29996 26022 30048
rect 27522 29996 27528 30048
rect 27580 30036 27586 30048
rect 27617 30039 27675 30045
rect 27617 30036 27629 30039
rect 27580 30008 27629 30036
rect 27580 29996 27586 30008
rect 27617 30005 27629 30008
rect 27663 30005 27675 30039
rect 27617 29999 27675 30005
rect 29914 29996 29920 30048
rect 29972 29996 29978 30048
rect 32217 30039 32275 30045
rect 32217 30005 32229 30039
rect 32263 30036 32275 30039
rect 37458 30036 37464 30048
rect 32263 30008 37464 30036
rect 32263 30005 32275 30008
rect 32217 29999 32275 30005
rect 37458 29996 37464 30008
rect 37516 29996 37522 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 12713 29835 12771 29841
rect 12713 29801 12725 29835
rect 12759 29832 12771 29835
rect 13354 29832 13360 29844
rect 12759 29804 13360 29832
rect 12759 29801 12771 29804
rect 12713 29795 12771 29801
rect 13354 29792 13360 29804
rect 13412 29792 13418 29844
rect 14369 29835 14427 29841
rect 14369 29801 14381 29835
rect 14415 29832 14427 29835
rect 14642 29832 14648 29844
rect 14415 29804 14648 29832
rect 14415 29801 14427 29804
rect 14369 29795 14427 29801
rect 14642 29792 14648 29804
rect 14700 29792 14706 29844
rect 17218 29792 17224 29844
rect 17276 29792 17282 29844
rect 17310 29792 17316 29844
rect 17368 29792 17374 29844
rect 17402 29792 17408 29844
rect 17460 29832 17466 29844
rect 17497 29835 17555 29841
rect 17497 29832 17509 29835
rect 17460 29804 17509 29832
rect 17460 29792 17466 29804
rect 17497 29801 17509 29804
rect 17543 29801 17555 29835
rect 17497 29795 17555 29801
rect 19337 29835 19395 29841
rect 19337 29801 19349 29835
rect 19383 29832 19395 29835
rect 19426 29832 19432 29844
rect 19383 29804 19432 29832
rect 19383 29801 19395 29804
rect 19337 29795 19395 29801
rect 19426 29792 19432 29804
rect 19484 29792 19490 29844
rect 22738 29832 22744 29844
rect 19720 29804 22744 29832
rect 11241 29767 11299 29773
rect 11241 29733 11253 29767
rect 11287 29764 11299 29767
rect 11517 29767 11575 29773
rect 11517 29764 11529 29767
rect 11287 29736 11529 29764
rect 11287 29733 11299 29736
rect 11241 29727 11299 29733
rect 11517 29733 11529 29736
rect 11563 29733 11575 29767
rect 11517 29727 11575 29733
rect 18322 29724 18328 29776
rect 18380 29764 18386 29776
rect 18877 29767 18935 29773
rect 18877 29764 18889 29767
rect 18380 29736 18889 29764
rect 18380 29724 18386 29736
rect 18877 29733 18889 29736
rect 18923 29764 18935 29767
rect 19720 29764 19748 29804
rect 22738 29792 22744 29804
rect 22796 29792 22802 29844
rect 24026 29792 24032 29844
rect 24084 29832 24090 29844
rect 24121 29835 24179 29841
rect 24121 29832 24133 29835
rect 24084 29804 24133 29832
rect 24084 29792 24090 29804
rect 24121 29801 24133 29804
rect 24167 29801 24179 29835
rect 24121 29795 24179 29801
rect 25961 29835 26019 29841
rect 25961 29801 25973 29835
rect 26007 29832 26019 29835
rect 26970 29832 26976 29844
rect 26007 29804 26976 29832
rect 26007 29801 26019 29804
rect 25961 29795 26019 29801
rect 26970 29792 26976 29804
rect 27028 29792 27034 29844
rect 28902 29792 28908 29844
rect 28960 29832 28966 29844
rect 30469 29835 30527 29841
rect 30469 29832 30481 29835
rect 28960 29804 30481 29832
rect 28960 29792 28966 29804
rect 30469 29801 30481 29804
rect 30515 29832 30527 29835
rect 30558 29832 30564 29844
rect 30515 29804 30564 29832
rect 30515 29801 30527 29804
rect 30469 29795 30527 29801
rect 30558 29792 30564 29804
rect 30616 29792 30622 29844
rect 31113 29835 31171 29841
rect 31113 29801 31125 29835
rect 31159 29801 31171 29835
rect 31113 29795 31171 29801
rect 32769 29835 32827 29841
rect 32769 29801 32781 29835
rect 32815 29832 32827 29835
rect 32950 29832 32956 29844
rect 32815 29804 32956 29832
rect 32815 29801 32827 29804
rect 32769 29795 32827 29801
rect 18923 29736 19748 29764
rect 18923 29733 18935 29736
rect 18877 29727 18935 29733
rect 23658 29724 23664 29776
rect 23716 29764 23722 29776
rect 24762 29764 24768 29776
rect 23716 29736 24768 29764
rect 23716 29724 23722 29736
rect 24762 29724 24768 29736
rect 24820 29724 24826 29776
rect 26050 29724 26056 29776
rect 26108 29724 26114 29776
rect 28534 29724 28540 29776
rect 28592 29724 28598 29776
rect 30282 29764 30288 29776
rect 28828 29736 30288 29764
rect 4525 29699 4583 29705
rect 4525 29665 4537 29699
rect 4571 29696 4583 29699
rect 4706 29696 4712 29708
rect 4571 29668 4712 29696
rect 4571 29665 4583 29668
rect 4525 29659 4583 29665
rect 4706 29656 4712 29668
rect 4764 29656 4770 29708
rect 4985 29699 5043 29705
rect 4985 29665 4997 29699
rect 5031 29696 5043 29699
rect 5258 29696 5264 29708
rect 5031 29668 5264 29696
rect 5031 29665 5043 29668
rect 4985 29659 5043 29665
rect 5258 29656 5264 29668
rect 5316 29656 5322 29708
rect 7929 29699 7987 29705
rect 7929 29696 7941 29699
rect 6380 29668 7941 29696
rect 842 29588 848 29640
rect 900 29628 906 29640
rect 1397 29631 1455 29637
rect 1397 29628 1409 29631
rect 900 29600 1409 29628
rect 900 29588 906 29600
rect 1397 29597 1409 29600
rect 1443 29597 1455 29631
rect 1397 29591 1455 29597
rect 3326 29588 3332 29640
rect 3384 29628 3390 29640
rect 3789 29631 3847 29637
rect 3789 29628 3801 29631
rect 3384 29600 3801 29628
rect 3384 29588 3390 29600
rect 3789 29597 3801 29600
rect 3835 29597 3847 29631
rect 3789 29591 3847 29597
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29628 4951 29631
rect 5353 29631 5411 29637
rect 5353 29628 5365 29631
rect 4939 29600 5365 29628
rect 4939 29597 4951 29600
rect 4893 29591 4951 29597
rect 5353 29597 5365 29600
rect 5399 29597 5411 29631
rect 5353 29591 5411 29597
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29628 6055 29631
rect 6178 29628 6184 29640
rect 6043 29600 6184 29628
rect 6043 29597 6055 29600
rect 5997 29591 6055 29597
rect 6178 29588 6184 29600
rect 6236 29588 6242 29640
rect 6380 29572 6408 29668
rect 7929 29665 7941 29668
rect 7975 29665 7987 29699
rect 7929 29659 7987 29665
rect 9214 29656 9220 29708
rect 9272 29656 9278 29708
rect 10410 29656 10416 29708
rect 10468 29696 10474 29708
rect 11333 29699 11391 29705
rect 11333 29696 11345 29699
rect 10468 29668 11345 29696
rect 10468 29656 10474 29668
rect 11333 29665 11345 29668
rect 11379 29665 11391 29699
rect 11333 29659 11391 29665
rect 15010 29656 15016 29708
rect 15068 29656 15074 29708
rect 15746 29656 15752 29708
rect 15804 29656 15810 29708
rect 23842 29656 23848 29708
rect 23900 29696 23906 29708
rect 24578 29696 24584 29708
rect 23900 29668 24584 29696
rect 23900 29656 23906 29668
rect 24578 29656 24584 29668
rect 24636 29696 24642 29708
rect 25501 29699 25559 29705
rect 24636 29668 25452 29696
rect 24636 29656 24642 29668
rect 7466 29588 7472 29640
rect 7524 29628 7530 29640
rect 7561 29631 7619 29637
rect 7561 29628 7573 29631
rect 7524 29600 7573 29628
rect 7524 29588 7530 29600
rect 7561 29597 7573 29600
rect 7607 29597 7619 29631
rect 7561 29591 7619 29597
rect 7650 29588 7656 29640
rect 7708 29628 7714 29640
rect 7837 29631 7895 29637
rect 7837 29628 7849 29631
rect 7708 29600 7849 29628
rect 7708 29588 7714 29600
rect 7837 29597 7849 29600
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 8110 29588 8116 29640
rect 8168 29628 8174 29640
rect 8665 29631 8723 29637
rect 8665 29628 8677 29631
rect 8168 29600 8677 29628
rect 8168 29588 8174 29600
rect 8665 29597 8677 29600
rect 8711 29597 8723 29631
rect 8665 29591 8723 29597
rect 8938 29588 8944 29640
rect 8996 29588 9002 29640
rect 10965 29631 11023 29637
rect 10965 29597 10977 29631
rect 11011 29628 11023 29631
rect 11146 29628 11152 29640
rect 11011 29600 11152 29628
rect 11011 29597 11023 29600
rect 10965 29591 11023 29597
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 11609 29631 11667 29637
rect 11609 29597 11621 29631
rect 11655 29628 11667 29631
rect 12618 29628 12624 29640
rect 11655 29600 12624 29628
rect 11655 29597 11667 29600
rect 11609 29591 11667 29597
rect 12618 29588 12624 29600
rect 12676 29588 12682 29640
rect 15194 29588 15200 29640
rect 15252 29628 15258 29640
rect 15473 29631 15531 29637
rect 15473 29628 15485 29631
rect 15252 29600 15485 29628
rect 15252 29588 15258 29600
rect 15473 29597 15485 29600
rect 15519 29597 15531 29631
rect 15473 29591 15531 29597
rect 17218 29588 17224 29640
rect 17276 29628 17282 29640
rect 17276 29600 17724 29628
rect 17276 29588 17282 29600
rect 3513 29563 3571 29569
rect 3513 29529 3525 29563
rect 3559 29560 3571 29563
rect 3878 29560 3884 29572
rect 3559 29532 3884 29560
rect 3559 29529 3571 29532
rect 3513 29523 3571 29529
rect 3878 29520 3884 29532
rect 3936 29520 3942 29572
rect 6362 29520 6368 29572
rect 6420 29520 6426 29572
rect 6822 29520 6828 29572
rect 6880 29560 6886 29572
rect 7193 29563 7251 29569
rect 7193 29560 7205 29563
rect 6880 29532 7205 29560
rect 6880 29520 6886 29532
rect 7193 29529 7205 29532
rect 7239 29560 7251 29563
rect 8956 29560 8984 29588
rect 7239 29532 8984 29560
rect 7239 29529 7251 29532
rect 7193 29523 7251 29529
rect 10226 29520 10232 29572
rect 10284 29520 10290 29572
rect 11241 29563 11299 29569
rect 11241 29529 11253 29563
rect 11287 29560 11299 29563
rect 11514 29560 11520 29572
rect 11287 29532 11520 29560
rect 11287 29529 11299 29532
rect 11241 29523 11299 29529
rect 11514 29520 11520 29532
rect 11572 29520 11578 29572
rect 17494 29569 17500 29572
rect 12437 29563 12495 29569
rect 12437 29529 12449 29563
rect 12483 29529 12495 29563
rect 17481 29563 17500 29569
rect 16974 29532 17448 29560
rect 12437 29523 12495 29529
rect 3418 29452 3424 29504
rect 3476 29452 3482 29504
rect 4246 29452 4252 29504
rect 4304 29492 4310 29504
rect 4433 29495 4491 29501
rect 4433 29492 4445 29495
rect 4304 29464 4445 29492
rect 4304 29452 4310 29464
rect 4433 29461 4445 29464
rect 4479 29461 4491 29495
rect 4433 29455 4491 29461
rect 7374 29452 7380 29504
rect 7432 29452 7438 29504
rect 7745 29495 7803 29501
rect 7745 29461 7757 29495
rect 7791 29492 7803 29495
rect 8113 29495 8171 29501
rect 8113 29492 8125 29495
rect 7791 29464 8125 29492
rect 7791 29461 7803 29464
rect 7745 29455 7803 29461
rect 8113 29461 8125 29464
rect 8159 29461 8171 29495
rect 8113 29455 8171 29461
rect 9398 29452 9404 29504
rect 9456 29492 9462 29504
rect 10689 29495 10747 29501
rect 10689 29492 10701 29495
rect 9456 29464 10701 29492
rect 9456 29452 9462 29464
rect 10689 29461 10701 29464
rect 10735 29492 10747 29495
rect 10870 29492 10876 29504
rect 10735 29464 10876 29492
rect 10735 29461 10747 29464
rect 10689 29455 10747 29461
rect 10870 29452 10876 29464
rect 10928 29492 10934 29504
rect 11057 29495 11115 29501
rect 11057 29492 11069 29495
rect 10928 29464 11069 29492
rect 10928 29452 10934 29464
rect 11057 29461 11069 29464
rect 11103 29461 11115 29495
rect 11057 29455 11115 29461
rect 11333 29495 11391 29501
rect 11333 29461 11345 29495
rect 11379 29492 11391 29495
rect 11422 29492 11428 29504
rect 11379 29464 11428 29492
rect 11379 29461 11391 29464
rect 11333 29455 11391 29461
rect 11422 29452 11428 29464
rect 11480 29452 11486 29504
rect 12452 29492 12480 29523
rect 12989 29495 13047 29501
rect 12989 29492 13001 29495
rect 12452 29464 13001 29492
rect 12989 29461 13001 29464
rect 13035 29492 13047 29495
rect 15102 29492 15108 29504
rect 13035 29464 15108 29492
rect 13035 29461 13047 29464
rect 12989 29455 13047 29461
rect 15102 29452 15108 29464
rect 15160 29452 15166 29504
rect 17420 29492 17448 29532
rect 17481 29529 17493 29563
rect 17481 29523 17500 29529
rect 17494 29520 17500 29523
rect 17552 29520 17558 29572
rect 17696 29569 17724 29600
rect 18782 29588 18788 29640
rect 18840 29628 18846 29640
rect 19242 29628 19248 29640
rect 18840 29600 19248 29628
rect 18840 29588 18846 29600
rect 19242 29588 19248 29600
rect 19300 29628 19306 29640
rect 19521 29631 19579 29637
rect 19521 29628 19533 29631
rect 19300 29600 19533 29628
rect 19300 29588 19306 29600
rect 19521 29597 19533 29600
rect 19567 29597 19579 29631
rect 19521 29591 19579 29597
rect 19613 29631 19671 29637
rect 19613 29597 19625 29631
rect 19659 29628 19671 29631
rect 19659 29600 19840 29628
rect 19659 29597 19671 29600
rect 19613 29591 19671 29597
rect 17681 29563 17739 29569
rect 17681 29529 17693 29563
rect 17727 29529 17739 29563
rect 17681 29523 17739 29529
rect 19702 29520 19708 29572
rect 19760 29520 19766 29572
rect 19812 29560 19840 29600
rect 19886 29588 19892 29640
rect 19944 29588 19950 29640
rect 20530 29588 20536 29640
rect 20588 29628 20594 29640
rect 21094 29631 21152 29637
rect 21094 29628 21106 29631
rect 20588 29600 21106 29628
rect 20588 29588 20594 29600
rect 21094 29597 21106 29600
rect 21140 29597 21152 29631
rect 21094 29591 21152 29597
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29628 21419 29631
rect 21729 29631 21787 29637
rect 21729 29628 21741 29631
rect 21407 29600 21741 29628
rect 21407 29597 21419 29600
rect 21361 29591 21419 29597
rect 21729 29597 21741 29600
rect 21775 29628 21787 29631
rect 22554 29628 22560 29640
rect 21775 29600 22560 29628
rect 21775 29597 21787 29600
rect 21729 29591 21787 29597
rect 22554 29588 22560 29600
rect 22612 29588 22618 29640
rect 23477 29631 23535 29637
rect 23477 29628 23489 29631
rect 22756 29600 23489 29628
rect 20254 29560 20260 29572
rect 19812 29532 20260 29560
rect 20254 29520 20260 29532
rect 20312 29560 20318 29572
rect 21996 29563 22054 29569
rect 20312 29532 20944 29560
rect 20312 29520 20318 29532
rect 17862 29492 17868 29504
rect 17420 29464 17868 29492
rect 17862 29452 17868 29464
rect 17920 29452 17926 29504
rect 19981 29495 20039 29501
rect 19981 29461 19993 29495
rect 20027 29492 20039 29495
rect 20806 29492 20812 29504
rect 20027 29464 20812 29492
rect 20027 29461 20039 29464
rect 19981 29455 20039 29461
rect 20806 29452 20812 29464
rect 20864 29452 20870 29504
rect 20916 29492 20944 29532
rect 21996 29529 22008 29563
rect 22042 29560 22054 29563
rect 22462 29560 22468 29572
rect 22042 29532 22468 29560
rect 22042 29529 22054 29532
rect 21996 29523 22054 29529
rect 22462 29520 22468 29532
rect 22520 29520 22526 29572
rect 22756 29492 22784 29600
rect 23477 29597 23489 29600
rect 23523 29597 23535 29631
rect 23937 29631 23995 29637
rect 23937 29628 23949 29631
rect 23477 29591 23535 29597
rect 23584 29600 23949 29628
rect 23290 29520 23296 29572
rect 23348 29520 23354 29572
rect 23584 29560 23612 29600
rect 23937 29597 23949 29600
rect 23983 29597 23995 29631
rect 23937 29591 23995 29597
rect 24118 29588 24124 29640
rect 24176 29628 24182 29640
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 24176 29600 24409 29628
rect 24176 29588 24182 29600
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 25222 29588 25228 29640
rect 25280 29588 25286 29640
rect 25424 29637 25452 29668
rect 25501 29665 25513 29699
rect 25547 29696 25559 29699
rect 25958 29696 25964 29708
rect 25547 29668 25964 29696
rect 25547 29665 25559 29668
rect 25501 29659 25559 29665
rect 25958 29656 25964 29668
rect 26016 29656 26022 29708
rect 27522 29656 27528 29708
rect 27580 29656 27586 29708
rect 27801 29699 27859 29705
rect 27801 29665 27813 29699
rect 27847 29696 27859 29699
rect 28828 29696 28856 29736
rect 30282 29724 30288 29736
rect 30340 29724 30346 29776
rect 27847 29668 28856 29696
rect 27847 29665 27859 29668
rect 27801 29659 27859 29665
rect 28902 29656 28908 29708
rect 28960 29656 28966 29708
rect 29089 29699 29147 29705
rect 29089 29665 29101 29699
rect 29135 29696 29147 29699
rect 29730 29696 29736 29708
rect 29135 29668 29736 29696
rect 29135 29665 29147 29668
rect 29089 29659 29147 29665
rect 25409 29631 25467 29637
rect 25409 29597 25421 29631
rect 25455 29597 25467 29631
rect 25409 29591 25467 29597
rect 25593 29631 25651 29637
rect 25593 29597 25605 29631
rect 25639 29597 25651 29631
rect 25593 29591 25651 29597
rect 23400 29532 23612 29560
rect 23753 29563 23811 29569
rect 20916 29464 22784 29492
rect 23106 29452 23112 29504
rect 23164 29492 23170 29504
rect 23400 29492 23428 29532
rect 23753 29529 23765 29563
rect 23799 29560 23811 29563
rect 24026 29560 24032 29572
rect 23799 29532 24032 29560
rect 23799 29529 23811 29532
rect 23753 29523 23811 29529
rect 24026 29520 24032 29532
rect 24084 29560 24090 29572
rect 24486 29560 24492 29572
rect 24084 29532 24492 29560
rect 24084 29520 24090 29532
rect 24486 29520 24492 29532
rect 24544 29520 24550 29572
rect 24762 29520 24768 29572
rect 24820 29560 24826 29572
rect 25608 29560 25636 29591
rect 25774 29588 25780 29640
rect 25832 29588 25838 29640
rect 28813 29631 28871 29637
rect 28813 29597 28825 29631
rect 28859 29628 28871 29631
rect 29104 29628 29132 29659
rect 29730 29656 29736 29668
rect 29788 29656 29794 29708
rect 31128 29696 31156 29795
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 33502 29792 33508 29844
rect 33560 29832 33566 29844
rect 34330 29832 34336 29844
rect 33560 29804 34336 29832
rect 33560 29792 33566 29804
rect 34330 29792 34336 29804
rect 34388 29792 34394 29844
rect 35434 29832 35440 29844
rect 34440 29804 35440 29832
rect 34440 29696 34468 29804
rect 35434 29792 35440 29804
rect 35492 29792 35498 29844
rect 36725 29767 36783 29773
rect 36725 29733 36737 29767
rect 36771 29764 36783 29767
rect 37274 29764 37280 29776
rect 36771 29736 37280 29764
rect 36771 29733 36783 29736
rect 36725 29727 36783 29733
rect 37274 29724 37280 29736
rect 37332 29724 37338 29776
rect 30116 29668 31156 29696
rect 33060 29668 34468 29696
rect 34701 29699 34759 29705
rect 28859 29600 29132 29628
rect 29181 29631 29239 29637
rect 28859 29597 28871 29600
rect 28813 29591 28871 29597
rect 29181 29597 29193 29631
rect 29227 29628 29239 29631
rect 29822 29628 29828 29640
rect 29227 29600 29828 29628
rect 29227 29597 29239 29600
rect 29181 29591 29239 29597
rect 29822 29588 29828 29600
rect 29880 29628 29886 29640
rect 30116 29637 30144 29668
rect 33060 29640 33088 29668
rect 34701 29665 34713 29699
rect 34747 29696 34759 29699
rect 35342 29696 35348 29708
rect 34747 29668 35348 29696
rect 34747 29665 34759 29668
rect 34701 29659 34759 29665
rect 35342 29656 35348 29668
rect 35400 29656 35406 29708
rect 30101 29631 30159 29637
rect 30101 29628 30113 29631
rect 29880 29600 30113 29628
rect 29880 29588 29886 29600
rect 30101 29597 30113 29600
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 30837 29631 30895 29637
rect 30837 29597 30849 29631
rect 30883 29597 30895 29631
rect 30837 29591 30895 29597
rect 24820 29532 25636 29560
rect 24820 29520 24826 29532
rect 26234 29520 26240 29572
rect 26292 29560 26298 29572
rect 28537 29563 28595 29569
rect 26292 29532 26358 29560
rect 26292 29520 26298 29532
rect 28537 29529 28549 29563
rect 28583 29529 28595 29563
rect 28537 29523 28595 29529
rect 28721 29563 28779 29569
rect 28721 29529 28733 29563
rect 28767 29560 28779 29563
rect 29549 29563 29607 29569
rect 29549 29560 29561 29563
rect 28767 29532 29561 29560
rect 28767 29529 28779 29532
rect 28721 29523 28779 29529
rect 29549 29529 29561 29532
rect 29595 29529 29607 29563
rect 30852 29560 30880 29591
rect 32122 29588 32128 29640
rect 32180 29628 32186 29640
rect 32953 29631 33011 29637
rect 32953 29628 32965 29631
rect 32180 29600 32965 29628
rect 32180 29588 32186 29600
rect 32953 29597 32965 29600
rect 32999 29597 33011 29631
rect 32953 29591 33011 29597
rect 33042 29588 33048 29640
rect 33100 29588 33106 29640
rect 33226 29588 33232 29640
rect 33284 29588 33290 29640
rect 33321 29631 33379 29637
rect 33321 29597 33333 29631
rect 33367 29628 33379 29631
rect 33686 29628 33692 29640
rect 33367 29600 33692 29628
rect 33367 29597 33379 29600
rect 33321 29591 33379 29597
rect 33686 29588 33692 29600
rect 33744 29588 33750 29640
rect 33870 29588 33876 29640
rect 33928 29628 33934 29640
rect 33965 29631 34023 29637
rect 33965 29628 33977 29631
rect 33928 29600 33977 29628
rect 33928 29588 33934 29600
rect 33965 29597 33977 29600
rect 34011 29597 34023 29631
rect 33965 29591 34023 29597
rect 36078 29588 36084 29640
rect 36136 29588 36142 29640
rect 36722 29588 36728 29640
rect 36780 29588 36786 29640
rect 36814 29588 36820 29640
rect 36872 29628 36878 29640
rect 37001 29631 37059 29637
rect 37001 29628 37013 29631
rect 36872 29600 37013 29628
rect 36872 29588 36878 29600
rect 37001 29597 37013 29600
rect 37047 29597 37059 29631
rect 37001 29591 37059 29597
rect 31297 29563 31355 29569
rect 30852 29532 31248 29560
rect 29549 29523 29607 29529
rect 23164 29464 23428 29492
rect 23661 29495 23719 29501
rect 23164 29452 23170 29464
rect 23661 29461 23673 29495
rect 23707 29492 23719 29495
rect 24394 29492 24400 29504
rect 23707 29464 24400 29492
rect 23707 29461 23719 29464
rect 23661 29455 23719 29461
rect 24394 29452 24400 29464
rect 24452 29452 24458 29504
rect 24854 29452 24860 29504
rect 24912 29492 24918 29504
rect 25041 29495 25099 29501
rect 25041 29492 25053 29495
rect 24912 29464 25053 29492
rect 24912 29452 24918 29464
rect 25041 29461 25053 29464
rect 25087 29461 25099 29495
rect 28552 29492 28580 29523
rect 28905 29495 28963 29501
rect 28905 29492 28917 29495
rect 28552 29464 28917 29492
rect 25041 29455 25099 29461
rect 28905 29461 28917 29464
rect 28951 29461 28963 29495
rect 28905 29455 28963 29461
rect 30285 29495 30343 29501
rect 30285 29461 30297 29495
rect 30331 29492 30343 29495
rect 30374 29492 30380 29504
rect 30331 29464 30380 29492
rect 30331 29461 30343 29464
rect 30285 29455 30343 29461
rect 30374 29452 30380 29464
rect 30432 29452 30438 29504
rect 30466 29452 30472 29504
rect 30524 29452 30530 29504
rect 30944 29501 30972 29532
rect 31110 29501 31116 29504
rect 30929 29495 30987 29501
rect 30929 29461 30941 29495
rect 30975 29461 30987 29495
rect 30929 29455 30987 29461
rect 31097 29495 31116 29501
rect 31097 29461 31109 29495
rect 31097 29455 31116 29461
rect 31110 29452 31116 29455
rect 31168 29452 31174 29504
rect 31220 29492 31248 29532
rect 31297 29529 31309 29563
rect 31343 29560 31355 29563
rect 31846 29560 31852 29572
rect 31343 29532 31852 29560
rect 31343 29529 31355 29532
rect 31297 29523 31355 29529
rect 31846 29520 31852 29532
rect 31904 29520 31910 29572
rect 34977 29563 35035 29569
rect 34977 29529 34989 29563
rect 35023 29529 35035 29563
rect 34977 29523 35035 29529
rect 34146 29492 34152 29504
rect 31220 29464 34152 29492
rect 34146 29452 34152 29464
rect 34204 29452 34210 29504
rect 34330 29452 34336 29504
rect 34388 29452 34394 29504
rect 34517 29495 34575 29501
rect 34517 29461 34529 29495
rect 34563 29492 34575 29495
rect 34992 29492 35020 29523
rect 34563 29464 35020 29492
rect 34563 29461 34575 29464
rect 34517 29455 34575 29461
rect 36446 29452 36452 29504
rect 36504 29452 36510 29504
rect 36909 29495 36967 29501
rect 36909 29461 36921 29495
rect 36955 29492 36967 29495
rect 37182 29492 37188 29504
rect 36955 29464 37188 29492
rect 36955 29461 36967 29464
rect 36909 29455 36967 29461
rect 37182 29452 37188 29464
rect 37240 29452 37246 29504
rect 1104 29402 38824 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 38824 29402
rect 1104 29328 38824 29350
rect 3896 29260 5856 29288
rect 3418 29220 3424 29232
rect 3266 29192 3424 29220
rect 3418 29180 3424 29192
rect 3476 29220 3482 29232
rect 3896 29220 3924 29260
rect 4798 29220 4804 29232
rect 3476 29192 3924 29220
rect 3988 29192 4804 29220
rect 3476 29180 3482 29192
rect 3988 29161 4016 29192
rect 3973 29155 4031 29161
rect 3973 29121 3985 29155
rect 4019 29121 4031 29155
rect 3973 29115 4031 29121
rect 4062 29112 4068 29164
rect 4120 29112 4126 29164
rect 4246 29112 4252 29164
rect 4304 29112 4310 29164
rect 4448 29161 4476 29192
rect 4798 29180 4804 29192
rect 4856 29180 4862 29232
rect 5828 29164 5856 29260
rect 8018 29248 8024 29300
rect 8076 29288 8082 29300
rect 8941 29291 8999 29297
rect 8076 29260 8432 29288
rect 8076 29248 8082 29260
rect 7101 29223 7159 29229
rect 7101 29189 7113 29223
rect 7147 29220 7159 29223
rect 7374 29220 7380 29232
rect 7147 29192 7380 29220
rect 7147 29189 7159 29192
rect 7101 29183 7159 29189
rect 7374 29180 7380 29192
rect 7432 29180 7438 29232
rect 8404 29220 8432 29260
rect 8941 29257 8953 29291
rect 8987 29288 8999 29291
rect 10226 29288 10232 29300
rect 8987 29260 10232 29288
rect 8987 29257 8999 29260
rect 8941 29251 8999 29257
rect 8956 29220 8984 29251
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 11514 29248 11520 29300
rect 11572 29248 11578 29300
rect 12618 29248 12624 29300
rect 12676 29248 12682 29300
rect 14826 29248 14832 29300
rect 14884 29248 14890 29300
rect 19242 29248 19248 29300
rect 19300 29288 19306 29300
rect 19300 29260 20208 29288
rect 19300 29248 19306 29260
rect 8326 29192 8984 29220
rect 10870 29180 10876 29232
rect 10928 29220 10934 29232
rect 12253 29223 12311 29229
rect 12253 29220 12265 29223
rect 10928 29192 12265 29220
rect 10928 29180 10934 29192
rect 12253 29189 12265 29192
rect 12299 29189 12311 29223
rect 12453 29223 12511 29229
rect 12453 29220 12465 29223
rect 12253 29183 12311 29189
rect 12452 29189 12465 29220
rect 12499 29189 12511 29223
rect 12452 29183 12511 29189
rect 4433 29155 4491 29161
rect 4433 29121 4445 29155
rect 4479 29121 4491 29155
rect 4433 29115 4491 29121
rect 5810 29112 5816 29164
rect 5868 29112 5874 29164
rect 6822 29112 6828 29164
rect 6880 29112 6886 29164
rect 9033 29155 9091 29161
rect 9033 29121 9045 29155
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 842 29044 848 29096
rect 900 29084 906 29096
rect 1397 29087 1455 29093
rect 1397 29084 1409 29087
rect 900 29056 1409 29084
rect 900 29044 906 29056
rect 1397 29053 1409 29056
rect 1443 29053 1455 29087
rect 1397 29047 1455 29053
rect 2225 29087 2283 29093
rect 2225 29053 2237 29087
rect 2271 29084 2283 29087
rect 3326 29084 3332 29096
rect 2271 29056 3332 29084
rect 2271 29053 2283 29056
rect 2225 29047 2283 29053
rect 3326 29044 3332 29056
rect 3384 29044 3390 29096
rect 3694 29044 3700 29096
rect 3752 29044 3758 29096
rect 4706 29044 4712 29096
rect 4764 29044 4770 29096
rect 4798 29044 4804 29096
rect 4856 29084 4862 29096
rect 6840 29084 6868 29112
rect 4856 29056 6868 29084
rect 4856 29044 4862 29056
rect 7098 29044 7104 29096
rect 7156 29084 7162 29096
rect 9048 29084 9076 29115
rect 9398 29112 9404 29164
rect 9456 29112 9462 29164
rect 10597 29155 10655 29161
rect 10597 29152 10609 29155
rect 9508 29124 10609 29152
rect 9508 29093 9536 29124
rect 10597 29121 10609 29124
rect 10643 29121 10655 29155
rect 10597 29115 10655 29121
rect 12161 29155 12219 29161
rect 12161 29121 12173 29155
rect 12207 29152 12219 29155
rect 12452 29152 12480 29183
rect 13354 29180 13360 29232
rect 13412 29220 13418 29232
rect 13412 29192 13846 29220
rect 13412 29180 13418 29192
rect 18322 29180 18328 29232
rect 18380 29180 18386 29232
rect 19334 29220 19340 29232
rect 18892 29192 19340 29220
rect 12894 29152 12900 29164
rect 12207 29124 12900 29152
rect 12207 29121 12219 29124
rect 12161 29115 12219 29121
rect 12894 29112 12900 29124
rect 12952 29112 12958 29164
rect 18892 29161 18920 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 20180 29220 20208 29260
rect 20254 29248 20260 29300
rect 20312 29248 20318 29300
rect 20346 29248 20352 29300
rect 20404 29248 20410 29300
rect 20714 29288 20720 29300
rect 20548 29260 20720 29288
rect 20548 29220 20576 29260
rect 20714 29248 20720 29260
rect 20772 29248 20778 29300
rect 21082 29248 21088 29300
rect 21140 29288 21146 29300
rect 24302 29288 24308 29300
rect 21140 29260 24308 29288
rect 21140 29248 21146 29260
rect 24302 29248 24308 29260
rect 24360 29248 24366 29300
rect 24670 29248 24676 29300
rect 24728 29288 24734 29300
rect 26418 29288 26424 29300
rect 24728 29260 24992 29288
rect 24728 29248 24734 29260
rect 20180 29192 20576 29220
rect 19150 29161 19156 29164
rect 15197 29155 15255 29161
rect 15197 29121 15209 29155
rect 15243 29121 15255 29155
rect 15197 29115 15255 29121
rect 18877 29155 18935 29161
rect 18877 29121 18889 29155
rect 18923 29121 18935 29155
rect 19144 29152 19156 29161
rect 19111 29124 19156 29152
rect 18877 29115 18935 29121
rect 19144 29115 19156 29124
rect 7156 29056 9076 29084
rect 9493 29087 9551 29093
rect 7156 29044 7162 29056
rect 9493 29053 9505 29087
rect 9539 29053 9551 29087
rect 9861 29087 9919 29093
rect 9861 29084 9873 29087
rect 9493 29047 9551 29053
rect 9784 29056 9873 29084
rect 8110 28976 8116 29028
rect 8168 29016 8174 29028
rect 9784 29025 9812 29056
rect 9861 29053 9873 29056
rect 9907 29053 9919 29087
rect 9861 29047 9919 29053
rect 11238 29044 11244 29096
rect 11296 29084 11302 29096
rect 11296 29056 12434 29084
rect 11296 29044 11302 29056
rect 8573 29019 8631 29025
rect 8573 29016 8585 29019
rect 8168 28988 8585 29016
rect 8168 28976 8174 28988
rect 8573 28985 8585 28988
rect 8619 28985 8631 29019
rect 8573 28979 8631 28985
rect 9769 29019 9827 29025
rect 9769 28985 9781 29019
rect 9815 28985 9827 29019
rect 9769 28979 9827 28985
rect 2958 28908 2964 28960
rect 3016 28948 3022 28960
rect 4065 28951 4123 28957
rect 4065 28948 4077 28951
rect 3016 28920 4077 28948
rect 3016 28908 3022 28920
rect 4065 28917 4077 28920
rect 4111 28917 4123 28951
rect 4065 28911 4123 28917
rect 6178 28908 6184 28960
rect 6236 28908 6242 28960
rect 10502 28908 10508 28960
rect 10560 28908 10566 28960
rect 12406 28957 12434 29056
rect 12618 29044 12624 29096
rect 12676 29084 12682 29096
rect 13081 29087 13139 29093
rect 13081 29084 13093 29087
rect 12676 29056 13093 29084
rect 12676 29044 12682 29056
rect 13081 29053 13093 29056
rect 13127 29053 13139 29087
rect 13081 29047 13139 29053
rect 13357 29087 13415 29093
rect 13357 29053 13369 29087
rect 13403 29084 13415 29087
rect 13998 29084 14004 29096
rect 13403 29056 14004 29084
rect 13403 29053 13415 29056
rect 13357 29047 13415 29053
rect 12397 28951 12455 28957
rect 12397 28917 12409 28951
rect 12443 28917 12455 28951
rect 13096 28948 13124 29047
rect 13998 29044 14004 29056
rect 14056 29044 14062 29096
rect 15212 29028 15240 29115
rect 19150 29112 19156 29115
rect 19208 29112 19214 29164
rect 19702 29112 19708 29164
rect 19760 29152 19766 29164
rect 20548 29161 20576 29192
rect 20625 29223 20683 29229
rect 20625 29189 20637 29223
rect 20671 29220 20683 29223
rect 20806 29220 20812 29232
rect 20671 29192 20812 29220
rect 20671 29189 20683 29192
rect 20625 29183 20683 29189
rect 20806 29180 20812 29192
rect 20864 29180 20870 29232
rect 21910 29220 21916 29232
rect 21284 29192 21916 29220
rect 20533 29155 20591 29161
rect 19760 29124 20484 29152
rect 19760 29112 19766 29124
rect 20456 29084 20484 29124
rect 20533 29121 20545 29155
rect 20579 29121 20591 29155
rect 20533 29115 20591 29121
rect 20717 29155 20775 29161
rect 20717 29121 20729 29155
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 20732 29084 20760 29115
rect 20898 29112 20904 29164
rect 20956 29112 20962 29164
rect 21174 29112 21180 29164
rect 21232 29112 21238 29164
rect 21284 29084 21312 29192
rect 21910 29180 21916 29192
rect 21968 29220 21974 29232
rect 22005 29223 22063 29229
rect 22005 29220 22017 29223
rect 21968 29192 22017 29220
rect 21968 29180 21974 29192
rect 22005 29189 22017 29192
rect 22051 29189 22063 29223
rect 22005 29183 22063 29189
rect 22097 29223 22155 29229
rect 22097 29189 22109 29223
rect 22143 29220 22155 29223
rect 23106 29220 23112 29232
rect 22143 29192 23112 29220
rect 22143 29189 22155 29192
rect 22097 29183 22155 29189
rect 23106 29180 23112 29192
rect 23164 29180 23170 29232
rect 23385 29223 23443 29229
rect 23385 29189 23397 29223
rect 23431 29220 23443 29223
rect 23474 29220 23480 29232
rect 23431 29192 23480 29220
rect 23431 29189 23443 29192
rect 23385 29183 23443 29189
rect 23474 29180 23480 29192
rect 23532 29220 23538 29232
rect 24026 29220 24032 29232
rect 23532 29192 24032 29220
rect 23532 29180 23538 29192
rect 24026 29180 24032 29192
rect 24084 29180 24090 29232
rect 24964 29220 24992 29260
rect 25240 29260 26424 29288
rect 25240 29220 25268 29260
rect 26418 29248 26424 29260
rect 26476 29248 26482 29300
rect 26510 29248 26516 29300
rect 26568 29248 26574 29300
rect 29733 29291 29791 29297
rect 29733 29257 29745 29291
rect 29779 29288 29791 29291
rect 29822 29288 29828 29300
rect 29779 29260 29828 29288
rect 29779 29257 29791 29260
rect 29733 29251 29791 29257
rect 29822 29248 29828 29260
rect 29880 29288 29886 29300
rect 30006 29288 30012 29300
rect 29880 29260 30012 29288
rect 29880 29248 29886 29260
rect 30006 29248 30012 29260
rect 30064 29248 30070 29300
rect 30834 29248 30840 29300
rect 30892 29248 30898 29300
rect 32677 29291 32735 29297
rect 32677 29257 32689 29291
rect 32723 29257 32735 29291
rect 32677 29251 32735 29257
rect 24886 29192 25268 29220
rect 25317 29223 25375 29229
rect 25317 29189 25329 29223
rect 25363 29220 25375 29223
rect 25685 29223 25743 29229
rect 25685 29220 25697 29223
rect 25363 29192 25697 29220
rect 25363 29189 25375 29192
rect 25317 29183 25375 29189
rect 25685 29189 25697 29192
rect 25731 29189 25743 29223
rect 25685 29183 25743 29189
rect 28261 29223 28319 29229
rect 28261 29189 28273 29223
rect 28307 29220 28319 29223
rect 28534 29220 28540 29232
rect 28307 29192 28540 29220
rect 28307 29189 28319 29192
rect 28261 29183 28319 29189
rect 28534 29180 28540 29192
rect 28592 29180 28598 29232
rect 29270 29180 29276 29232
rect 29328 29180 29334 29232
rect 30374 29180 30380 29232
rect 30432 29220 30438 29232
rect 30469 29223 30527 29229
rect 30469 29220 30481 29223
rect 30432 29192 30481 29220
rect 30432 29180 30438 29192
rect 30469 29189 30481 29192
rect 30515 29189 30527 29223
rect 30852 29220 30880 29248
rect 32692 29220 32720 29251
rect 32858 29248 32864 29300
rect 32916 29288 32922 29300
rect 33045 29291 33103 29297
rect 33045 29288 33057 29291
rect 32916 29260 33057 29288
rect 32916 29248 32922 29260
rect 33045 29257 33057 29260
rect 33091 29257 33103 29291
rect 33045 29251 33103 29257
rect 33870 29248 33876 29300
rect 33928 29248 33934 29300
rect 34330 29248 34336 29300
rect 34388 29288 34394 29300
rect 34517 29291 34575 29297
rect 34517 29288 34529 29291
rect 34388 29260 34529 29288
rect 34388 29248 34394 29260
rect 34517 29257 34529 29260
rect 34563 29257 34575 29291
rect 34517 29251 34575 29257
rect 36630 29248 36636 29300
rect 36688 29288 36694 29300
rect 36688 29260 37044 29288
rect 36688 29248 36694 29260
rect 33134 29220 33140 29232
rect 30852 29192 30958 29220
rect 32692 29192 33140 29220
rect 30469 29183 30527 29189
rect 33134 29180 33140 29192
rect 33192 29180 33198 29232
rect 33505 29223 33563 29229
rect 33505 29220 33517 29223
rect 33428 29192 33517 29220
rect 21634 29112 21640 29164
rect 21692 29152 21698 29164
rect 21821 29155 21879 29161
rect 21692 29124 21772 29152
rect 21692 29112 21698 29124
rect 20456 29056 21312 29084
rect 15194 29016 15200 29028
rect 14752 28988 15200 29016
rect 14752 28948 14780 28988
rect 15194 28976 15200 28988
rect 15252 28976 15258 29028
rect 18138 28976 18144 29028
rect 18196 28976 18202 29028
rect 21174 28976 21180 29028
rect 21232 29016 21238 29028
rect 21453 29019 21511 29025
rect 21453 29016 21465 29019
rect 21232 28988 21465 29016
rect 21232 28976 21238 28988
rect 21453 28985 21465 28988
rect 21499 29016 21511 29019
rect 21634 29016 21640 29028
rect 21499 28988 21640 29016
rect 21499 28985 21511 28988
rect 21453 28979 21511 28985
rect 21634 28976 21640 28988
rect 21692 28976 21698 29028
rect 21744 29016 21772 29124
rect 21821 29121 21833 29155
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29121 22247 29155
rect 22649 29155 22707 29161
rect 22649 29152 22661 29155
rect 22189 29115 22247 29121
rect 22296 29124 22661 29152
rect 21836 29084 21864 29115
rect 22094 29084 22100 29096
rect 21836 29056 22100 29084
rect 22094 29044 22100 29056
rect 22152 29044 22158 29096
rect 21744 28988 21956 29016
rect 13096 28920 14780 28948
rect 21928 28948 21956 28988
rect 22002 28976 22008 29028
rect 22060 29016 22066 29028
rect 22204 29016 22232 29115
rect 22060 28988 22232 29016
rect 22296 29016 22324 29124
rect 22649 29121 22661 29124
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 23566 29112 23572 29164
rect 23624 29112 23630 29164
rect 26786 29112 26792 29164
rect 26844 29152 26850 29164
rect 26844 29124 27660 29152
rect 26844 29112 26850 29124
rect 27632 29096 27660 29124
rect 30190 29112 30196 29164
rect 30248 29112 30254 29164
rect 32766 29112 32772 29164
rect 32824 29152 32830 29164
rect 33428 29152 33456 29192
rect 33505 29189 33517 29192
rect 33551 29189 33563 29223
rect 33505 29183 33563 29189
rect 33594 29180 33600 29232
rect 33652 29220 33658 29232
rect 33705 29223 33763 29229
rect 33705 29220 33717 29223
rect 33652 29192 33717 29220
rect 33652 29180 33658 29192
rect 33705 29189 33717 29192
rect 33751 29189 33763 29223
rect 33705 29183 33763 29189
rect 34146 29180 34152 29232
rect 34204 29220 34210 29232
rect 34204 29192 34376 29220
rect 34204 29180 34210 29192
rect 34348 29161 34376 29192
rect 35986 29180 35992 29232
rect 36044 29220 36050 29232
rect 36449 29223 36507 29229
rect 36449 29220 36461 29223
rect 36044 29192 36461 29220
rect 36044 29180 36050 29192
rect 36449 29189 36461 29192
rect 36495 29220 36507 29223
rect 36495 29192 36952 29220
rect 36495 29189 36507 29192
rect 36449 29183 36507 29189
rect 32824 29124 33456 29152
rect 32824 29112 32830 29124
rect 22833 29087 22891 29093
rect 22833 29053 22845 29087
rect 22879 29053 22891 29087
rect 22833 29047 22891 29053
rect 23753 29087 23811 29093
rect 23753 29053 23765 29087
rect 23799 29084 23811 29087
rect 25222 29084 25228 29096
rect 23799 29056 25228 29084
rect 23799 29053 23811 29056
rect 23753 29047 23811 29053
rect 22373 29019 22431 29025
rect 22373 29016 22385 29019
rect 22296 28988 22385 29016
rect 22060 28976 22066 28988
rect 22373 28985 22385 28988
rect 22419 28985 22431 29019
rect 22373 28979 22431 28985
rect 22462 28976 22468 29028
rect 22520 28976 22526 29028
rect 22848 29016 22876 29047
rect 25222 29044 25228 29056
rect 25280 29044 25286 29096
rect 25590 29044 25596 29096
rect 25648 29044 25654 29096
rect 26326 29044 26332 29096
rect 26384 29044 26390 29096
rect 27525 29087 27583 29093
rect 27525 29053 27537 29087
rect 27571 29053 27583 29087
rect 27525 29047 27583 29053
rect 22572 28988 22876 29016
rect 23845 29019 23903 29025
rect 22572 28948 22600 28988
rect 23845 28985 23857 29019
rect 23891 29016 23903 29019
rect 24118 29016 24124 29028
rect 23891 28988 24124 29016
rect 23891 28985 23903 28988
rect 23845 28979 23903 28985
rect 24118 28976 24124 28988
rect 24176 28976 24182 29028
rect 25774 28976 25780 29028
rect 25832 29016 25838 29028
rect 27540 29016 27568 29047
rect 27614 29044 27620 29096
rect 27672 29084 27678 29096
rect 27985 29087 28043 29093
rect 27985 29084 27997 29087
rect 27672 29056 27997 29084
rect 27672 29044 27678 29056
rect 27985 29053 27997 29056
rect 28031 29053 28043 29087
rect 27985 29047 28043 29053
rect 31478 29044 31484 29096
rect 31536 29084 31542 29096
rect 32401 29087 32459 29093
rect 32401 29084 32413 29087
rect 31536 29056 32413 29084
rect 31536 29044 31542 29056
rect 32401 29053 32413 29056
rect 32447 29053 32459 29087
rect 32401 29047 32459 29053
rect 32493 29087 32551 29093
rect 32493 29053 32505 29087
rect 32539 29053 32551 29087
rect 32493 29047 32551 29053
rect 32861 29087 32919 29093
rect 32861 29053 32873 29087
rect 32907 29084 32919 29087
rect 33042 29084 33048 29096
rect 32907 29056 33048 29084
rect 32907 29053 32919 29056
rect 32861 29047 32919 29053
rect 32508 29016 32536 29047
rect 33042 29044 33048 29056
rect 33100 29044 33106 29096
rect 25832 28988 27568 29016
rect 31956 28988 32536 29016
rect 33428 29016 33456 29124
rect 34333 29155 34391 29161
rect 34333 29121 34345 29155
rect 34379 29152 34391 29155
rect 34422 29152 34428 29164
rect 34379 29124 34428 29152
rect 34379 29121 34391 29124
rect 34333 29115 34391 29121
rect 34422 29112 34428 29124
rect 34480 29112 34486 29164
rect 34606 29112 34612 29164
rect 34664 29112 34670 29164
rect 36630 29112 36636 29164
rect 36688 29112 36694 29164
rect 36924 29161 36952 29192
rect 36909 29155 36967 29161
rect 36909 29121 36921 29155
rect 36955 29121 36967 29155
rect 37016 29152 37044 29260
rect 37093 29155 37151 29161
rect 37093 29152 37105 29155
rect 37016 29124 37105 29152
rect 36909 29115 36967 29121
rect 37093 29121 37105 29124
rect 37139 29121 37151 29155
rect 37093 29115 37151 29121
rect 37182 29112 37188 29164
rect 37240 29152 37246 29164
rect 37461 29155 37519 29161
rect 37461 29152 37473 29155
rect 37240 29124 37473 29152
rect 37240 29112 37246 29124
rect 37461 29121 37473 29124
rect 37507 29121 37519 29155
rect 37461 29115 37519 29121
rect 34054 29044 34060 29096
rect 34112 29044 34118 29096
rect 34149 29087 34207 29093
rect 34149 29053 34161 29087
rect 34195 29053 34207 29087
rect 34149 29047 34207 29053
rect 34241 29087 34299 29093
rect 34241 29053 34253 29087
rect 34287 29053 34299 29087
rect 34241 29047 34299 29053
rect 34164 29016 34192 29047
rect 33428 28988 34192 29016
rect 34256 29016 34284 29047
rect 35434 29044 35440 29096
rect 35492 29044 35498 29096
rect 37369 29087 37427 29093
rect 37369 29084 37381 29087
rect 36832 29056 37381 29084
rect 34330 29016 34336 29028
rect 34256 28988 34336 29016
rect 25832 28976 25838 28988
rect 21928 28920 22600 28948
rect 12397 28911 12455 28917
rect 26234 28908 26240 28960
rect 26292 28948 26298 28960
rect 26973 28951 27031 28957
rect 26973 28948 26985 28951
rect 26292 28920 26985 28948
rect 26292 28908 26298 28920
rect 26973 28917 26985 28920
rect 27019 28917 27031 28951
rect 26973 28911 27031 28917
rect 31846 28908 31852 28960
rect 31904 28948 31910 28960
rect 31956 28957 31984 28988
rect 31941 28951 31999 28957
rect 31941 28948 31953 28951
rect 31904 28920 31953 28948
rect 31904 28908 31910 28920
rect 31941 28917 31953 28920
rect 31987 28917 31999 28951
rect 31941 28911 31999 28917
rect 33134 28908 33140 28960
rect 33192 28948 33198 28960
rect 33689 28951 33747 28957
rect 33689 28948 33701 28951
rect 33192 28920 33701 28948
rect 33192 28908 33198 28920
rect 33689 28917 33701 28920
rect 33735 28948 33747 28951
rect 34054 28948 34060 28960
rect 33735 28920 34060 28948
rect 33735 28917 33747 28920
rect 33689 28911 33747 28917
rect 34054 28908 34060 28920
rect 34112 28908 34118 28960
rect 34164 28948 34192 28988
rect 34330 28976 34336 28988
rect 34388 28976 34394 29028
rect 36832 28960 36860 29056
rect 37369 29053 37381 29056
rect 37415 29053 37427 29087
rect 37369 29047 37427 29053
rect 34790 28948 34796 28960
rect 34164 28920 34796 28948
rect 34790 28908 34796 28920
rect 34848 28908 34854 28960
rect 36814 28908 36820 28960
rect 36872 28908 36878 28960
rect 36998 28908 37004 28960
rect 37056 28908 37062 28960
rect 37642 28908 37648 28960
rect 37700 28948 37706 28960
rect 37737 28951 37795 28957
rect 37737 28948 37749 28951
rect 37700 28920 37749 28948
rect 37700 28908 37706 28920
rect 37737 28917 37749 28920
rect 37783 28917 37795 28951
rect 37737 28911 37795 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 3145 28747 3203 28753
rect 3145 28713 3157 28747
rect 3191 28744 3203 28747
rect 3694 28744 3700 28756
rect 3191 28716 3700 28744
rect 3191 28713 3203 28716
rect 3145 28707 3203 28713
rect 3694 28704 3700 28716
rect 3752 28704 3758 28756
rect 3973 28747 4031 28753
rect 3973 28713 3985 28747
rect 4019 28744 4031 28747
rect 7377 28747 7435 28753
rect 4019 28716 4384 28744
rect 4019 28713 4031 28716
rect 3973 28707 4031 28713
rect 4062 28676 4068 28688
rect 3620 28648 4068 28676
rect 3620 28552 3648 28648
rect 4062 28636 4068 28648
rect 4120 28636 4126 28688
rect 4356 28676 4384 28716
rect 7377 28713 7389 28747
rect 7423 28744 7435 28747
rect 7466 28744 7472 28756
rect 7423 28716 7472 28744
rect 7423 28713 7435 28716
rect 7377 28707 7435 28713
rect 7466 28704 7472 28716
rect 7524 28704 7530 28756
rect 7561 28747 7619 28753
rect 7561 28713 7573 28747
rect 7607 28744 7619 28747
rect 8202 28744 8208 28756
rect 7607 28716 8208 28744
rect 7607 28713 7619 28716
rect 7561 28707 7619 28713
rect 4356 28648 4936 28676
rect 3712 28580 4476 28608
rect 2958 28500 2964 28552
rect 3016 28500 3022 28552
rect 3145 28543 3203 28549
rect 3145 28509 3157 28543
rect 3191 28509 3203 28543
rect 3145 28503 3203 28509
rect 3160 28472 3188 28503
rect 3326 28500 3332 28552
rect 3384 28500 3390 28552
rect 3421 28543 3479 28549
rect 3421 28509 3433 28543
rect 3467 28540 3479 28543
rect 3602 28540 3608 28552
rect 3467 28512 3608 28540
rect 3467 28509 3479 28512
rect 3421 28503 3479 28509
rect 3602 28500 3608 28512
rect 3660 28500 3666 28552
rect 3712 28472 3740 28580
rect 3786 28500 3792 28552
rect 3844 28500 3850 28552
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28509 4031 28543
rect 3973 28503 4031 28509
rect 3160 28444 3740 28472
rect 3605 28407 3663 28413
rect 3605 28373 3617 28407
rect 3651 28404 3663 28407
rect 3712 28404 3740 28444
rect 3651 28376 3740 28404
rect 3988 28404 4016 28503
rect 4062 28500 4068 28552
rect 4120 28500 4126 28552
rect 4448 28472 4476 28580
rect 4798 28568 4804 28620
rect 4856 28568 4862 28620
rect 4908 28608 4936 28648
rect 7006 28636 7012 28688
rect 7064 28676 7070 28688
rect 7576 28676 7604 28707
rect 8202 28704 8208 28716
rect 8260 28704 8266 28756
rect 11057 28747 11115 28753
rect 11057 28713 11069 28747
rect 11103 28744 11115 28747
rect 11238 28744 11244 28756
rect 11103 28716 11244 28744
rect 11103 28713 11115 28716
rect 11057 28707 11115 28713
rect 11238 28704 11244 28716
rect 11296 28704 11302 28756
rect 12894 28704 12900 28756
rect 12952 28704 12958 28756
rect 21821 28747 21879 28753
rect 21821 28713 21833 28747
rect 21867 28744 21879 28747
rect 21910 28744 21916 28756
rect 21867 28716 21916 28744
rect 21867 28713 21879 28716
rect 21821 28707 21879 28713
rect 21910 28704 21916 28716
rect 21968 28704 21974 28756
rect 25774 28704 25780 28756
rect 25832 28744 25838 28756
rect 26053 28747 26111 28753
rect 26053 28744 26065 28747
rect 25832 28716 26065 28744
rect 25832 28704 25838 28716
rect 26053 28713 26065 28716
rect 26099 28713 26111 28747
rect 26053 28707 26111 28713
rect 30006 28704 30012 28756
rect 30064 28744 30070 28756
rect 30377 28747 30435 28753
rect 30064 28716 30328 28744
rect 30064 28704 30070 28716
rect 7064 28648 7604 28676
rect 13648 28648 16068 28676
rect 7064 28636 7070 28648
rect 5077 28611 5135 28617
rect 5077 28608 5089 28611
rect 4908 28580 5089 28608
rect 5077 28577 5089 28580
rect 5123 28577 5135 28611
rect 5077 28571 5135 28577
rect 6549 28611 6607 28617
rect 6549 28577 6561 28611
rect 6595 28608 6607 28611
rect 6730 28608 6736 28620
rect 6595 28580 6736 28608
rect 6595 28577 6607 28580
rect 6549 28571 6607 28577
rect 6730 28568 6736 28580
rect 6788 28608 6794 28620
rect 7193 28611 7251 28617
rect 7193 28608 7205 28611
rect 6788 28580 7205 28608
rect 6788 28568 6794 28580
rect 7193 28577 7205 28580
rect 7239 28577 7251 28611
rect 7193 28571 7251 28577
rect 7374 28568 7380 28620
rect 7432 28608 7438 28620
rect 8389 28611 8447 28617
rect 8389 28608 8401 28611
rect 7432 28580 8401 28608
rect 7432 28568 7438 28580
rect 8389 28577 8401 28580
rect 8435 28577 8447 28611
rect 8389 28571 8447 28577
rect 8938 28568 8944 28620
rect 8996 28608 9002 28620
rect 9309 28611 9367 28617
rect 9309 28608 9321 28611
rect 8996 28580 9321 28608
rect 8996 28568 9002 28580
rect 9309 28577 9321 28580
rect 9355 28577 9367 28611
rect 9309 28571 9367 28577
rect 11422 28568 11428 28620
rect 11480 28568 11486 28620
rect 13538 28568 13544 28620
rect 13596 28608 13602 28620
rect 13648 28617 13676 28648
rect 16040 28620 16068 28648
rect 24670 28636 24676 28688
rect 24728 28636 24734 28688
rect 30190 28676 30196 28688
rect 29012 28648 30196 28676
rect 13633 28611 13691 28617
rect 13633 28608 13645 28611
rect 13596 28580 13645 28608
rect 13596 28568 13602 28580
rect 13633 28577 13645 28580
rect 13679 28577 13691 28611
rect 13633 28571 13691 28577
rect 15194 28568 15200 28620
rect 15252 28568 15258 28620
rect 16022 28568 16028 28620
rect 16080 28608 16086 28620
rect 16298 28608 16304 28620
rect 16080 28580 16304 28608
rect 16080 28568 16086 28580
rect 16298 28568 16304 28580
rect 16356 28568 16362 28620
rect 23566 28568 23572 28620
rect 23624 28608 23630 28620
rect 23934 28608 23940 28620
rect 23624 28580 23940 28608
rect 23624 28568 23630 28580
rect 23934 28568 23940 28580
rect 23992 28568 23998 28620
rect 24210 28568 24216 28620
rect 24268 28608 24274 28620
rect 26510 28608 26516 28620
rect 24268 28580 24532 28608
rect 24268 28568 24274 28580
rect 4706 28500 4712 28552
rect 4764 28500 4770 28552
rect 6914 28500 6920 28552
rect 6972 28540 6978 28552
rect 7929 28543 7987 28549
rect 7929 28540 7941 28543
rect 6972 28512 7941 28540
rect 6972 28500 6978 28512
rect 7929 28509 7941 28512
rect 7975 28540 7987 28543
rect 8110 28540 8116 28552
rect 7975 28512 8116 28540
rect 7975 28509 7987 28512
rect 7929 28503 7987 28509
rect 8110 28500 8116 28512
rect 8168 28500 8174 28552
rect 11146 28500 11152 28552
rect 11204 28500 11210 28552
rect 13354 28540 13360 28552
rect 12558 28512 13360 28540
rect 13354 28500 13360 28512
rect 13412 28500 13418 28552
rect 15212 28540 15240 28568
rect 16942 28540 16948 28552
rect 15212 28512 16948 28540
rect 16942 28500 16948 28512
rect 17000 28540 17006 28552
rect 17037 28543 17095 28549
rect 17037 28540 17049 28543
rect 17000 28512 17049 28540
rect 17000 28500 17006 28512
rect 17037 28509 17049 28512
rect 17083 28509 17095 28543
rect 17037 28503 17095 28509
rect 21542 28500 21548 28552
rect 21600 28540 21606 28552
rect 21729 28543 21787 28549
rect 21729 28540 21741 28543
rect 21600 28512 21741 28540
rect 21600 28500 21606 28512
rect 21729 28509 21741 28512
rect 21775 28509 21787 28543
rect 21729 28503 21787 28509
rect 22370 28500 22376 28552
rect 22428 28500 22434 28552
rect 22557 28543 22615 28549
rect 22557 28509 22569 28543
rect 22603 28509 22615 28543
rect 22557 28503 22615 28509
rect 5166 28472 5172 28484
rect 4448 28444 5172 28472
rect 5166 28432 5172 28444
rect 5224 28432 5230 28484
rect 5810 28432 5816 28484
rect 5868 28432 5874 28484
rect 7466 28472 7472 28484
rect 6472 28444 7472 28472
rect 5442 28404 5448 28416
rect 3988 28376 5448 28404
rect 3651 28373 3663 28376
rect 3605 28367 3663 28373
rect 5442 28364 5448 28376
rect 5500 28404 5506 28416
rect 6472 28404 6500 28444
rect 7466 28432 7472 28444
rect 7524 28472 7530 28484
rect 7561 28475 7619 28481
rect 7561 28472 7573 28475
rect 7524 28444 7573 28472
rect 7524 28432 7530 28444
rect 7561 28441 7573 28444
rect 7607 28472 7619 28475
rect 8021 28475 8079 28481
rect 8021 28472 8033 28475
rect 7607 28444 8033 28472
rect 7607 28441 7619 28444
rect 7561 28435 7619 28441
rect 8021 28441 8033 28444
rect 8067 28441 8079 28475
rect 8021 28435 8079 28441
rect 8202 28432 8208 28484
rect 8260 28432 8266 28484
rect 9582 28432 9588 28484
rect 9640 28432 9646 28484
rect 10226 28432 10232 28484
rect 10284 28432 10290 28484
rect 13446 28432 13452 28484
rect 13504 28432 13510 28484
rect 14369 28475 14427 28481
rect 14369 28441 14381 28475
rect 14415 28441 14427 28475
rect 14369 28435 14427 28441
rect 17313 28475 17371 28481
rect 17313 28441 17325 28475
rect 17359 28472 17371 28475
rect 17586 28472 17592 28484
rect 17359 28444 17592 28472
rect 17359 28441 17371 28444
rect 17313 28435 17371 28441
rect 5500 28376 6500 28404
rect 5500 28364 5506 28376
rect 6638 28364 6644 28416
rect 6696 28364 6702 28416
rect 12986 28364 12992 28416
rect 13044 28364 13050 28416
rect 13357 28407 13415 28413
rect 13357 28373 13369 28407
rect 13403 28404 13415 28407
rect 13906 28404 13912 28416
rect 13403 28376 13912 28404
rect 13403 28373 13415 28376
rect 13357 28367 13415 28373
rect 13906 28364 13912 28376
rect 13964 28364 13970 28416
rect 14182 28364 14188 28416
rect 14240 28404 14246 28416
rect 14384 28404 14412 28435
rect 17586 28432 17592 28444
rect 17644 28432 17650 28484
rect 17954 28432 17960 28484
rect 18012 28432 18018 28484
rect 19058 28432 19064 28484
rect 19116 28432 19122 28484
rect 22572 28472 22600 28503
rect 22646 28500 22652 28552
rect 22704 28500 22710 28552
rect 24504 28549 24532 28580
rect 24964 28580 26516 28608
rect 24964 28549 24992 28580
rect 26510 28568 26516 28580
rect 26568 28568 26574 28620
rect 27525 28611 27583 28617
rect 27525 28577 27537 28611
rect 27571 28608 27583 28611
rect 27893 28611 27951 28617
rect 27893 28608 27905 28611
rect 27571 28580 27905 28608
rect 27571 28577 27583 28580
rect 27525 28571 27583 28577
rect 27893 28577 27905 28580
rect 27939 28577 27951 28611
rect 27893 28571 27951 28577
rect 29012 28552 29040 28648
rect 30190 28636 30196 28648
rect 30248 28636 30254 28688
rect 30300 28676 30328 28716
rect 30377 28713 30389 28747
rect 30423 28744 30435 28747
rect 30466 28744 30472 28756
rect 30423 28716 30472 28744
rect 30423 28713 30435 28716
rect 30377 28707 30435 28713
rect 30466 28704 30472 28716
rect 30524 28704 30530 28756
rect 31297 28747 31355 28753
rect 31297 28713 31309 28747
rect 31343 28744 31355 28747
rect 31478 28744 31484 28756
rect 31343 28716 31484 28744
rect 31343 28713 31355 28716
rect 31297 28707 31355 28713
rect 31478 28704 31484 28716
rect 31536 28704 31542 28756
rect 31662 28704 31668 28756
rect 31720 28744 31726 28756
rect 34517 28747 34575 28753
rect 34517 28744 34529 28747
rect 31720 28716 34529 28744
rect 31720 28704 31726 28716
rect 34517 28713 34529 28716
rect 34563 28744 34575 28747
rect 34606 28744 34612 28756
rect 34563 28716 34612 28744
rect 34563 28713 34575 28716
rect 34517 28707 34575 28713
rect 34606 28704 34612 28716
rect 34664 28704 34670 28756
rect 34793 28747 34851 28753
rect 34793 28713 34805 28747
rect 34839 28744 34851 28747
rect 34882 28744 34888 28756
rect 34839 28716 34888 28744
rect 34839 28713 34851 28716
rect 34793 28707 34851 28713
rect 34882 28704 34888 28716
rect 34940 28704 34946 28756
rect 34977 28747 35035 28753
rect 34977 28713 34989 28747
rect 35023 28744 35035 28747
rect 35023 28716 35664 28744
rect 35023 28713 35035 28716
rect 34977 28707 35035 28713
rect 33689 28679 33747 28685
rect 30300 28648 31248 28676
rect 29641 28611 29699 28617
rect 29641 28608 29653 28611
rect 29104 28580 29653 28608
rect 22741 28543 22799 28549
rect 22741 28509 22753 28543
rect 22787 28540 22799 28543
rect 23385 28543 23443 28549
rect 23385 28540 23397 28543
rect 22787 28512 23397 28540
rect 22787 28509 22799 28512
rect 22741 28503 22799 28509
rect 23385 28509 23397 28512
rect 23431 28509 23443 28543
rect 23385 28503 23443 28509
rect 24489 28543 24547 28549
rect 24489 28509 24501 28543
rect 24535 28509 24547 28543
rect 24489 28503 24547 28509
rect 24949 28543 25007 28549
rect 24949 28509 24961 28543
rect 24995 28509 25007 28543
rect 24949 28503 25007 28509
rect 26418 28500 26424 28552
rect 26476 28500 26482 28552
rect 27801 28543 27859 28549
rect 27801 28509 27813 28543
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 22922 28472 22928 28484
rect 22572 28444 22928 28472
rect 22922 28432 22928 28444
rect 22980 28432 22986 28484
rect 24210 28432 24216 28484
rect 24268 28472 24274 28484
rect 25590 28472 25596 28484
rect 24268 28444 25596 28472
rect 24268 28432 24274 28444
rect 25590 28432 25596 28444
rect 25648 28472 25654 28484
rect 25685 28475 25743 28481
rect 25685 28472 25697 28475
rect 25648 28444 25697 28472
rect 25648 28432 25654 28444
rect 25685 28441 25697 28444
rect 25731 28441 25743 28475
rect 27816 28472 27844 28503
rect 28442 28500 28448 28552
rect 28500 28500 28506 28552
rect 28905 28543 28963 28549
rect 28905 28509 28917 28543
rect 28951 28509 28963 28543
rect 28905 28503 28963 28509
rect 25685 28435 25743 28441
rect 27632 28444 27844 28472
rect 28920 28472 28948 28503
rect 28994 28500 29000 28552
rect 29052 28500 29058 28552
rect 29104 28549 29132 28580
rect 29641 28577 29653 28580
rect 29687 28577 29699 28611
rect 30101 28611 30159 28617
rect 30101 28608 30113 28611
rect 29641 28571 29699 28577
rect 29840 28580 30113 28608
rect 29089 28543 29147 28549
rect 29089 28509 29101 28543
rect 29135 28509 29147 28543
rect 29089 28503 29147 28509
rect 29178 28500 29184 28552
rect 29236 28540 29242 28552
rect 29273 28543 29331 28549
rect 29273 28540 29285 28543
rect 29236 28512 29285 28540
rect 29236 28500 29242 28512
rect 29273 28509 29285 28512
rect 29319 28509 29331 28543
rect 29273 28503 29331 28509
rect 29730 28500 29736 28552
rect 29788 28500 29794 28552
rect 29840 28472 29868 28580
rect 30101 28577 30113 28580
rect 30147 28608 30159 28611
rect 30837 28611 30895 28617
rect 30837 28608 30849 28611
rect 30147 28580 30849 28608
rect 30147 28577 30159 28580
rect 30101 28571 30159 28577
rect 30837 28577 30849 28580
rect 30883 28608 30895 28611
rect 30883 28580 30972 28608
rect 30883 28577 30895 28580
rect 30837 28571 30895 28577
rect 29917 28543 29975 28549
rect 29917 28509 29929 28543
rect 29963 28509 29975 28543
rect 29917 28503 29975 28509
rect 28920 28444 29868 28472
rect 29932 28472 29960 28503
rect 30006 28500 30012 28552
rect 30064 28500 30070 28552
rect 30190 28500 30196 28552
rect 30248 28540 30254 28552
rect 30944 28549 30972 28580
rect 31110 28568 31116 28620
rect 31168 28568 31174 28620
rect 30653 28543 30711 28549
rect 30653 28540 30665 28543
rect 30248 28512 30665 28540
rect 30248 28500 30254 28512
rect 30653 28509 30665 28512
rect 30699 28509 30711 28543
rect 30653 28503 30711 28509
rect 30929 28543 30987 28549
rect 30929 28509 30941 28543
rect 30975 28509 30987 28543
rect 31128 28540 31156 28568
rect 30929 28503 30987 28509
rect 31036 28512 31156 28540
rect 30742 28472 30748 28484
rect 29932 28444 30748 28472
rect 14240 28376 14412 28404
rect 15381 28407 15439 28413
rect 14240 28364 14246 28376
rect 15381 28373 15393 28407
rect 15427 28404 15439 28407
rect 15470 28404 15476 28416
rect 15427 28376 15476 28404
rect 15427 28373 15439 28376
rect 15381 28367 15439 28373
rect 15470 28364 15476 28376
rect 15528 28364 15534 28416
rect 15746 28364 15752 28416
rect 15804 28364 15810 28416
rect 15838 28364 15844 28416
rect 15896 28364 15902 28416
rect 22830 28364 22836 28416
rect 22888 28404 22894 28416
rect 23017 28407 23075 28413
rect 23017 28404 23029 28407
rect 22888 28376 23029 28404
rect 22888 28364 22894 28376
rect 23017 28373 23029 28376
rect 23063 28373 23075 28407
rect 25700 28404 25728 28435
rect 27632 28416 27660 28444
rect 29748 28416 29776 28444
rect 30742 28432 30748 28444
rect 30800 28432 30806 28484
rect 27614 28404 27620 28416
rect 25700 28376 27620 28404
rect 23017 28367 23075 28373
rect 27614 28364 27620 28376
rect 27672 28364 27678 28416
rect 28258 28364 28264 28416
rect 28316 28404 28322 28416
rect 28629 28407 28687 28413
rect 28629 28404 28641 28407
rect 28316 28376 28641 28404
rect 28316 28364 28322 28376
rect 28629 28373 28641 28376
rect 28675 28373 28687 28407
rect 28629 28367 28687 28373
rect 29730 28364 29736 28416
rect 29788 28364 29794 28416
rect 29822 28364 29828 28416
rect 29880 28404 29886 28416
rect 30469 28407 30527 28413
rect 30469 28404 30481 28407
rect 29880 28376 30481 28404
rect 29880 28364 29886 28376
rect 30469 28373 30481 28376
rect 30515 28404 30527 28407
rect 31036 28404 31064 28512
rect 31110 28432 31116 28484
rect 31168 28472 31174 28484
rect 31220 28472 31248 28648
rect 33689 28645 33701 28679
rect 33735 28676 33747 28679
rect 33962 28676 33968 28688
rect 33735 28648 33968 28676
rect 33735 28645 33747 28648
rect 33689 28639 33747 28645
rect 33962 28636 33968 28648
rect 34020 28636 34026 28688
rect 34054 28636 34060 28688
rect 34112 28676 34118 28688
rect 34992 28676 35020 28707
rect 34112 28648 35020 28676
rect 34112 28636 34118 28648
rect 35526 28636 35532 28688
rect 35584 28636 35590 28688
rect 32769 28611 32827 28617
rect 32769 28577 32781 28611
rect 32815 28608 32827 28611
rect 33502 28608 33508 28620
rect 32815 28580 33508 28608
rect 32815 28577 32827 28580
rect 32769 28571 32827 28577
rect 33502 28568 33508 28580
rect 33560 28568 33566 28620
rect 34241 28611 34299 28617
rect 34241 28608 34253 28611
rect 33796 28580 34253 28608
rect 33796 28552 33824 28580
rect 34241 28577 34253 28580
rect 34287 28608 34299 28611
rect 34330 28608 34336 28620
rect 34287 28580 34336 28608
rect 34287 28577 34299 28580
rect 34241 28571 34299 28577
rect 34330 28568 34336 28580
rect 34388 28608 34394 28620
rect 34388 28580 34744 28608
rect 34388 28568 34394 28580
rect 33134 28500 33140 28552
rect 33192 28540 33198 28552
rect 33229 28543 33287 28549
rect 33229 28540 33241 28543
rect 33192 28512 33241 28540
rect 33192 28500 33198 28512
rect 33229 28509 33241 28512
rect 33275 28509 33287 28543
rect 33229 28503 33287 28509
rect 31168 28444 31248 28472
rect 31168 28432 31174 28444
rect 32766 28432 32772 28484
rect 32824 28472 32830 28484
rect 33244 28472 33272 28503
rect 33778 28500 33784 28552
rect 33836 28500 33842 28552
rect 33962 28500 33968 28552
rect 34020 28540 34026 28552
rect 34057 28543 34115 28549
rect 34057 28540 34069 28543
rect 34020 28512 34069 28540
rect 34020 28500 34026 28512
rect 34057 28509 34069 28512
rect 34103 28540 34115 28543
rect 34146 28540 34152 28552
rect 34103 28512 34152 28540
rect 34103 28509 34115 28512
rect 34057 28503 34115 28509
rect 34146 28500 34152 28512
rect 34204 28500 34210 28552
rect 33594 28472 33600 28484
rect 32824 28444 33180 28472
rect 33244 28444 33600 28472
rect 32824 28432 32830 28444
rect 30515 28376 31064 28404
rect 30515 28373 30527 28376
rect 30469 28367 30527 28373
rect 33042 28364 33048 28416
rect 33100 28364 33106 28416
rect 33152 28413 33180 28444
rect 33594 28432 33600 28444
rect 33652 28472 33658 28484
rect 33873 28475 33931 28481
rect 33873 28472 33885 28475
rect 33652 28444 33885 28472
rect 33652 28432 33658 28444
rect 33873 28441 33885 28444
rect 33919 28472 33931 28475
rect 34330 28472 34336 28484
rect 33919 28444 34336 28472
rect 33919 28441 33931 28444
rect 33873 28435 33931 28441
rect 34330 28432 34336 28444
rect 34388 28432 34394 28484
rect 34716 28472 34744 28580
rect 34882 28568 34888 28620
rect 34940 28608 34946 28620
rect 35437 28611 35495 28617
rect 35437 28608 35449 28611
rect 34940 28580 35449 28608
rect 34940 28568 34946 28580
rect 35437 28577 35449 28580
rect 35483 28608 35495 28611
rect 35544 28608 35572 28636
rect 35483 28580 35572 28608
rect 35483 28577 35495 28580
rect 35437 28571 35495 28577
rect 34992 28512 35296 28540
rect 34992 28481 35020 28512
rect 34961 28475 35020 28481
rect 34961 28472 34973 28475
rect 34716 28444 34973 28472
rect 34961 28441 34973 28444
rect 35007 28444 35020 28475
rect 35161 28475 35219 28481
rect 35007 28441 35019 28444
rect 34961 28435 35019 28441
rect 35161 28441 35173 28475
rect 35207 28441 35219 28475
rect 35268 28472 35296 28512
rect 35342 28500 35348 28552
rect 35400 28540 35406 28552
rect 35526 28540 35532 28552
rect 35400 28512 35532 28540
rect 35400 28500 35406 28512
rect 35526 28500 35532 28512
rect 35584 28500 35590 28552
rect 35636 28540 35664 28716
rect 35986 28704 35992 28756
rect 36044 28704 36050 28756
rect 35897 28611 35955 28617
rect 35897 28577 35909 28611
rect 35943 28608 35955 28611
rect 36004 28608 36032 28704
rect 36446 28608 36452 28620
rect 35943 28580 36032 28608
rect 36096 28580 36452 28608
rect 35943 28577 35955 28580
rect 35897 28571 35955 28577
rect 36096 28540 36124 28580
rect 36446 28568 36452 28580
rect 36504 28568 36510 28620
rect 36814 28568 36820 28620
rect 36872 28568 36878 28620
rect 35636 28512 36124 28540
rect 36170 28500 36176 28552
rect 36228 28500 36234 28552
rect 36265 28543 36323 28549
rect 36265 28509 36277 28543
rect 36311 28509 36323 28543
rect 36265 28503 36323 28509
rect 36280 28472 36308 28503
rect 36354 28500 36360 28552
rect 36412 28500 36418 28552
rect 36998 28500 37004 28552
rect 37056 28500 37062 28552
rect 37458 28500 37464 28552
rect 37516 28500 37522 28552
rect 37734 28500 37740 28552
rect 37792 28500 37798 28552
rect 37918 28500 37924 28552
rect 37976 28500 37982 28552
rect 35268 28444 36308 28472
rect 37185 28475 37243 28481
rect 35161 28435 35219 28441
rect 37185 28441 37197 28475
rect 37231 28472 37243 28475
rect 37550 28472 37556 28484
rect 37231 28444 37556 28472
rect 37231 28441 37243 28444
rect 37185 28435 37243 28441
rect 33137 28407 33195 28413
rect 33137 28373 33149 28407
rect 33183 28373 33195 28407
rect 33137 28367 33195 28373
rect 33505 28407 33563 28413
rect 33505 28373 33517 28407
rect 33551 28404 33563 28407
rect 33686 28404 33692 28416
rect 33551 28376 33692 28404
rect 33551 28373 33563 28376
rect 33505 28367 33563 28373
rect 33686 28364 33692 28376
rect 33744 28364 33750 28416
rect 34790 28364 34796 28416
rect 34848 28404 34854 28416
rect 35176 28404 35204 28435
rect 37550 28432 37556 28444
rect 37608 28432 37614 28484
rect 34848 28376 35204 28404
rect 35253 28407 35311 28413
rect 34848 28364 34854 28376
rect 35253 28373 35265 28407
rect 35299 28404 35311 28407
rect 35342 28404 35348 28416
rect 35299 28376 35348 28404
rect 35299 28373 35311 28376
rect 35253 28367 35311 28373
rect 35342 28364 35348 28376
rect 35400 28364 35406 28416
rect 35526 28364 35532 28416
rect 35584 28404 35590 28416
rect 36170 28404 36176 28416
rect 35584 28376 36176 28404
rect 35584 28364 35590 28376
rect 36170 28364 36176 28376
rect 36228 28364 36234 28416
rect 37277 28407 37335 28413
rect 37277 28373 37289 28407
rect 37323 28404 37335 28407
rect 38010 28404 38016 28416
rect 37323 28376 38016 28404
rect 37323 28373 37335 28376
rect 37277 28367 37335 28373
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 1104 28314 38824 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 38824 28314
rect 1104 28240 38824 28262
rect 4893 28203 4951 28209
rect 4893 28200 4905 28203
rect 2148 28172 4905 28200
rect 2148 28141 2176 28172
rect 4893 28169 4905 28172
rect 4939 28169 4951 28203
rect 6638 28200 6644 28212
rect 4893 28163 4951 28169
rect 5368 28172 6644 28200
rect 2133 28135 2191 28141
rect 2133 28101 2145 28135
rect 2179 28101 2191 28135
rect 2133 28095 2191 28101
rect 2774 28092 2780 28144
rect 2832 28092 2838 28144
rect 3602 28092 3608 28144
rect 3660 28132 3666 28144
rect 5258 28132 5264 28144
rect 3660 28104 4844 28132
rect 3660 28092 3666 28104
rect 3970 28024 3976 28076
rect 4028 28064 4034 28076
rect 4249 28067 4307 28073
rect 4249 28064 4261 28067
rect 4028 28036 4261 28064
rect 4028 28024 4034 28036
rect 4249 28033 4261 28036
rect 4295 28033 4307 28067
rect 4249 28027 4307 28033
rect 4433 28067 4491 28073
rect 4433 28033 4445 28067
rect 4479 28033 4491 28067
rect 4433 28027 4491 28033
rect 4525 28067 4583 28073
rect 4525 28033 4537 28067
rect 4571 28064 4583 28067
rect 4614 28064 4620 28076
rect 4571 28036 4620 28064
rect 4571 28033 4583 28036
rect 4525 28027 4583 28033
rect 1394 27956 1400 28008
rect 1452 27996 1458 28008
rect 1857 27999 1915 28005
rect 1857 27996 1869 27999
rect 1452 27968 1869 27996
rect 1452 27956 1458 27968
rect 1857 27965 1869 27968
rect 1903 27965 1915 27999
rect 1857 27959 1915 27965
rect 3418 27956 3424 28008
rect 3476 27996 3482 28008
rect 3605 27999 3663 28005
rect 3605 27996 3617 27999
rect 3476 27968 3617 27996
rect 3476 27956 3482 27968
rect 3605 27965 3617 27968
rect 3651 27996 3663 27999
rect 4062 27996 4068 28008
rect 3651 27968 4068 27996
rect 3651 27965 3663 27968
rect 3605 27959 3663 27965
rect 4062 27956 4068 27968
rect 4120 27956 4126 28008
rect 3142 27888 3148 27940
rect 3200 27928 3206 27940
rect 4448 27928 4476 28027
rect 4614 28024 4620 28036
rect 4672 28024 4678 28076
rect 4706 28024 4712 28076
rect 4764 28024 4770 28076
rect 4816 28073 4844 28104
rect 5092 28104 5264 28132
rect 5092 28073 5120 28104
rect 5258 28092 5264 28104
rect 5316 28092 5322 28144
rect 5368 28141 5396 28172
rect 6638 28160 6644 28172
rect 6696 28160 6702 28212
rect 7558 28200 7564 28212
rect 7300 28172 7564 28200
rect 5353 28135 5411 28141
rect 5353 28101 5365 28135
rect 5399 28101 5411 28135
rect 5597 28135 5655 28141
rect 5597 28132 5609 28135
rect 5353 28095 5411 28101
rect 5460 28104 5609 28132
rect 4801 28067 4859 28073
rect 4801 28033 4813 28067
rect 4847 28033 4859 28067
rect 4801 28027 4859 28033
rect 4985 28067 5043 28073
rect 4985 28033 4997 28067
rect 5031 28033 5043 28067
rect 4985 28027 5043 28033
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28033 5135 28067
rect 5077 28027 5135 28033
rect 5169 28067 5227 28073
rect 5169 28033 5181 28067
rect 5215 28033 5227 28067
rect 5276 28064 5304 28092
rect 5460 28064 5488 28104
rect 5597 28101 5609 28104
rect 5643 28101 5655 28135
rect 5597 28095 5655 28101
rect 5813 28135 5871 28141
rect 5813 28101 5825 28135
rect 5859 28101 5871 28135
rect 5813 28095 5871 28101
rect 5276 28036 5488 28064
rect 5828 28064 5856 28095
rect 7006 28092 7012 28144
rect 7064 28092 7070 28144
rect 6730 28064 6736 28076
rect 5828 28036 6736 28064
rect 5169 28027 5227 28033
rect 5000 27996 5028 28027
rect 4724 27968 5028 27996
rect 4724 27937 4752 27968
rect 3200 27900 4476 27928
rect 4709 27931 4767 27937
rect 3200 27888 3206 27900
rect 4709 27897 4721 27931
rect 4755 27897 4767 27931
rect 5184 27928 5212 28027
rect 6730 28024 6736 28036
rect 6788 28024 6794 28076
rect 7300 28073 7328 28172
rect 7558 28160 7564 28172
rect 7616 28160 7622 28212
rect 8846 28200 8852 28212
rect 7668 28172 8852 28200
rect 7668 28132 7696 28172
rect 8846 28160 8852 28172
rect 8904 28160 8910 28212
rect 9582 28160 9588 28212
rect 9640 28200 9646 28212
rect 10413 28203 10471 28209
rect 10413 28200 10425 28203
rect 9640 28172 10425 28200
rect 9640 28160 9646 28172
rect 10413 28169 10425 28172
rect 10459 28169 10471 28203
rect 10413 28163 10471 28169
rect 15286 28160 15292 28212
rect 15344 28200 15350 28212
rect 15746 28200 15752 28212
rect 15344 28172 15752 28200
rect 15344 28160 15350 28172
rect 15746 28160 15752 28172
rect 15804 28200 15810 28212
rect 16025 28203 16083 28209
rect 16025 28200 16037 28203
rect 15804 28172 16037 28200
rect 15804 28160 15810 28172
rect 16025 28169 16037 28172
rect 16071 28169 16083 28203
rect 16025 28163 16083 28169
rect 17586 28160 17592 28212
rect 17644 28160 17650 28212
rect 17957 28203 18015 28209
rect 17957 28169 17969 28203
rect 18003 28200 18015 28203
rect 19058 28200 19064 28212
rect 18003 28172 19064 28200
rect 18003 28169 18015 28172
rect 17957 28163 18015 28169
rect 10226 28132 10232 28144
rect 7576 28104 7696 28132
rect 9062 28104 10232 28132
rect 7576 28073 7604 28104
rect 10226 28092 10232 28104
rect 10284 28092 10290 28144
rect 12618 28132 12624 28144
rect 12084 28104 12624 28132
rect 7285 28067 7343 28073
rect 7285 28033 7297 28067
rect 7331 28033 7343 28067
rect 7285 28027 7343 28033
rect 7561 28067 7619 28073
rect 7561 28033 7573 28067
rect 7607 28033 7619 28067
rect 7561 28027 7619 28033
rect 10410 28024 10416 28076
rect 10468 28024 10474 28076
rect 10502 28024 10508 28076
rect 10560 28064 10566 28076
rect 10597 28067 10655 28073
rect 10597 28064 10609 28067
rect 10560 28036 10609 28064
rect 10560 28024 10566 28036
rect 10597 28033 10609 28036
rect 10643 28033 10655 28067
rect 10597 28027 10655 28033
rect 11146 28024 11152 28076
rect 11204 28064 11210 28076
rect 12084 28073 12112 28104
rect 12618 28092 12624 28104
rect 12676 28092 12682 28144
rect 13630 28132 13636 28144
rect 13570 28104 13636 28132
rect 13630 28092 13636 28104
rect 13688 28132 13694 28144
rect 13688 28104 14306 28132
rect 13688 28092 13694 28104
rect 15194 28092 15200 28144
rect 15252 28132 15258 28144
rect 15252 28104 15792 28132
rect 15252 28092 15258 28104
rect 15764 28073 15792 28104
rect 16482 28092 16488 28144
rect 16540 28132 16546 28144
rect 17972 28132 18000 28163
rect 19058 28160 19064 28172
rect 19116 28160 19122 28212
rect 20257 28203 20315 28209
rect 20257 28169 20269 28203
rect 20303 28200 20315 28203
rect 20898 28200 20904 28212
rect 20303 28172 20904 28200
rect 20303 28169 20315 28172
rect 20257 28163 20315 28169
rect 20898 28160 20904 28172
rect 20956 28160 20962 28212
rect 21361 28203 21419 28209
rect 21361 28169 21373 28203
rect 21407 28200 21419 28203
rect 21818 28200 21824 28212
rect 21407 28172 21824 28200
rect 21407 28169 21419 28172
rect 21361 28163 21419 28169
rect 21818 28160 21824 28172
rect 21876 28160 21882 28212
rect 23934 28160 23940 28212
rect 23992 28160 23998 28212
rect 25961 28203 26019 28209
rect 25961 28169 25973 28203
rect 26007 28200 26019 28203
rect 28442 28200 28448 28212
rect 26007 28172 28448 28200
rect 26007 28169 26019 28172
rect 25961 28163 26019 28169
rect 28442 28160 28448 28172
rect 28500 28160 28506 28212
rect 29730 28160 29736 28212
rect 29788 28160 29794 28212
rect 30742 28160 30748 28212
rect 30800 28200 30806 28212
rect 31846 28200 31852 28212
rect 30800 28172 31852 28200
rect 30800 28160 30806 28172
rect 16540 28104 18000 28132
rect 16540 28092 16546 28104
rect 19334 28092 19340 28144
rect 19392 28132 19398 28144
rect 19705 28135 19763 28141
rect 19705 28132 19717 28135
rect 19392 28104 19717 28132
rect 19392 28092 19398 28104
rect 19705 28101 19717 28104
rect 19751 28101 19763 28135
rect 19705 28095 19763 28101
rect 20714 28092 20720 28144
rect 20772 28132 20778 28144
rect 22002 28132 22008 28144
rect 20772 28104 22008 28132
rect 20772 28092 20778 28104
rect 22002 28092 22008 28104
rect 22060 28092 22066 28144
rect 24210 28132 24216 28144
rect 22572 28104 24216 28132
rect 22572 28076 22600 28104
rect 24210 28092 24216 28104
rect 24268 28092 24274 28144
rect 26234 28132 26240 28144
rect 24596 28104 25452 28132
rect 24596 28076 24624 28104
rect 12069 28067 12127 28073
rect 12069 28064 12081 28067
rect 11204 28036 12081 28064
rect 11204 28024 11210 28036
rect 12069 28033 12081 28036
rect 12115 28033 12127 28067
rect 12069 28027 12127 28033
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28033 15899 28067
rect 15841 28027 15899 28033
rect 6914 27956 6920 28008
rect 6972 27956 6978 28008
rect 7101 27999 7159 28005
rect 7101 27965 7113 27999
rect 7147 27996 7159 27999
rect 7374 27996 7380 28008
rect 7147 27968 7380 27996
rect 7147 27965 7159 27968
rect 7101 27959 7159 27965
rect 7374 27956 7380 27968
rect 7432 27956 7438 28008
rect 7469 27999 7527 28005
rect 7469 27965 7481 27999
rect 7515 27996 7527 27999
rect 7837 27999 7895 28005
rect 7837 27996 7849 27999
rect 7515 27968 7849 27996
rect 7515 27965 7527 27968
rect 7469 27959 7527 27965
rect 7837 27965 7849 27968
rect 7883 27965 7895 27999
rect 7837 27959 7895 27965
rect 8202 27956 8208 28008
rect 8260 27996 8266 28008
rect 9309 27999 9367 28005
rect 9309 27996 9321 27999
rect 8260 27968 9321 27996
rect 8260 27956 8266 27968
rect 9309 27965 9321 27968
rect 9355 27965 9367 27999
rect 9309 27959 9367 27965
rect 12345 27999 12403 28005
rect 12345 27965 12357 27999
rect 12391 27996 12403 27999
rect 12986 27996 12992 28008
rect 12391 27968 12992 27996
rect 12391 27965 12403 27968
rect 12345 27959 12403 27965
rect 12986 27956 12992 27968
rect 13044 27956 13050 28008
rect 13814 27956 13820 28008
rect 13872 27996 13878 28008
rect 14001 27999 14059 28005
rect 14001 27996 14013 27999
rect 13872 27968 14013 27996
rect 13872 27956 13878 27968
rect 14001 27965 14013 27968
rect 14047 27965 14059 27999
rect 14001 27959 14059 27965
rect 6178 27928 6184 27940
rect 5184 27900 6184 27928
rect 4709 27891 4767 27897
rect 2866 27820 2872 27872
rect 2924 27860 2930 27872
rect 3697 27863 3755 27869
rect 3697 27860 3709 27863
rect 2924 27832 3709 27860
rect 2924 27820 2930 27832
rect 3697 27829 3709 27832
rect 3743 27829 3755 27863
rect 3697 27823 3755 27829
rect 3786 27820 3792 27872
rect 3844 27860 3850 27872
rect 5353 27863 5411 27869
rect 5353 27860 5365 27863
rect 3844 27832 5365 27860
rect 3844 27820 3850 27832
rect 5353 27829 5365 27832
rect 5399 27829 5411 27863
rect 5353 27823 5411 27829
rect 5442 27820 5448 27872
rect 5500 27820 5506 27872
rect 5644 27869 5672 27900
rect 6178 27888 6184 27900
rect 6236 27928 6242 27940
rect 6236 27900 7052 27928
rect 6236 27888 6242 27900
rect 5629 27863 5687 27869
rect 5629 27829 5641 27863
rect 5675 27829 5687 27863
rect 5629 27823 5687 27829
rect 6549 27863 6607 27869
rect 6549 27829 6561 27863
rect 6595 27860 6607 27863
rect 6914 27860 6920 27872
rect 6595 27832 6920 27860
rect 6595 27829 6607 27832
rect 6549 27823 6607 27829
rect 6914 27820 6920 27832
rect 6972 27820 6978 27872
rect 7024 27869 7052 27900
rect 7009 27863 7067 27869
rect 7009 27829 7021 27863
rect 7055 27829 7067 27863
rect 7009 27823 7067 27829
rect 13817 27863 13875 27869
rect 13817 27829 13829 27863
rect 13863 27860 13875 27863
rect 13906 27860 13912 27872
rect 13863 27832 13912 27860
rect 13863 27829 13875 27832
rect 13817 27823 13875 27829
rect 13906 27820 13912 27832
rect 13964 27820 13970 27872
rect 14016 27860 14044 27959
rect 15470 27956 15476 28008
rect 15528 27956 15534 28008
rect 15856 27860 15884 28027
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 17037 28067 17095 28073
rect 17037 28064 17049 28067
rect 15988 28036 17049 28064
rect 15988 28024 15994 28036
rect 17037 28033 17049 28036
rect 17083 28033 17095 28067
rect 17037 28027 17095 28033
rect 17129 28067 17187 28073
rect 17129 28033 17141 28067
rect 17175 28064 17187 28067
rect 17954 28064 17960 28076
rect 17175 28036 17960 28064
rect 17175 28033 17187 28036
rect 17129 28027 17187 28033
rect 17954 28024 17960 28036
rect 18012 28064 18018 28076
rect 18874 28064 18880 28076
rect 18012 28036 18880 28064
rect 18012 28024 18018 28036
rect 18874 28024 18880 28036
rect 18932 28024 18938 28076
rect 19518 28024 19524 28076
rect 19576 28024 19582 28076
rect 19981 28067 20039 28073
rect 19981 28064 19993 28067
rect 19904 28036 19993 28064
rect 16022 27956 16028 28008
rect 16080 27996 16086 28008
rect 17221 27999 17279 28005
rect 17221 27996 17233 27999
rect 16080 27968 17233 27996
rect 16080 27956 16086 27968
rect 17221 27965 17233 27968
rect 17267 27965 17279 27999
rect 17221 27959 17279 27965
rect 17236 27928 17264 27959
rect 18046 27956 18052 28008
rect 18104 27956 18110 28008
rect 18138 27956 18144 28008
rect 18196 27956 18202 28008
rect 18156 27928 18184 27956
rect 17236 27900 18184 27928
rect 14016 27832 15884 27860
rect 16669 27863 16727 27869
rect 16669 27829 16681 27863
rect 16715 27860 16727 27863
rect 16850 27860 16856 27872
rect 16715 27832 16856 27860
rect 16715 27829 16727 27832
rect 16669 27823 16727 27829
rect 16850 27820 16856 27832
rect 16908 27820 16914 27872
rect 19610 27820 19616 27872
rect 19668 27860 19674 27872
rect 19904 27869 19932 28036
rect 19981 28033 19993 28036
rect 20027 28033 20039 28067
rect 20993 28067 21051 28073
rect 20993 28064 21005 28067
rect 19981 28027 20039 28033
rect 20272 28036 21005 28064
rect 20272 28005 20300 28036
rect 20993 28033 21005 28036
rect 21039 28064 21051 28067
rect 21266 28064 21272 28076
rect 21039 28036 21272 28064
rect 21039 28033 21051 28036
rect 20993 28027 21051 28033
rect 21266 28024 21272 28036
rect 21324 28024 21330 28076
rect 22186 28024 22192 28076
rect 22244 28024 22250 28076
rect 22554 28024 22560 28076
rect 22612 28024 22618 28076
rect 22830 28073 22836 28076
rect 22824 28064 22836 28073
rect 22791 28036 22836 28064
rect 22824 28027 22836 28036
rect 22830 28024 22836 28027
rect 22888 28024 22894 28076
rect 24394 28024 24400 28076
rect 24452 28024 24458 28076
rect 24578 28024 24584 28076
rect 24636 28024 24642 28076
rect 24673 28067 24731 28073
rect 24673 28033 24685 28067
rect 24719 28064 24731 28067
rect 24854 28064 24860 28076
rect 24719 28036 24860 28064
rect 24719 28033 24731 28036
rect 24673 28027 24731 28033
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 24946 28024 24952 28076
rect 25004 28024 25010 28076
rect 25222 28024 25228 28076
rect 25280 28024 25286 28076
rect 25424 28073 25452 28104
rect 25516 28104 26240 28132
rect 25516 28073 25544 28104
rect 26234 28092 26240 28104
rect 26292 28092 26298 28144
rect 28258 28092 28264 28144
rect 28316 28092 28322 28144
rect 29270 28092 29276 28144
rect 29328 28092 29334 28144
rect 25409 28067 25467 28073
rect 25409 28033 25421 28067
rect 25455 28033 25467 28067
rect 25409 28027 25467 28033
rect 25501 28067 25559 28073
rect 25501 28033 25513 28067
rect 25547 28033 25559 28067
rect 25501 28027 25559 28033
rect 25682 28024 25688 28076
rect 25740 28064 25746 28076
rect 25777 28067 25835 28073
rect 25777 28064 25789 28067
rect 25740 28036 25789 28064
rect 25740 28024 25746 28036
rect 25777 28033 25789 28036
rect 25823 28064 25835 28067
rect 26053 28067 26111 28073
rect 26053 28064 26065 28067
rect 25823 28036 26065 28064
rect 25823 28033 25835 28036
rect 25777 28027 25835 28033
rect 26053 28033 26065 28036
rect 26099 28033 26111 28067
rect 26053 28027 26111 28033
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 27985 28067 28043 28073
rect 27985 28064 27997 28067
rect 27672 28036 27997 28064
rect 27672 28024 27678 28036
rect 27985 28033 27997 28036
rect 28031 28033 28043 28067
rect 27985 28027 28043 28033
rect 20257 27999 20315 28005
rect 20257 27965 20269 27999
rect 20303 27965 20315 27999
rect 20257 27959 20315 27965
rect 20714 27956 20720 28008
rect 20772 27996 20778 28008
rect 20901 27999 20959 28005
rect 20901 27996 20913 27999
rect 20772 27968 20913 27996
rect 20772 27956 20778 27968
rect 20901 27965 20913 27968
rect 20947 27965 20959 27999
rect 20901 27959 20959 27965
rect 21082 27956 21088 28008
rect 21140 27956 21146 28008
rect 21174 27956 21180 28008
rect 21232 27956 21238 28008
rect 24762 27956 24768 28008
rect 24820 27996 24826 28008
rect 25593 27999 25651 28005
rect 25593 27996 25605 27999
rect 24820 27968 25605 27996
rect 24820 27956 24826 27968
rect 25593 27965 25605 27968
rect 25639 27965 25651 27999
rect 25593 27959 25651 27965
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 26605 27999 26663 28005
rect 26605 27996 26617 27999
rect 26292 27968 26617 27996
rect 26292 27956 26298 27968
rect 26605 27965 26617 27968
rect 26651 27965 26663 27999
rect 26605 27959 26663 27965
rect 26970 27956 26976 28008
rect 27028 27956 27034 28008
rect 29288 27996 29316 28092
rect 29748 28064 29776 28160
rect 29914 28092 29920 28144
rect 29972 28132 29978 28144
rect 30193 28135 30251 28141
rect 30193 28132 30205 28135
rect 29972 28104 30205 28132
rect 29972 28092 29978 28104
rect 30193 28101 30205 28104
rect 30239 28101 30251 28135
rect 30193 28095 30251 28101
rect 31478 28092 31484 28144
rect 31536 28132 31542 28144
rect 31536 28104 31616 28132
rect 31536 28092 31542 28104
rect 30653 28067 30711 28073
rect 30653 28064 30665 28067
rect 29748 28036 30665 28064
rect 30653 28033 30665 28036
rect 30699 28064 30711 28067
rect 30742 28064 30748 28076
rect 30699 28036 30748 28064
rect 30699 28033 30711 28036
rect 30653 28027 30711 28033
rect 30742 28024 30748 28036
rect 30800 28024 30806 28076
rect 31588 28073 31616 28104
rect 31573 28067 31631 28073
rect 31573 28033 31585 28067
rect 31619 28033 31631 28067
rect 31680 28064 31708 28172
rect 31846 28160 31852 28172
rect 31904 28160 31910 28212
rect 34790 28160 34796 28212
rect 34848 28200 34854 28212
rect 36354 28200 36360 28212
rect 34848 28172 36360 28200
rect 34848 28160 34854 28172
rect 36354 28160 36360 28172
rect 36412 28160 36418 28212
rect 37734 28160 37740 28212
rect 37792 28200 37798 28212
rect 37921 28203 37979 28209
rect 37921 28200 37933 28203
rect 37792 28172 37933 28200
rect 37792 28160 37798 28172
rect 37921 28169 37933 28172
rect 37967 28169 37979 28203
rect 37921 28163 37979 28169
rect 32950 28092 32956 28144
rect 33008 28092 33014 28144
rect 33686 28092 33692 28144
rect 33744 28132 33750 28144
rect 33744 28104 34560 28132
rect 33744 28092 33750 28104
rect 31757 28067 31815 28073
rect 31757 28064 31769 28067
rect 31680 28036 31769 28064
rect 31573 28027 31631 28033
rect 31757 28033 31769 28036
rect 31803 28033 31815 28067
rect 31757 28027 31815 28033
rect 34330 28024 34336 28076
rect 34388 28024 34394 28076
rect 34532 28073 34560 28104
rect 37550 28092 37556 28144
rect 37608 28092 37614 28144
rect 37642 28092 37648 28144
rect 37700 28092 37706 28144
rect 34517 28067 34575 28073
rect 34517 28033 34529 28067
rect 34563 28033 34575 28067
rect 34517 28027 34575 28033
rect 37274 28024 37280 28076
rect 37332 28024 37338 28076
rect 37425 28067 37483 28073
rect 37425 28033 37437 28067
rect 37471 28064 37483 28067
rect 37471 28036 37596 28064
rect 37471 28033 37483 28036
rect 37425 28027 37483 28033
rect 29917 27999 29975 28005
rect 29917 27996 29929 27999
rect 29288 27968 29929 27996
rect 29917 27965 29929 27968
rect 29963 27965 29975 27999
rect 29917 27959 29975 27965
rect 30834 27956 30840 28008
rect 30892 27956 30898 28008
rect 30929 27999 30987 28005
rect 30929 27965 30941 27999
rect 30975 27996 30987 27999
rect 31110 27996 31116 28008
rect 30975 27968 31116 27996
rect 30975 27965 30987 27968
rect 30929 27959 30987 27965
rect 31110 27956 31116 27968
rect 31168 27956 31174 28008
rect 31481 27999 31539 28005
rect 31481 27965 31493 27999
rect 31527 27965 31539 27999
rect 31481 27959 31539 27965
rect 32217 27999 32275 28005
rect 32217 27965 32229 27999
rect 32263 27996 32275 27999
rect 32766 27996 32772 28008
rect 32263 27968 32772 27996
rect 32263 27965 32275 27968
rect 32217 27959 32275 27965
rect 25133 27931 25191 27937
rect 25133 27897 25145 27931
rect 25179 27928 25191 27931
rect 26326 27928 26332 27940
rect 25179 27900 26332 27928
rect 25179 27897 25191 27900
rect 25133 27891 25191 27897
rect 26326 27888 26332 27900
rect 26384 27888 26390 27940
rect 30745 27931 30803 27937
rect 30745 27897 30757 27931
rect 30791 27928 30803 27931
rect 30852 27928 30880 27956
rect 31496 27928 31524 27959
rect 32766 27956 32772 27968
rect 32824 27956 32830 28008
rect 33962 27956 33968 28008
rect 34020 27956 34026 28008
rect 34241 27999 34299 28005
rect 34241 27965 34253 27999
rect 34287 27996 34299 27999
rect 35434 27996 35440 28008
rect 34287 27968 35440 27996
rect 34287 27965 34299 27968
rect 34241 27959 34299 27965
rect 35434 27956 35440 27968
rect 35492 27956 35498 28008
rect 35250 27928 35256 27940
rect 30791 27900 31524 27928
rect 34440 27900 35256 27928
rect 30791 27897 30803 27900
rect 30745 27891 30803 27897
rect 19889 27863 19947 27869
rect 19889 27860 19901 27863
rect 19668 27832 19901 27860
rect 19668 27820 19674 27832
rect 19889 27829 19901 27832
rect 19935 27829 19947 27863
rect 19889 27823 19947 27829
rect 20070 27820 20076 27872
rect 20128 27820 20134 27872
rect 21542 27820 21548 27872
rect 21600 27860 21606 27872
rect 21821 27863 21879 27869
rect 21821 27860 21833 27863
rect 21600 27832 21833 27860
rect 21600 27820 21606 27832
rect 21821 27829 21833 27832
rect 21867 27829 21879 27863
rect 21821 27823 21879 27829
rect 27522 27820 27528 27872
rect 27580 27860 27586 27872
rect 27617 27863 27675 27869
rect 27617 27860 27629 27863
rect 27580 27832 27629 27860
rect 27580 27820 27586 27832
rect 27617 27829 27629 27832
rect 27663 27829 27675 27863
rect 27617 27823 27675 27829
rect 30837 27863 30895 27869
rect 30837 27829 30849 27863
rect 30883 27860 30895 27863
rect 31478 27860 31484 27872
rect 30883 27832 31484 27860
rect 30883 27829 30895 27832
rect 30837 27823 30895 27829
rect 31478 27820 31484 27832
rect 31536 27820 31542 27872
rect 31941 27863 31999 27869
rect 31941 27829 31953 27863
rect 31987 27860 31999 27863
rect 32674 27860 32680 27872
rect 31987 27832 32680 27860
rect 31987 27829 31999 27832
rect 31941 27823 31999 27829
rect 32674 27820 32680 27832
rect 32732 27860 32738 27872
rect 34440 27860 34468 27900
rect 35250 27888 35256 27900
rect 35308 27888 35314 27940
rect 37568 27928 37596 28036
rect 37734 28024 37740 28076
rect 37792 28073 37798 28076
rect 37792 28027 37800 28073
rect 37792 28024 37798 28027
rect 38010 28024 38016 28076
rect 38068 28024 38074 28076
rect 38010 27928 38016 27940
rect 37568 27900 38016 27928
rect 38010 27888 38016 27900
rect 38068 27888 38074 27940
rect 32732 27832 34468 27860
rect 32732 27820 32738 27832
rect 34514 27820 34520 27872
rect 34572 27820 34578 27872
rect 38194 27820 38200 27872
rect 38252 27820 38258 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 3418 27616 3424 27668
rect 3476 27616 3482 27668
rect 3602 27616 3608 27668
rect 3660 27616 3666 27668
rect 3970 27616 3976 27668
rect 4028 27616 4034 27668
rect 7377 27659 7435 27665
rect 7377 27625 7389 27659
rect 7423 27656 7435 27659
rect 7558 27656 7564 27668
rect 7423 27628 7564 27656
rect 7423 27625 7435 27628
rect 7377 27619 7435 27625
rect 7558 27616 7564 27628
rect 7616 27616 7622 27668
rect 11320 27659 11378 27665
rect 11320 27625 11332 27659
rect 11366 27656 11378 27659
rect 11366 27628 13032 27656
rect 11366 27625 11378 27628
rect 11320 27619 11378 27625
rect 4249 27591 4307 27597
rect 4249 27557 4261 27591
rect 4295 27588 4307 27591
rect 7282 27588 7288 27600
rect 4295 27560 7288 27588
rect 4295 27557 4307 27560
rect 4249 27551 4307 27557
rect 7282 27548 7288 27560
rect 7340 27548 7346 27600
rect 13004 27597 13032 27628
rect 13906 27616 13912 27668
rect 13964 27656 13970 27668
rect 14366 27656 14372 27668
rect 13964 27628 14372 27656
rect 13964 27616 13970 27628
rect 14366 27616 14372 27628
rect 14424 27616 14430 27668
rect 16390 27656 16396 27668
rect 15948 27628 16396 27656
rect 12989 27591 13047 27597
rect 12989 27557 13001 27591
rect 13035 27557 13047 27591
rect 12989 27551 13047 27557
rect 14550 27548 14556 27600
rect 14608 27588 14614 27600
rect 15102 27588 15108 27600
rect 14608 27560 15108 27588
rect 14608 27548 14614 27560
rect 15102 27548 15108 27560
rect 15160 27588 15166 27600
rect 15948 27588 15976 27628
rect 16390 27616 16396 27628
rect 16448 27616 16454 27668
rect 16850 27616 16856 27668
rect 16908 27656 16914 27668
rect 16957 27659 17015 27665
rect 16957 27656 16969 27659
rect 16908 27628 16969 27656
rect 16908 27616 16914 27628
rect 16957 27625 16969 27628
rect 17003 27625 17015 27659
rect 16957 27619 17015 27625
rect 17770 27616 17776 27668
rect 17828 27656 17834 27668
rect 18782 27656 18788 27668
rect 17828 27628 18788 27656
rect 17828 27616 17834 27628
rect 15160 27560 15976 27588
rect 15160 27548 15166 27560
rect 17586 27548 17592 27600
rect 17644 27548 17650 27600
rect 3326 27480 3332 27532
rect 3384 27520 3390 27532
rect 3881 27523 3939 27529
rect 3881 27520 3893 27523
rect 3384 27492 3893 27520
rect 3384 27480 3390 27492
rect 3881 27489 3893 27492
rect 3927 27489 3939 27523
rect 3881 27483 3939 27489
rect 13538 27480 13544 27532
rect 13596 27480 13602 27532
rect 15286 27520 15292 27532
rect 14292 27492 15292 27520
rect 1394 27412 1400 27464
rect 1452 27412 1458 27464
rect 2774 27412 2780 27464
rect 2832 27452 2838 27464
rect 3050 27452 3056 27464
rect 2832 27424 3056 27452
rect 2832 27412 2838 27424
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 3142 27412 3148 27464
rect 3200 27452 3206 27464
rect 3200 27424 3372 27452
rect 3200 27412 3206 27424
rect 1670 27344 1676 27396
rect 1728 27344 1734 27396
rect 3237 27387 3295 27393
rect 3237 27353 3249 27387
rect 3283 27353 3295 27387
rect 3344 27384 3372 27424
rect 3602 27412 3608 27464
rect 3660 27452 3666 27464
rect 3789 27455 3847 27461
rect 3789 27452 3801 27455
rect 3660 27424 3801 27452
rect 3660 27412 3666 27424
rect 3789 27421 3801 27424
rect 3835 27421 3847 27455
rect 3789 27415 3847 27421
rect 4065 27455 4123 27461
rect 4065 27421 4077 27455
rect 4111 27452 4123 27455
rect 4614 27452 4620 27464
rect 4111 27424 4620 27452
rect 4111 27421 4123 27424
rect 4065 27415 4123 27421
rect 3437 27387 3495 27393
rect 3437 27384 3449 27387
rect 3344 27356 3449 27384
rect 3237 27347 3295 27353
rect 3437 27353 3449 27356
rect 3483 27353 3495 27387
rect 3437 27347 3495 27353
rect 3145 27319 3203 27325
rect 3145 27285 3157 27319
rect 3191 27316 3203 27319
rect 3252 27316 3280 27347
rect 3326 27316 3332 27328
rect 3191 27288 3332 27316
rect 3191 27285 3203 27288
rect 3145 27279 3203 27285
rect 3326 27276 3332 27288
rect 3384 27316 3390 27328
rect 4080 27316 4108 27415
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 7006 27412 7012 27464
rect 7064 27452 7070 27464
rect 7285 27455 7343 27461
rect 7285 27452 7297 27455
rect 7064 27424 7297 27452
rect 7064 27412 7070 27424
rect 7285 27421 7297 27424
rect 7331 27421 7343 27455
rect 7285 27415 7343 27421
rect 7466 27412 7472 27464
rect 7524 27412 7530 27464
rect 10226 27412 10232 27464
rect 10284 27452 10290 27464
rect 14292 27461 14320 27492
rect 15286 27480 15292 27492
rect 15344 27480 15350 27532
rect 15654 27520 15660 27532
rect 15396 27492 15660 27520
rect 11057 27455 11115 27461
rect 11057 27452 11069 27455
rect 10284 27424 11069 27452
rect 10284 27412 10290 27424
rect 11057 27421 11069 27424
rect 11103 27421 11115 27455
rect 11057 27415 11115 27421
rect 14277 27455 14335 27461
rect 14277 27421 14289 27455
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27452 14703 27455
rect 14691 27424 15148 27452
rect 14691 27421 14703 27424
rect 14645 27415 14703 27421
rect 4341 27387 4399 27393
rect 4341 27353 4353 27387
rect 4387 27353 4399 27387
rect 4341 27347 4399 27353
rect 5169 27387 5227 27393
rect 5169 27353 5181 27387
rect 5215 27384 5227 27387
rect 5258 27384 5264 27396
rect 5215 27356 5264 27384
rect 5215 27353 5227 27356
rect 5169 27347 5227 27353
rect 3384 27288 4108 27316
rect 4356 27316 4384 27347
rect 5258 27344 5264 27356
rect 5316 27344 5322 27396
rect 12618 27384 12624 27396
rect 12558 27356 12624 27384
rect 12618 27344 12624 27356
rect 12676 27384 12682 27396
rect 13630 27384 13636 27396
rect 12676 27356 13636 27384
rect 12676 27344 12682 27356
rect 13630 27344 13636 27356
rect 13688 27344 13694 27396
rect 5442 27316 5448 27328
rect 4356 27288 5448 27316
rect 3384 27276 3390 27288
rect 5442 27276 5448 27288
rect 5500 27316 5506 27328
rect 6362 27316 6368 27328
rect 5500 27288 6368 27316
rect 5500 27276 5506 27288
rect 6362 27276 6368 27288
rect 6420 27276 6426 27328
rect 12805 27319 12863 27325
rect 12805 27285 12817 27319
rect 12851 27316 12863 27319
rect 13078 27316 13084 27328
rect 12851 27288 13084 27316
rect 12851 27285 12863 27288
rect 12805 27279 12863 27285
rect 13078 27276 13084 27288
rect 13136 27316 13142 27328
rect 13357 27319 13415 27325
rect 13357 27316 13369 27319
rect 13136 27288 13369 27316
rect 13136 27276 13142 27288
rect 13357 27285 13369 27288
rect 13403 27285 13415 27319
rect 13357 27279 13415 27285
rect 13446 27276 13452 27328
rect 13504 27276 13510 27328
rect 14826 27276 14832 27328
rect 14884 27276 14890 27328
rect 15120 27316 15148 27424
rect 15194 27412 15200 27464
rect 15252 27452 15258 27464
rect 15396 27452 15424 27492
rect 15654 27480 15660 27492
rect 15712 27520 15718 27532
rect 15930 27520 15936 27532
rect 15712 27492 15936 27520
rect 15712 27480 15718 27492
rect 15930 27480 15936 27492
rect 15988 27480 15994 27532
rect 16942 27480 16948 27532
rect 17000 27520 17006 27532
rect 17221 27523 17279 27529
rect 17221 27520 17233 27523
rect 17000 27492 17233 27520
rect 17000 27480 17006 27492
rect 17221 27489 17233 27492
rect 17267 27489 17279 27523
rect 17221 27483 17279 27489
rect 17605 27461 17633 27548
rect 18248 27471 18276 27628
rect 18782 27616 18788 27628
rect 18840 27656 18846 27668
rect 18840 27628 19334 27656
rect 18840 27616 18846 27628
rect 19306 27600 19334 27628
rect 19518 27616 19524 27668
rect 19576 27656 19582 27668
rect 20073 27659 20131 27665
rect 20073 27656 20085 27659
rect 19576 27628 20085 27656
rect 19576 27616 19582 27628
rect 20073 27625 20085 27628
rect 20119 27625 20131 27659
rect 22830 27656 22836 27668
rect 20073 27619 20131 27625
rect 22066 27628 22836 27656
rect 19306 27560 19340 27600
rect 19334 27548 19340 27560
rect 19392 27548 19398 27600
rect 19426 27548 19432 27600
rect 19484 27588 19490 27600
rect 20441 27591 20499 27597
rect 19484 27560 20300 27588
rect 19484 27548 19490 27560
rect 19058 27480 19064 27532
rect 19116 27520 19122 27532
rect 19705 27523 19763 27529
rect 19705 27520 19717 27523
rect 19116 27492 19717 27520
rect 19116 27480 19122 27492
rect 19705 27489 19717 27492
rect 19751 27489 19763 27523
rect 19705 27483 19763 27489
rect 18233 27465 18291 27471
rect 17486 27455 17544 27461
rect 17486 27452 17498 27455
rect 15252 27424 15424 27452
rect 15252 27412 15258 27424
rect 17482 27421 17498 27452
rect 17532 27421 17544 27455
rect 17482 27415 17544 27421
rect 17590 27455 17648 27461
rect 17590 27421 17602 27455
rect 17636 27421 17648 27455
rect 17590 27415 17648 27421
rect 16390 27344 16396 27396
rect 16448 27344 16454 27396
rect 17482 27384 17510 27415
rect 17678 27412 17684 27464
rect 17736 27452 17742 27464
rect 18049 27455 18107 27461
rect 18049 27452 18061 27455
rect 17736 27424 18061 27452
rect 17736 27412 17742 27424
rect 18049 27421 18061 27424
rect 18095 27421 18107 27455
rect 18233 27431 18245 27465
rect 18279 27431 18291 27465
rect 18233 27425 18291 27431
rect 18417 27455 18475 27461
rect 18049 27415 18107 27421
rect 18417 27421 18429 27455
rect 18463 27452 18475 27455
rect 18966 27452 18972 27464
rect 18463 27424 18972 27452
rect 18463 27421 18475 27424
rect 18417 27415 18475 27421
rect 17954 27384 17960 27396
rect 17482 27356 17960 27384
rect 17954 27344 17960 27356
rect 18012 27344 18018 27396
rect 18064 27384 18092 27415
rect 18432 27384 18460 27415
rect 18966 27412 18972 27424
rect 19024 27412 19030 27464
rect 19334 27412 19340 27464
rect 19392 27412 19398 27464
rect 19518 27412 19524 27464
rect 19576 27412 19582 27464
rect 20272 27461 20300 27560
rect 20441 27557 20453 27591
rect 20487 27588 20499 27591
rect 21174 27588 21180 27600
rect 20487 27560 21180 27588
rect 20487 27557 20499 27560
rect 20441 27551 20499 27557
rect 21174 27548 21180 27560
rect 21232 27548 21238 27600
rect 22066 27588 22094 27628
rect 22830 27616 22836 27628
rect 22888 27616 22894 27668
rect 27359 27659 27417 27665
rect 27359 27625 27371 27659
rect 27405 27656 27417 27659
rect 27522 27656 27528 27668
rect 27405 27628 27528 27656
rect 27405 27625 27417 27628
rect 27359 27619 27417 27625
rect 27522 27616 27528 27628
rect 27580 27616 27586 27668
rect 27706 27616 27712 27668
rect 27764 27656 27770 27668
rect 28169 27659 28227 27665
rect 28169 27656 28181 27659
rect 27764 27628 28181 27656
rect 27764 27616 27770 27628
rect 28169 27625 28181 27628
rect 28215 27656 28227 27659
rect 28718 27656 28724 27668
rect 28215 27628 28724 27656
rect 28215 27625 28227 27628
rect 28169 27619 28227 27625
rect 28718 27616 28724 27628
rect 28776 27616 28782 27668
rect 28813 27659 28871 27665
rect 28813 27625 28825 27659
rect 28859 27656 28871 27659
rect 29822 27656 29828 27668
rect 28859 27628 29828 27656
rect 28859 27625 28871 27628
rect 28813 27619 28871 27625
rect 29822 27616 29828 27628
rect 29880 27616 29886 27668
rect 31297 27659 31355 27665
rect 31297 27625 31309 27659
rect 31343 27656 31355 27659
rect 31386 27656 31392 27668
rect 31343 27628 31392 27656
rect 31343 27625 31355 27628
rect 31297 27619 31355 27625
rect 31386 27616 31392 27628
rect 31444 27616 31450 27668
rect 31754 27616 31760 27668
rect 31812 27616 31818 27668
rect 33229 27659 33287 27665
rect 33229 27625 33241 27659
rect 33275 27656 33287 27659
rect 33962 27656 33968 27668
rect 33275 27628 33968 27656
rect 33275 27625 33287 27628
rect 33229 27619 33287 27625
rect 33962 27616 33968 27628
rect 34020 27616 34026 27668
rect 37734 27656 37740 27668
rect 37476 27628 37740 27656
rect 24762 27588 24768 27600
rect 21284 27560 22094 27588
rect 23952 27560 24768 27588
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27421 19671 27455
rect 19797 27455 19855 27461
rect 19797 27452 19809 27455
rect 19613 27415 19671 27421
rect 19720 27424 19809 27452
rect 18064 27356 18460 27384
rect 18690 27344 18696 27396
rect 18748 27344 18754 27396
rect 18874 27344 18880 27396
rect 18932 27384 18938 27396
rect 19426 27384 19432 27396
rect 18932 27356 19432 27384
rect 18932 27344 18938 27356
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 16298 27316 16304 27328
rect 15120 27288 16304 27316
rect 16298 27276 16304 27288
rect 16356 27276 16362 27328
rect 17862 27276 17868 27328
rect 17920 27276 17926 27328
rect 18138 27276 18144 27328
rect 18196 27276 18202 27328
rect 18414 27276 18420 27328
rect 18472 27316 18478 27328
rect 18509 27319 18567 27325
rect 18509 27316 18521 27319
rect 18472 27288 18521 27316
rect 18472 27276 18478 27288
rect 18509 27285 18521 27288
rect 18555 27285 18567 27319
rect 18509 27279 18567 27285
rect 19061 27319 19119 27325
rect 19061 27285 19073 27319
rect 19107 27316 19119 27319
rect 19628 27316 19656 27415
rect 19720 27396 19748 27424
rect 19797 27421 19809 27424
rect 19843 27452 19855 27455
rect 20073 27455 20131 27461
rect 20073 27452 20085 27455
rect 19843 27424 20085 27452
rect 19843 27421 19855 27424
rect 19797 27415 19855 27421
rect 20073 27421 20085 27424
rect 20119 27421 20131 27455
rect 20073 27415 20131 27421
rect 20257 27455 20315 27461
rect 20257 27421 20269 27455
rect 20303 27452 20315 27455
rect 20438 27452 20444 27464
rect 20303 27424 20444 27452
rect 20303 27421 20315 27424
rect 20257 27415 20315 27421
rect 20438 27412 20444 27424
rect 20496 27412 20502 27464
rect 21284 27461 21312 27560
rect 21542 27480 21548 27532
rect 21600 27480 21606 27532
rect 21269 27455 21327 27461
rect 21269 27421 21281 27455
rect 21315 27421 21327 27455
rect 21269 27415 21327 27421
rect 21450 27412 21456 27464
rect 21508 27412 21514 27464
rect 21637 27455 21695 27461
rect 21637 27421 21649 27455
rect 21683 27421 21695 27455
rect 21637 27415 21695 27421
rect 19702 27344 19708 27396
rect 19760 27344 19766 27396
rect 20809 27387 20867 27393
rect 20809 27384 20821 27387
rect 19996 27356 20821 27384
rect 19794 27316 19800 27328
rect 19107 27288 19800 27316
rect 19107 27285 19119 27288
rect 19061 27279 19119 27285
rect 19794 27276 19800 27288
rect 19852 27276 19858 27328
rect 19996 27325 20024 27356
rect 20809 27353 20821 27356
rect 20855 27353 20867 27387
rect 20809 27347 20867 27353
rect 20901 27387 20959 27393
rect 20901 27353 20913 27387
rect 20947 27384 20959 27387
rect 21082 27384 21088 27396
rect 20947 27356 21088 27384
rect 20947 27353 20959 27356
rect 20901 27347 20959 27353
rect 21082 27344 21088 27356
rect 21140 27344 21146 27396
rect 21177 27387 21235 27393
rect 21177 27353 21189 27387
rect 21223 27384 21235 27387
rect 21542 27384 21548 27396
rect 21223 27356 21548 27384
rect 21223 27353 21235 27356
rect 21177 27347 21235 27353
rect 21542 27344 21548 27356
rect 21600 27344 21606 27396
rect 19981 27319 20039 27325
rect 19981 27285 19993 27319
rect 20027 27285 20039 27319
rect 19981 27279 20039 27285
rect 20622 27276 20628 27328
rect 20680 27276 20686 27328
rect 20993 27319 21051 27325
rect 20993 27285 21005 27319
rect 21039 27316 21051 27319
rect 21358 27316 21364 27328
rect 21039 27288 21364 27316
rect 21039 27285 21051 27288
rect 20993 27279 21051 27285
rect 21358 27276 21364 27288
rect 21416 27276 21422 27328
rect 21652 27316 21680 27415
rect 21818 27412 21824 27464
rect 21876 27412 21882 27464
rect 22097 27455 22155 27461
rect 22097 27421 22109 27455
rect 22143 27452 22155 27455
rect 22922 27452 22928 27464
rect 22143 27424 22928 27452
rect 22143 27421 22155 27424
rect 22097 27415 22155 27421
rect 22922 27412 22928 27424
rect 22980 27412 22986 27464
rect 23952 27461 23980 27560
rect 24762 27548 24768 27560
rect 24820 27548 24826 27600
rect 25869 27591 25927 27597
rect 25869 27557 25881 27591
rect 25915 27588 25927 27591
rect 26234 27588 26240 27600
rect 25915 27560 26240 27588
rect 25915 27557 25927 27560
rect 25869 27551 25927 27557
rect 26234 27548 26240 27560
rect 26292 27548 26298 27600
rect 28537 27591 28595 27597
rect 28537 27557 28549 27591
rect 28583 27588 28595 27591
rect 28629 27591 28687 27597
rect 28629 27588 28641 27591
rect 28583 27560 28641 27588
rect 28583 27557 28595 27560
rect 28537 27551 28595 27557
rect 28629 27557 28641 27560
rect 28675 27588 28687 27591
rect 28994 27588 29000 27600
rect 28675 27560 29000 27588
rect 28675 27557 28687 27560
rect 28629 27551 28687 27557
rect 28994 27548 29000 27560
rect 29052 27548 29058 27600
rect 31404 27588 31432 27616
rect 31404 27560 31800 27588
rect 24213 27523 24271 27529
rect 24213 27489 24225 27523
rect 24259 27520 24271 27523
rect 24578 27520 24584 27532
rect 24259 27492 24584 27520
rect 24259 27489 24271 27492
rect 24213 27483 24271 27489
rect 24578 27480 24584 27492
rect 24636 27520 24642 27532
rect 25317 27523 25375 27529
rect 24636 27492 25268 27520
rect 24636 27480 24642 27492
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 24026 27412 24032 27464
rect 24084 27452 24090 27464
rect 25240 27461 25268 27492
rect 25317 27489 25329 27523
rect 25363 27520 25375 27523
rect 25682 27520 25688 27532
rect 25363 27492 25688 27520
rect 25363 27489 25375 27492
rect 25317 27483 25375 27489
rect 25682 27480 25688 27492
rect 25740 27480 25746 27532
rect 25777 27523 25835 27529
rect 25777 27489 25789 27523
rect 25823 27520 25835 27523
rect 26970 27520 26976 27532
rect 25823 27492 26976 27520
rect 25823 27489 25835 27492
rect 25777 27483 25835 27489
rect 26970 27480 26976 27492
rect 27028 27480 27034 27532
rect 27614 27480 27620 27532
rect 27672 27480 27678 27532
rect 30834 27480 30840 27532
rect 30892 27480 30898 27532
rect 31110 27480 31116 27532
rect 31168 27480 31174 27532
rect 24121 27455 24179 27461
rect 24121 27452 24133 27455
rect 24084 27424 24133 27452
rect 24084 27412 24090 27424
rect 24121 27421 24133 27424
rect 24167 27421 24179 27455
rect 24121 27415 24179 27421
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27452 24823 27455
rect 25041 27455 25099 27461
rect 25041 27452 25053 27455
rect 24811 27424 25053 27452
rect 24811 27421 24823 27424
rect 24765 27415 24823 27421
rect 25041 27421 25053 27424
rect 25087 27421 25099 27455
rect 25041 27415 25099 27421
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 25593 27455 25651 27461
rect 25593 27421 25605 27455
rect 25639 27452 25651 27455
rect 25866 27452 25872 27464
rect 25639 27424 25872 27452
rect 25639 27421 25651 27424
rect 25593 27415 25651 27421
rect 22005 27387 22063 27393
rect 22005 27353 22017 27387
rect 22051 27384 22063 27387
rect 22342 27387 22400 27393
rect 22342 27384 22354 27387
rect 22051 27356 22354 27384
rect 22051 27353 22063 27356
rect 22005 27347 22063 27353
rect 22342 27353 22354 27356
rect 22388 27353 22400 27387
rect 24136 27384 24164 27415
rect 24302 27384 24308 27396
rect 24136 27356 24308 27384
rect 22342 27347 22400 27353
rect 24302 27344 24308 27356
rect 24360 27384 24366 27396
rect 24397 27387 24455 27393
rect 24397 27384 24409 27387
rect 24360 27356 24409 27384
rect 24360 27344 24366 27356
rect 24397 27353 24409 27356
rect 24443 27353 24455 27387
rect 24397 27347 24455 27353
rect 24581 27387 24639 27393
rect 24581 27353 24593 27387
rect 24627 27353 24639 27387
rect 24581 27347 24639 27353
rect 22738 27316 22744 27328
rect 21652 27288 22744 27316
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 23290 27276 23296 27328
rect 23348 27316 23354 27328
rect 23477 27319 23535 27325
rect 23477 27316 23489 27319
rect 23348 27288 23489 27316
rect 23348 27276 23354 27288
rect 23477 27285 23489 27288
rect 23523 27316 23535 27319
rect 24596 27316 24624 27347
rect 24854 27344 24860 27396
rect 24912 27384 24918 27396
rect 25424 27384 25452 27415
rect 25866 27412 25872 27424
rect 25924 27412 25930 27464
rect 30742 27412 30748 27464
rect 30800 27412 30806 27464
rect 30852 27452 30880 27480
rect 31205 27455 31263 27461
rect 31205 27452 31217 27455
rect 30852 27424 31217 27452
rect 31205 27421 31217 27424
rect 31251 27421 31263 27455
rect 31205 27415 31263 27421
rect 31478 27412 31484 27464
rect 31536 27412 31542 27464
rect 31772 27461 31800 27560
rect 32122 27548 32128 27600
rect 32180 27548 32186 27600
rect 32861 27591 32919 27597
rect 32861 27557 32873 27591
rect 32907 27588 32919 27591
rect 33134 27588 33140 27600
rect 32907 27560 33140 27588
rect 32907 27557 32919 27560
rect 32861 27551 32919 27557
rect 33134 27548 33140 27560
rect 33192 27548 33198 27600
rect 35342 27548 35348 27600
rect 35400 27548 35406 27600
rect 37093 27591 37151 27597
rect 37093 27557 37105 27591
rect 37139 27588 37151 27591
rect 37476 27588 37504 27628
rect 37734 27616 37740 27628
rect 37792 27616 37798 27668
rect 37918 27616 37924 27668
rect 37976 27656 37982 27668
rect 38381 27659 38439 27665
rect 38381 27656 38393 27659
rect 37976 27628 38393 27656
rect 37976 27616 37982 27628
rect 38381 27625 38393 27628
rect 38427 27625 38439 27659
rect 38381 27619 38439 27625
rect 37139 27560 37504 27588
rect 37139 27557 37151 27560
rect 37093 27551 37151 27557
rect 37550 27548 37556 27600
rect 37608 27548 37614 27600
rect 31846 27480 31852 27532
rect 31904 27480 31910 27532
rect 32766 27480 32772 27532
rect 32824 27480 32830 27532
rect 35360 27520 35388 27548
rect 37568 27520 37596 27548
rect 35360 27492 36952 27520
rect 37568 27492 38148 27520
rect 31757 27455 31815 27461
rect 31757 27421 31769 27455
rect 31803 27421 31815 27455
rect 31757 27415 31815 27421
rect 33042 27412 33048 27464
rect 33100 27412 33106 27464
rect 35161 27455 35219 27461
rect 35161 27421 35173 27455
rect 35207 27421 35219 27455
rect 35161 27415 35219 27421
rect 24912 27356 25452 27384
rect 24912 27344 24918 27356
rect 23523 27288 24624 27316
rect 25424 27316 25452 27356
rect 26878 27344 26884 27396
rect 26936 27344 26942 27396
rect 28258 27344 28264 27396
rect 28316 27384 28322 27396
rect 28997 27387 29055 27393
rect 28997 27384 29009 27387
rect 28316 27356 29009 27384
rect 28316 27344 28322 27356
rect 28997 27353 29009 27356
rect 29043 27353 29055 27387
rect 28997 27347 29055 27353
rect 31665 27387 31723 27393
rect 31665 27353 31677 27387
rect 31711 27384 31723 27387
rect 32398 27384 32404 27396
rect 31711 27356 32404 27384
rect 31711 27353 31723 27356
rect 31665 27347 31723 27353
rect 32398 27344 32404 27356
rect 32456 27344 32462 27396
rect 35176 27384 35204 27415
rect 35250 27412 35256 27464
rect 35308 27452 35314 27464
rect 35345 27455 35403 27461
rect 35345 27452 35357 27455
rect 35308 27424 35357 27452
rect 35308 27412 35314 27424
rect 35345 27421 35357 27424
rect 35391 27421 35403 27455
rect 35345 27415 35403 27421
rect 35176 27356 35388 27384
rect 35360 27328 35388 27356
rect 26418 27316 26424 27328
rect 25424 27288 26424 27316
rect 23523 27285 23535 27288
rect 23477 27279 23535 27285
rect 26418 27276 26424 27288
rect 26476 27276 26482 27328
rect 27982 27276 27988 27328
rect 28040 27276 28046 27328
rect 28166 27276 28172 27328
rect 28224 27276 28230 27328
rect 28810 27325 28816 27328
rect 28797 27319 28816 27325
rect 28797 27285 28809 27319
rect 28797 27279 28816 27285
rect 28810 27276 28816 27279
rect 28868 27276 28874 27328
rect 29638 27276 29644 27328
rect 29696 27316 29702 27328
rect 32950 27316 32956 27328
rect 29696 27288 32956 27316
rect 29696 27276 29702 27288
rect 32950 27276 32956 27288
rect 33008 27276 33014 27328
rect 34790 27276 34796 27328
rect 34848 27316 34854 27328
rect 35253 27319 35311 27325
rect 35253 27316 35265 27319
rect 34848 27288 35265 27316
rect 34848 27276 34854 27288
rect 35253 27285 35265 27288
rect 35299 27285 35311 27319
rect 35253 27279 35311 27285
rect 35342 27276 35348 27328
rect 35400 27276 35406 27328
rect 36924 27316 36952 27492
rect 37001 27455 37059 27461
rect 37001 27421 37013 27455
rect 37047 27452 37059 27455
rect 37366 27452 37372 27464
rect 37047 27424 37372 27452
rect 37047 27421 37059 27424
rect 37001 27415 37059 27421
rect 37366 27412 37372 27424
rect 37424 27412 37430 27464
rect 37520 27455 37578 27461
rect 37520 27421 37532 27455
rect 37566 27452 37578 27455
rect 37737 27455 37795 27461
rect 37737 27452 37749 27455
rect 37566 27421 37596 27452
rect 37520 27415 37596 27421
rect 37568 27328 37596 27415
rect 37660 27424 37749 27452
rect 37458 27316 37464 27328
rect 36924 27288 37464 27316
rect 37458 27276 37464 27288
rect 37516 27276 37522 27328
rect 37550 27276 37556 27328
rect 37608 27276 37614 27328
rect 37660 27325 37688 27424
rect 37737 27421 37749 27424
rect 37783 27421 37795 27455
rect 37737 27415 37795 27421
rect 37918 27412 37924 27464
rect 37976 27412 37982 27464
rect 38010 27412 38016 27464
rect 38068 27412 38074 27464
rect 38120 27461 38148 27492
rect 38105 27455 38163 27461
rect 38105 27421 38117 27455
rect 38151 27421 38163 27455
rect 38105 27415 38163 27421
rect 37645 27319 37703 27325
rect 37645 27285 37657 27319
rect 37691 27285 37703 27319
rect 37645 27279 37703 27285
rect 1104 27226 38824 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 38824 27226
rect 1104 27152 38824 27174
rect 3418 27072 3424 27124
rect 3476 27112 3482 27124
rect 3513 27115 3571 27121
rect 3513 27112 3525 27115
rect 3476 27084 3525 27112
rect 3476 27072 3482 27084
rect 3513 27081 3525 27084
rect 3559 27112 3571 27115
rect 3970 27112 3976 27124
rect 3559 27084 3976 27112
rect 3559 27081 3571 27084
rect 3513 27075 3571 27081
rect 3970 27072 3976 27084
rect 4028 27072 4034 27124
rect 12989 27115 13047 27121
rect 8220 27084 9674 27112
rect 6270 27044 6276 27056
rect 4554 27016 6276 27044
rect 6270 27004 6276 27016
rect 6328 27044 6334 27056
rect 8220 27044 8248 27084
rect 9646 27044 9674 27084
rect 12989 27081 13001 27115
rect 13035 27112 13047 27115
rect 13446 27112 13452 27124
rect 13035 27084 13452 27112
rect 13035 27081 13047 27084
rect 12989 27075 13047 27081
rect 13446 27072 13452 27084
rect 13504 27112 13510 27124
rect 17770 27112 17776 27124
rect 13504 27084 17776 27112
rect 13504 27072 13510 27084
rect 17770 27072 17776 27084
rect 17828 27072 17834 27124
rect 18414 27072 18420 27124
rect 18472 27112 18478 27124
rect 19518 27112 19524 27124
rect 18472 27084 19524 27112
rect 18472 27072 18478 27084
rect 19518 27072 19524 27084
rect 19576 27072 19582 27124
rect 21358 27072 21364 27124
rect 21416 27072 21422 27124
rect 21818 27072 21824 27124
rect 21876 27112 21882 27124
rect 22649 27115 22707 27121
rect 22649 27112 22661 27115
rect 21876 27084 22661 27112
rect 21876 27072 21882 27084
rect 22649 27081 22661 27084
rect 22695 27081 22707 27115
rect 22649 27075 22707 27081
rect 25961 27115 26019 27121
rect 25961 27081 25973 27115
rect 26007 27112 26019 27115
rect 33689 27115 33747 27121
rect 26007 27084 26556 27112
rect 26007 27081 26019 27084
rect 25961 27075 26019 27081
rect 12897 27047 12955 27053
rect 6328 27016 8326 27044
rect 9646 27016 10166 27044
rect 6328 27004 6334 27016
rect 12897 27013 12909 27047
rect 12943 27044 12955 27047
rect 13262 27044 13268 27056
rect 12943 27016 13268 27044
rect 12943 27013 12955 27016
rect 12897 27007 12955 27013
rect 13262 27004 13268 27016
rect 13320 27004 13326 27056
rect 15197 27047 15255 27053
rect 15197 27013 15209 27047
rect 15243 27044 15255 27047
rect 15565 27047 15623 27053
rect 15243 27016 15516 27044
rect 15243 27013 15255 27016
rect 15197 27007 15255 27013
rect 15488 26988 15516 27016
rect 15565 27013 15577 27047
rect 15611 27044 15623 27047
rect 16209 27047 16267 27053
rect 15611 27016 15976 27044
rect 15611 27013 15623 27016
rect 15565 27007 15623 27013
rect 2317 26979 2375 26985
rect 2317 26945 2329 26979
rect 2363 26976 2375 26979
rect 2777 26979 2835 26985
rect 2777 26976 2789 26979
rect 2363 26948 2789 26976
rect 2363 26945 2375 26948
rect 2317 26939 2375 26945
rect 2777 26945 2789 26948
rect 2823 26945 2835 26979
rect 2777 26939 2835 26945
rect 3326 26936 3332 26988
rect 3384 26936 3390 26988
rect 5353 26979 5411 26985
rect 5353 26945 5365 26979
rect 5399 26945 5411 26979
rect 5353 26939 5411 26945
rect 5997 26979 6055 26985
rect 5997 26945 6009 26979
rect 6043 26976 6055 26979
rect 6086 26976 6092 26988
rect 6043 26948 6092 26976
rect 6043 26945 6055 26948
rect 5997 26939 6055 26945
rect 1670 26868 1676 26920
rect 1728 26908 1734 26920
rect 1949 26911 2007 26917
rect 1949 26908 1961 26911
rect 1728 26880 1961 26908
rect 1728 26868 1734 26880
rect 1949 26877 1961 26880
rect 1995 26877 2007 26911
rect 1949 26871 2007 26877
rect 2409 26911 2467 26917
rect 2409 26877 2421 26911
rect 2455 26908 2467 26911
rect 3142 26908 3148 26920
rect 2455 26880 3148 26908
rect 2455 26877 2467 26880
rect 2409 26871 2467 26877
rect 3142 26868 3148 26880
rect 3200 26868 3206 26920
rect 3970 26868 3976 26920
rect 4028 26908 4034 26920
rect 4985 26911 5043 26917
rect 4985 26908 4997 26911
rect 4028 26880 4997 26908
rect 4028 26868 4034 26880
rect 4985 26877 4997 26880
rect 5031 26877 5043 26911
rect 4985 26871 5043 26877
rect 5258 26868 5264 26920
rect 5316 26908 5322 26920
rect 5368 26908 5396 26939
rect 6086 26936 6092 26948
rect 6144 26936 6150 26988
rect 6181 26979 6239 26985
rect 6181 26945 6193 26979
rect 6227 26976 6239 26979
rect 6362 26976 6368 26988
rect 6227 26948 6368 26976
rect 6227 26945 6239 26948
rect 6181 26939 6239 26945
rect 6362 26936 6368 26948
rect 6420 26936 6426 26988
rect 13170 26936 13176 26988
rect 13228 26976 13234 26988
rect 13817 26979 13875 26985
rect 13817 26976 13829 26979
rect 13228 26948 13829 26976
rect 13228 26936 13234 26948
rect 13817 26945 13829 26948
rect 13863 26945 13875 26979
rect 13817 26939 13875 26945
rect 13998 26936 14004 26988
rect 14056 26936 14062 26988
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 14277 26979 14335 26985
rect 14277 26945 14289 26979
rect 14323 26976 14335 26979
rect 14366 26976 14372 26988
rect 14323 26948 14372 26976
rect 14323 26945 14335 26948
rect 14277 26939 14335 26945
rect 7561 26911 7619 26917
rect 7561 26908 7573 26911
rect 5316 26880 7573 26908
rect 5316 26868 5322 26880
rect 7561 26877 7573 26880
rect 7607 26877 7619 26911
rect 7561 26871 7619 26877
rect 7837 26911 7895 26917
rect 7837 26877 7849 26911
rect 7883 26908 7895 26911
rect 8294 26908 8300 26920
rect 7883 26880 8300 26908
rect 7883 26877 7895 26880
rect 7837 26871 7895 26877
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 9401 26911 9459 26917
rect 9401 26877 9413 26911
rect 9447 26908 9459 26911
rect 9447 26880 9536 26908
rect 9447 26877 9459 26880
rect 9401 26871 9459 26877
rect 5810 26732 5816 26784
rect 5868 26772 5874 26784
rect 5997 26775 6055 26781
rect 5997 26772 6009 26775
rect 5868 26744 6009 26772
rect 5868 26732 5874 26744
rect 5997 26741 6009 26744
rect 6043 26741 6055 26775
rect 5997 26735 6055 26741
rect 9309 26775 9367 26781
rect 9309 26741 9321 26775
rect 9355 26772 9367 26775
rect 9398 26772 9404 26784
rect 9355 26744 9404 26772
rect 9355 26741 9367 26744
rect 9309 26735 9367 26741
rect 9398 26732 9404 26744
rect 9456 26732 9462 26784
rect 9508 26772 9536 26880
rect 9674 26868 9680 26920
rect 9732 26868 9738 26920
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 12069 26911 12127 26917
rect 12069 26908 12081 26911
rect 11204 26880 12081 26908
rect 11204 26868 11210 26880
rect 12069 26877 12081 26880
rect 12115 26877 12127 26911
rect 12069 26871 12127 26877
rect 13722 26868 13728 26920
rect 13780 26908 13786 26920
rect 14108 26908 14136 26939
rect 13780 26880 14136 26908
rect 13780 26868 13786 26880
rect 13446 26800 13452 26852
rect 13504 26840 13510 26852
rect 14292 26840 14320 26939
rect 14366 26936 14372 26948
rect 14424 26936 14430 26988
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 14476 26948 15117 26976
rect 13504 26812 14320 26840
rect 13504 26800 13510 26812
rect 14476 26784 14504 26948
rect 15105 26945 15117 26948
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 15286 26936 15292 26988
rect 15344 26936 15350 26988
rect 15470 26936 15476 26988
rect 15528 26936 15534 26988
rect 15654 26936 15660 26988
rect 15712 26936 15718 26988
rect 15948 26985 15976 27016
rect 16209 27013 16221 27047
rect 16255 27013 16267 27047
rect 16209 27007 16267 27013
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26945 15991 26979
rect 16224 26976 16252 27007
rect 17862 27004 17868 27056
rect 17920 27044 17926 27056
rect 18877 27047 18935 27053
rect 18877 27044 18889 27047
rect 17920 27016 18889 27044
rect 17920 27004 17926 27016
rect 18877 27013 18889 27016
rect 18923 27013 18935 27047
rect 18877 27007 18935 27013
rect 19245 27047 19303 27053
rect 19245 27013 19257 27047
rect 19291 27044 19303 27047
rect 19334 27044 19340 27056
rect 19291 27016 19340 27044
rect 19291 27013 19303 27016
rect 19245 27007 19303 27013
rect 19334 27004 19340 27016
rect 19392 27044 19398 27056
rect 21913 27047 21971 27053
rect 19392 27016 20116 27044
rect 19392 27004 19398 27016
rect 20088 26988 20116 27016
rect 21913 27013 21925 27047
rect 21959 27044 21971 27047
rect 22370 27044 22376 27056
rect 21959 27016 22376 27044
rect 21959 27013 21971 27016
rect 21913 27007 21971 27013
rect 22370 27004 22376 27016
rect 22428 27004 22434 27056
rect 25866 27004 25872 27056
rect 25924 27044 25930 27056
rect 25924 27016 26372 27044
rect 25924 27004 25930 27016
rect 17954 26976 17960 26988
rect 16224 26948 17960 26976
rect 15933 26939 15991 26945
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 19061 26979 19119 26985
rect 19061 26976 19073 26979
rect 18104 26948 19073 26976
rect 18104 26936 18110 26948
rect 19061 26945 19073 26948
rect 19107 26976 19119 26979
rect 19107 26948 19334 26976
rect 19107 26945 19119 26948
rect 19061 26939 19119 26945
rect 14826 26868 14832 26920
rect 14884 26908 14890 26920
rect 15749 26911 15807 26917
rect 15749 26908 15761 26911
rect 14884 26880 15761 26908
rect 14884 26868 14890 26880
rect 15749 26877 15761 26880
rect 15795 26877 15807 26911
rect 15749 26871 15807 26877
rect 16206 26868 16212 26920
rect 16264 26908 16270 26920
rect 16301 26911 16359 26917
rect 16301 26908 16313 26911
rect 16264 26880 16313 26908
rect 16264 26868 16270 26880
rect 16301 26877 16313 26880
rect 16347 26877 16359 26911
rect 19306 26908 19334 26948
rect 19610 26936 19616 26988
rect 19668 26936 19674 26988
rect 19794 26936 19800 26988
rect 19852 26976 19858 26988
rect 19852 26948 20024 26976
rect 19852 26936 19858 26948
rect 19702 26908 19708 26920
rect 19306 26880 19708 26908
rect 16301 26871 16359 26877
rect 19702 26868 19708 26880
rect 19760 26868 19766 26920
rect 19996 26840 20024 26948
rect 20070 26936 20076 26988
rect 20128 26936 20134 26988
rect 21450 26936 21456 26988
rect 21508 26936 21514 26988
rect 21542 26936 21548 26988
rect 21600 26976 21606 26988
rect 21818 26976 21824 26988
rect 21600 26948 21824 26976
rect 21600 26936 21606 26948
rect 21818 26936 21824 26948
rect 21876 26936 21882 26988
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26976 22063 26979
rect 22738 26976 22744 26988
rect 22051 26948 22744 26976
rect 22051 26945 22063 26948
rect 22005 26939 22063 26945
rect 22738 26936 22744 26948
rect 22796 26936 22802 26988
rect 23290 26936 23296 26988
rect 23348 26936 23354 26988
rect 24210 26936 24216 26988
rect 24268 26936 24274 26988
rect 25590 26936 25596 26988
rect 25648 26936 25654 26988
rect 26050 26936 26056 26988
rect 26108 26936 26114 26988
rect 26237 26979 26295 26985
rect 26237 26945 26249 26979
rect 26283 26945 26295 26979
rect 26237 26939 26295 26945
rect 20622 26868 20628 26920
rect 20680 26908 20686 26920
rect 22186 26908 22192 26920
rect 20680 26880 22192 26908
rect 20680 26868 20686 26880
rect 22186 26868 22192 26880
rect 22244 26868 22250 26920
rect 23566 26868 23572 26920
rect 23624 26868 23630 26920
rect 24121 26911 24179 26917
rect 24121 26877 24133 26911
rect 24167 26908 24179 26911
rect 24489 26911 24547 26917
rect 24489 26908 24501 26911
rect 24167 26880 24501 26908
rect 24167 26877 24179 26880
rect 24121 26871 24179 26877
rect 24489 26877 24501 26880
rect 24535 26877 24547 26911
rect 24489 26871 24547 26877
rect 24578 26868 24584 26920
rect 24636 26908 24642 26920
rect 26252 26908 26280 26939
rect 26344 26917 26372 27016
rect 26418 26936 26424 26988
rect 26476 26936 26482 26988
rect 26528 26976 26556 27084
rect 33689 27081 33701 27115
rect 33735 27112 33747 27115
rect 33778 27112 33784 27124
rect 33735 27084 33784 27112
rect 33735 27081 33747 27084
rect 33689 27075 33747 27081
rect 33778 27072 33784 27084
rect 33836 27072 33842 27124
rect 34882 27072 34888 27124
rect 34940 27112 34946 27124
rect 37001 27115 37059 27121
rect 34940 27084 35756 27112
rect 34940 27072 34946 27084
rect 26694 27004 26700 27056
rect 26752 27044 26758 27056
rect 27709 27047 27767 27053
rect 27709 27044 27721 27047
rect 26752 27016 27721 27044
rect 26752 27004 26758 27016
rect 27709 27013 27721 27016
rect 27755 27013 27767 27047
rect 27709 27007 27767 27013
rect 27982 27004 27988 27056
rect 28040 27044 28046 27056
rect 28905 27047 28963 27053
rect 28905 27044 28917 27047
rect 28040 27016 28917 27044
rect 28040 27004 28046 27016
rect 28905 27013 28917 27016
rect 28951 27013 28963 27047
rect 28905 27007 28963 27013
rect 29638 27004 29644 27056
rect 29696 27004 29702 27056
rect 30837 27047 30895 27053
rect 30837 27013 30849 27047
rect 30883 27044 30895 27047
rect 31202 27044 31208 27056
rect 30883 27016 31208 27044
rect 30883 27013 30895 27016
rect 30837 27007 30895 27013
rect 31202 27004 31208 27016
rect 31260 27044 31266 27056
rect 31260 27016 31754 27044
rect 31260 27004 31266 27016
rect 26605 26979 26663 26985
rect 26605 26976 26617 26979
rect 26528 26948 26617 26976
rect 26605 26945 26617 26948
rect 26651 26976 26663 26979
rect 27525 26979 27583 26985
rect 27525 26976 27537 26979
rect 26651 26948 27537 26976
rect 26651 26945 26663 26948
rect 26605 26939 26663 26945
rect 27525 26945 27537 26948
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 28074 26936 28080 26988
rect 28132 26976 28138 26988
rect 28629 26979 28687 26985
rect 28629 26976 28641 26979
rect 28132 26948 28641 26976
rect 28132 26936 28138 26948
rect 28629 26945 28641 26948
rect 28675 26945 28687 26979
rect 31018 26976 31024 26988
rect 28629 26939 28687 26945
rect 30392 26948 31024 26976
rect 24636 26880 26280 26908
rect 26329 26911 26387 26917
rect 24636 26868 24642 26880
rect 26329 26877 26341 26911
rect 26375 26877 26387 26911
rect 26329 26871 26387 26877
rect 20990 26840 20996 26852
rect 19996 26812 20996 26840
rect 20990 26800 20996 26812
rect 21048 26800 21054 26852
rect 26344 26840 26372 26871
rect 26510 26868 26516 26920
rect 26568 26908 26574 26920
rect 28261 26911 28319 26917
rect 28261 26908 28273 26911
rect 26568 26880 28273 26908
rect 26568 26868 26574 26880
rect 28261 26877 28273 26880
rect 28307 26877 28319 26911
rect 28261 26871 28319 26877
rect 26694 26840 26700 26852
rect 25516 26812 26096 26840
rect 26344 26812 26700 26840
rect 10226 26772 10232 26784
rect 9508 26744 10232 26772
rect 10226 26732 10232 26744
rect 10284 26732 10290 26784
rect 11514 26732 11520 26784
rect 11572 26732 11578 26784
rect 13909 26775 13967 26781
rect 13909 26741 13921 26775
rect 13955 26772 13967 26775
rect 14090 26772 14096 26784
rect 13955 26744 14096 26772
rect 13955 26741 13967 26744
rect 13909 26735 13967 26741
rect 14090 26732 14096 26744
rect 14148 26732 14154 26784
rect 14277 26775 14335 26781
rect 14277 26741 14289 26775
rect 14323 26772 14335 26775
rect 14458 26772 14464 26784
rect 14323 26744 14464 26772
rect 14323 26741 14335 26744
rect 14277 26735 14335 26741
rect 14458 26732 14464 26744
rect 14516 26732 14522 26784
rect 19429 26775 19487 26781
rect 19429 26741 19441 26775
rect 19475 26772 19487 26775
rect 19518 26772 19524 26784
rect 19475 26744 19524 26772
rect 19475 26741 19487 26744
rect 19429 26735 19487 26741
rect 19518 26732 19524 26744
rect 19576 26732 19582 26784
rect 19981 26775 20039 26781
rect 19981 26741 19993 26775
rect 20027 26772 20039 26775
rect 20162 26772 20168 26784
rect 20027 26744 20168 26772
rect 20027 26741 20039 26744
rect 19981 26735 20039 26741
rect 20162 26732 20168 26744
rect 20220 26732 20226 26784
rect 24854 26732 24860 26784
rect 24912 26772 24918 26784
rect 25516 26772 25544 26812
rect 24912 26744 25544 26772
rect 26068 26772 26096 26812
rect 26694 26800 26700 26812
rect 26752 26800 26758 26852
rect 26789 26843 26847 26849
rect 26789 26809 26801 26843
rect 26835 26840 26847 26843
rect 27890 26840 27896 26852
rect 26835 26812 27896 26840
rect 26835 26809 26847 26812
rect 26789 26803 26847 26809
rect 27890 26800 27896 26812
rect 27948 26800 27954 26852
rect 26973 26775 27031 26781
rect 26973 26772 26985 26775
rect 26068 26744 26985 26772
rect 24912 26732 24918 26744
rect 26973 26741 26985 26744
rect 27019 26741 27031 26775
rect 26973 26735 27031 26741
rect 28258 26732 28264 26784
rect 28316 26772 28322 26784
rect 30392 26781 30420 26948
rect 31018 26936 31024 26948
rect 31076 26976 31082 26988
rect 31726 26976 31754 27016
rect 32122 27004 32128 27056
rect 32180 27044 32186 27056
rect 32180 27016 32444 27044
rect 32180 27004 32186 27016
rect 32416 26985 32444 27016
rect 32950 27004 32956 27056
rect 33008 27044 33014 27056
rect 33008 27016 33994 27044
rect 33008 27004 33014 27016
rect 35250 27004 35256 27056
rect 35308 27044 35314 27056
rect 35308 27016 35664 27044
rect 35308 27004 35314 27016
rect 32217 26979 32275 26985
rect 32217 26976 32229 26979
rect 31076 26948 31616 26976
rect 31726 26948 32229 26976
rect 31076 26936 31082 26948
rect 31588 26908 31616 26948
rect 32217 26945 32229 26948
rect 32263 26945 32275 26979
rect 32217 26939 32275 26945
rect 32401 26979 32459 26985
rect 32401 26945 32413 26979
rect 32447 26945 32459 26979
rect 32401 26939 32459 26945
rect 32674 26936 32680 26988
rect 32732 26936 32738 26988
rect 35434 26936 35440 26988
rect 35492 26936 35498 26988
rect 35636 26920 35664 27016
rect 35728 26985 35756 27084
rect 37001 27081 37013 27115
rect 37047 27112 37059 27115
rect 37918 27112 37924 27124
rect 37047 27084 37924 27112
rect 37047 27081 37059 27084
rect 37001 27075 37059 27081
rect 37918 27072 37924 27084
rect 37976 27072 37982 27124
rect 38378 27072 38384 27124
rect 38436 27072 38442 27124
rect 38013 27047 38071 27053
rect 38013 27044 38025 27047
rect 36464 27016 38025 27044
rect 36464 26985 36492 27016
rect 38013 27013 38025 27016
rect 38059 27013 38071 27047
rect 38013 27007 38071 27013
rect 35713 26979 35771 26985
rect 35713 26945 35725 26979
rect 35759 26945 35771 26979
rect 35713 26939 35771 26945
rect 36449 26979 36507 26985
rect 36449 26945 36461 26979
rect 36495 26945 36507 26979
rect 36449 26939 36507 26945
rect 36538 26936 36544 26988
rect 36596 26936 36602 26988
rect 36722 26936 36728 26988
rect 36780 26936 36786 26988
rect 36817 26979 36875 26985
rect 36817 26945 36829 26979
rect 36863 26945 36875 26979
rect 36817 26939 36875 26945
rect 31754 26908 31760 26920
rect 31588 26880 31760 26908
rect 31754 26868 31760 26880
rect 31812 26868 31818 26920
rect 34514 26868 34520 26920
rect 34572 26908 34578 26920
rect 35161 26911 35219 26917
rect 35161 26908 35173 26911
rect 34572 26880 35173 26908
rect 34572 26868 34578 26880
rect 35161 26877 35173 26880
rect 35207 26877 35219 26911
rect 35161 26871 35219 26877
rect 35618 26868 35624 26920
rect 35676 26868 35682 26920
rect 36081 26911 36139 26917
rect 36081 26877 36093 26911
rect 36127 26908 36139 26911
rect 36170 26908 36176 26920
rect 36127 26880 36176 26908
rect 36127 26877 36139 26880
rect 36081 26871 36139 26877
rect 36170 26868 36176 26880
rect 36228 26908 36234 26920
rect 36832 26908 36860 26939
rect 37642 26936 37648 26988
rect 37700 26936 37706 26988
rect 37921 26979 37979 26985
rect 37921 26976 37933 26979
rect 37752 26948 37933 26976
rect 36228 26880 36860 26908
rect 36228 26868 36234 26880
rect 37366 26868 37372 26920
rect 37424 26868 37430 26920
rect 37458 26868 37464 26920
rect 37516 26908 37522 26920
rect 37752 26908 37780 26948
rect 37921 26945 37933 26948
rect 37967 26945 37979 26979
rect 37921 26939 37979 26945
rect 38105 26979 38163 26985
rect 38105 26945 38117 26979
rect 38151 26945 38163 26979
rect 38105 26939 38163 26945
rect 37516 26880 37780 26908
rect 37829 26911 37887 26917
rect 37516 26868 37522 26880
rect 37829 26877 37841 26911
rect 37875 26908 37887 26911
rect 38010 26908 38016 26920
rect 37875 26880 38016 26908
rect 37875 26877 37887 26880
rect 37829 26871 37887 26877
rect 38010 26868 38016 26880
rect 38068 26868 38074 26920
rect 37550 26800 37556 26852
rect 37608 26840 37614 26852
rect 38120 26840 38148 26939
rect 38194 26936 38200 26988
rect 38252 26936 38258 26988
rect 37608 26812 38148 26840
rect 37608 26800 37614 26812
rect 30377 26775 30435 26781
rect 30377 26772 30389 26775
rect 28316 26744 30389 26772
rect 28316 26732 28322 26744
rect 30377 26741 30389 26744
rect 30423 26741 30435 26775
rect 30377 26735 30435 26741
rect 30742 26732 30748 26784
rect 30800 26772 30806 26784
rect 31113 26775 31171 26781
rect 31113 26772 31125 26775
rect 30800 26744 31125 26772
rect 30800 26732 30806 26744
rect 31113 26741 31125 26744
rect 31159 26741 31171 26775
rect 31113 26735 31171 26741
rect 32861 26775 32919 26781
rect 32861 26741 32873 26775
rect 32907 26772 32919 26775
rect 33594 26772 33600 26784
rect 32907 26744 33600 26772
rect 32907 26741 32919 26744
rect 32861 26735 32919 26741
rect 33594 26732 33600 26744
rect 33652 26732 33658 26784
rect 37458 26732 37464 26784
rect 37516 26732 37522 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 3053 26571 3111 26577
rect 3053 26537 3065 26571
rect 3099 26568 3111 26571
rect 3142 26568 3148 26580
rect 3099 26540 3148 26568
rect 3099 26537 3111 26540
rect 3053 26531 3111 26537
rect 3142 26528 3148 26540
rect 3200 26528 3206 26580
rect 3970 26528 3976 26580
rect 4028 26528 4034 26580
rect 5258 26528 5264 26580
rect 5316 26568 5322 26580
rect 5316 26540 6500 26568
rect 5316 26528 5322 26540
rect 3160 26500 3188 26528
rect 3160 26472 4016 26500
rect 2869 26435 2927 26441
rect 2869 26401 2881 26435
rect 2915 26432 2927 26435
rect 2915 26404 3832 26432
rect 2915 26401 2927 26404
rect 2869 26395 2927 26401
rect 2774 26324 2780 26376
rect 2832 26324 2838 26376
rect 2961 26367 3019 26373
rect 2961 26333 2973 26367
rect 3007 26364 3019 26367
rect 3237 26367 3295 26373
rect 3237 26364 3249 26367
rect 3007 26336 3249 26364
rect 3007 26333 3019 26336
rect 2961 26327 3019 26333
rect 3237 26333 3249 26336
rect 3283 26364 3295 26367
rect 3326 26364 3332 26376
rect 3283 26336 3332 26364
rect 3283 26333 3295 26336
rect 3237 26327 3295 26333
rect 3326 26324 3332 26336
rect 3384 26324 3390 26376
rect 3418 26324 3424 26376
rect 3476 26324 3482 26376
rect 3804 26373 3832 26404
rect 3988 26373 4016 26472
rect 5258 26432 5264 26444
rect 4632 26404 5264 26432
rect 4632 26373 4660 26404
rect 5258 26392 5264 26404
rect 5316 26392 5322 26444
rect 6472 26441 6500 26540
rect 8294 26528 8300 26580
rect 8352 26528 8358 26580
rect 9674 26528 9680 26580
rect 9732 26568 9738 26580
rect 9861 26571 9919 26577
rect 9861 26568 9873 26571
rect 9732 26540 9873 26568
rect 9732 26528 9738 26540
rect 9861 26537 9873 26540
rect 9907 26537 9919 26571
rect 9861 26531 9919 26537
rect 13170 26528 13176 26580
rect 13228 26528 13234 26580
rect 13262 26528 13268 26580
rect 13320 26568 13326 26580
rect 19429 26571 19487 26577
rect 19429 26568 19441 26571
rect 13320 26540 19441 26568
rect 13320 26528 13326 26540
rect 19429 26537 19441 26540
rect 19475 26537 19487 26571
rect 19429 26531 19487 26537
rect 19702 26528 19708 26580
rect 19760 26568 19766 26580
rect 20346 26568 20352 26580
rect 19760 26540 20352 26568
rect 19760 26528 19766 26540
rect 20346 26528 20352 26540
rect 20404 26528 20410 26580
rect 20438 26528 20444 26580
rect 20496 26528 20502 26580
rect 23566 26528 23572 26580
rect 23624 26568 23630 26580
rect 24397 26571 24455 26577
rect 24397 26568 24409 26571
rect 23624 26540 24409 26568
rect 23624 26528 23630 26540
rect 24397 26537 24409 26540
rect 24443 26537 24455 26571
rect 24397 26531 24455 26537
rect 25501 26571 25559 26577
rect 25501 26537 25513 26571
rect 25547 26568 25559 26571
rect 26510 26568 26516 26580
rect 25547 26540 26516 26568
rect 25547 26537 25559 26540
rect 25501 26531 25559 26537
rect 26510 26528 26516 26540
rect 26568 26528 26574 26580
rect 28077 26571 28135 26577
rect 28077 26537 28089 26571
rect 28123 26568 28135 26571
rect 28166 26568 28172 26580
rect 28123 26540 28172 26568
rect 28123 26537 28135 26540
rect 28077 26531 28135 26537
rect 28166 26528 28172 26540
rect 28224 26528 28230 26580
rect 29638 26528 29644 26580
rect 29696 26568 29702 26580
rect 30193 26571 30251 26577
rect 30193 26568 30205 26571
rect 29696 26540 30205 26568
rect 29696 26528 29702 26540
rect 30193 26537 30205 26540
rect 30239 26537 30251 26571
rect 30193 26531 30251 26537
rect 35253 26571 35311 26577
rect 35253 26537 35265 26571
rect 35299 26568 35311 26571
rect 35342 26568 35348 26580
rect 35299 26540 35348 26568
rect 35299 26537 35311 26540
rect 35253 26531 35311 26537
rect 35342 26528 35348 26540
rect 35400 26528 35406 26580
rect 35437 26571 35495 26577
rect 35437 26537 35449 26571
rect 35483 26568 35495 26571
rect 35618 26568 35624 26580
rect 35483 26540 35624 26568
rect 35483 26537 35495 26540
rect 35437 26531 35495 26537
rect 35618 26528 35624 26540
rect 35676 26528 35682 26580
rect 36538 26528 36544 26580
rect 36596 26528 36602 26580
rect 37461 26571 37519 26577
rect 37461 26537 37473 26571
rect 37507 26568 37519 26571
rect 37734 26568 37740 26580
rect 37507 26540 37740 26568
rect 37507 26537 37519 26540
rect 37461 26531 37519 26537
rect 37734 26528 37740 26540
rect 37792 26528 37798 26580
rect 15378 26500 15384 26512
rect 13306 26472 15384 26500
rect 6457 26435 6515 26441
rect 6457 26401 6469 26435
rect 6503 26401 6515 26435
rect 6457 26395 6515 26401
rect 8110 26392 8116 26444
rect 8168 26432 8174 26444
rect 8205 26435 8263 26441
rect 8205 26432 8217 26435
rect 8168 26404 8217 26432
rect 8168 26392 8174 26404
rect 8205 26401 8217 26404
rect 8251 26401 8263 26435
rect 8205 26395 8263 26401
rect 10226 26392 10232 26444
rect 10284 26392 10290 26444
rect 3789 26367 3847 26373
rect 3789 26333 3801 26367
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26333 4675 26367
rect 4617 26327 4675 26333
rect 2682 26256 2688 26308
rect 2740 26296 2746 26308
rect 4632 26296 4660 26327
rect 8478 26324 8484 26376
rect 8536 26324 8542 26376
rect 8570 26324 8576 26376
rect 8628 26364 8634 26376
rect 8665 26367 8723 26373
rect 8665 26364 8677 26367
rect 8628 26336 8677 26364
rect 8628 26324 8634 26336
rect 8665 26333 8677 26336
rect 8711 26333 8723 26367
rect 8665 26327 8723 26333
rect 8757 26367 8815 26373
rect 8757 26333 8769 26367
rect 8803 26364 8815 26367
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8803 26336 9137 26364
rect 8803 26333 8815 26336
rect 8757 26327 8815 26333
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 2740 26268 4660 26296
rect 4893 26299 4951 26305
rect 2740 26256 2746 26268
rect 4893 26265 4905 26299
rect 4939 26296 4951 26299
rect 6270 26296 6276 26308
rect 4939 26268 5304 26296
rect 6118 26268 6276 26296
rect 4939 26265 4951 26268
rect 4893 26259 4951 26265
rect 5276 26228 5304 26268
rect 6270 26256 6276 26268
rect 6328 26296 6334 26308
rect 6733 26299 6791 26305
rect 6328 26268 6684 26296
rect 6328 26256 6334 26268
rect 5626 26228 5632 26240
rect 5276 26200 5632 26228
rect 5626 26188 5632 26200
rect 5684 26188 5690 26240
rect 6362 26188 6368 26240
rect 6420 26188 6426 26240
rect 6656 26228 6684 26268
rect 6733 26265 6745 26299
rect 6779 26296 6791 26299
rect 7006 26296 7012 26308
rect 6779 26268 7012 26296
rect 6779 26265 6791 26268
rect 6733 26259 6791 26265
rect 7006 26256 7012 26268
rect 7064 26256 7070 26308
rect 8680 26296 8708 26327
rect 9490 26324 9496 26376
rect 9548 26364 9554 26376
rect 9677 26367 9735 26373
rect 9677 26364 9689 26367
rect 9548 26336 9689 26364
rect 9548 26324 9554 26336
rect 9677 26333 9689 26336
rect 9723 26333 9735 26367
rect 9677 26327 9735 26333
rect 9766 26324 9772 26376
rect 9824 26364 9830 26376
rect 9861 26367 9919 26373
rect 9861 26364 9873 26367
rect 9824 26336 9873 26364
rect 9824 26324 9830 26336
rect 9861 26333 9873 26336
rect 9907 26333 9919 26367
rect 10042 26364 10048 26376
rect 9861 26327 9919 26333
rect 9968 26336 10048 26364
rect 9968 26296 9996 26336
rect 10042 26324 10048 26336
rect 10100 26324 10106 26376
rect 13306 26373 13334 26472
rect 15378 26460 15384 26472
rect 15436 26460 15442 26512
rect 15470 26460 15476 26512
rect 15528 26500 15534 26512
rect 17865 26503 17923 26509
rect 15528 26472 16252 26500
rect 15528 26460 15534 26472
rect 14090 26392 14096 26444
rect 14148 26392 14154 26444
rect 14553 26435 14611 26441
rect 14553 26401 14565 26435
rect 14599 26432 14611 26435
rect 15562 26432 15568 26444
rect 14599 26404 15568 26432
rect 14599 26401 14611 26404
rect 14553 26395 14611 26401
rect 15562 26392 15568 26404
rect 15620 26392 15626 26444
rect 15746 26392 15752 26444
rect 15804 26432 15810 26444
rect 16224 26441 16252 26472
rect 17865 26469 17877 26503
rect 17911 26500 17923 26503
rect 18874 26500 18880 26512
rect 17911 26472 18880 26500
rect 17911 26469 17923 26472
rect 17865 26463 17923 26469
rect 18874 26460 18880 26472
rect 18932 26460 18938 26512
rect 19058 26460 19064 26512
rect 19116 26500 19122 26512
rect 19116 26472 20392 26500
rect 19116 26460 19122 26472
rect 15841 26435 15899 26441
rect 15841 26432 15853 26435
rect 15804 26404 15853 26432
rect 15804 26392 15810 26404
rect 15841 26401 15853 26404
rect 15887 26401 15899 26435
rect 15841 26395 15899 26401
rect 16209 26435 16267 26441
rect 16209 26401 16221 26435
rect 16255 26401 16267 26435
rect 16209 26395 16267 26401
rect 16326 26435 16384 26441
rect 16326 26401 16338 26435
rect 16372 26432 16384 26435
rect 16482 26432 16488 26444
rect 16372 26404 16488 26432
rect 16372 26401 16384 26404
rect 16326 26395 16384 26401
rect 16482 26392 16488 26404
rect 16540 26392 16546 26444
rect 17681 26435 17739 26441
rect 17681 26401 17693 26435
rect 17727 26432 17739 26435
rect 19521 26435 19579 26441
rect 19521 26432 19533 26435
rect 17727 26404 19533 26432
rect 17727 26401 17739 26404
rect 17681 26395 17739 26401
rect 18340 26376 18368 26404
rect 19521 26401 19533 26404
rect 19567 26401 19579 26435
rect 19521 26395 19579 26401
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 13265 26367 13334 26373
rect 13265 26333 13277 26367
rect 13311 26338 13334 26367
rect 13311 26333 13323 26338
rect 13265 26327 13323 26333
rect 7116 26268 7222 26296
rect 8680 26268 9996 26296
rect 7116 26228 7144 26268
rect 10502 26256 10508 26308
rect 10560 26256 10566 26308
rect 11790 26296 11796 26308
rect 11730 26268 11796 26296
rect 11790 26256 11796 26268
rect 11848 26296 11854 26308
rect 12618 26296 12624 26308
rect 11848 26268 12624 26296
rect 11848 26256 11854 26268
rect 12618 26256 12624 26268
rect 12676 26256 12682 26308
rect 13096 26296 13124 26327
rect 13446 26324 13452 26376
rect 13504 26364 13510 26376
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 13504 26336 13553 26364
rect 13504 26324 13510 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13634 26367 13692 26373
rect 13634 26333 13646 26367
rect 13680 26364 13692 26367
rect 13722 26364 13728 26376
rect 13680 26336 13728 26364
rect 13680 26333 13692 26336
rect 13634 26327 13692 26333
rect 13464 26296 13492 26324
rect 13648 26296 13676 26327
rect 13722 26324 13728 26336
rect 13780 26324 13786 26376
rect 14458 26324 14464 26376
rect 14516 26324 14522 26376
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26333 15347 26367
rect 15289 26327 15347 26333
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26364 15531 26367
rect 15654 26364 15660 26376
rect 15519 26336 15660 26364
rect 15519 26333 15531 26336
rect 15473 26327 15531 26333
rect 14185 26299 14243 26305
rect 14185 26296 14197 26299
rect 13096 26268 13492 26296
rect 13556 26268 13676 26296
rect 13832 26268 14197 26296
rect 6656 26200 7144 26228
rect 9582 26188 9588 26240
rect 9640 26228 9646 26240
rect 11974 26228 11980 26240
rect 9640 26200 11980 26228
rect 9640 26188 9646 26200
rect 11974 26188 11980 26200
rect 12032 26188 12038 26240
rect 13078 26188 13084 26240
rect 13136 26228 13142 26240
rect 13556 26228 13584 26268
rect 13136 26200 13584 26228
rect 13136 26188 13142 26200
rect 13630 26188 13636 26240
rect 13688 26228 13694 26240
rect 13832 26228 13860 26268
rect 14185 26265 14197 26268
rect 14231 26296 14243 26299
rect 15194 26296 15200 26308
rect 14231 26268 15200 26296
rect 14231 26265 14243 26268
rect 14185 26259 14243 26265
rect 15194 26256 15200 26268
rect 15252 26256 15258 26308
rect 15304 26296 15332 26327
rect 15654 26324 15660 26336
rect 15712 26324 15718 26376
rect 17310 26324 17316 26376
rect 17368 26324 17374 26376
rect 17494 26373 17500 26376
rect 17467 26367 17500 26373
rect 17467 26333 17479 26367
rect 17467 26327 17500 26333
rect 17494 26324 17500 26327
rect 17552 26324 17558 26376
rect 17773 26367 17831 26373
rect 17773 26363 17785 26367
rect 17696 26335 17785 26363
rect 17328 26296 17356 26324
rect 17696 26296 17724 26335
rect 17773 26333 17785 26335
rect 17819 26333 17831 26367
rect 17773 26327 17831 26333
rect 17954 26324 17960 26376
rect 18012 26324 18018 26376
rect 18138 26324 18144 26376
rect 18196 26324 18202 26376
rect 18322 26324 18328 26376
rect 18380 26324 18386 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18601 26367 18659 26373
rect 18601 26364 18613 26367
rect 18472 26336 18613 26364
rect 18472 26324 18478 26336
rect 18601 26333 18613 26336
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 18782 26324 18788 26376
rect 18840 26324 18846 26376
rect 18966 26324 18972 26376
rect 19024 26364 19030 26376
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 19024 26336 19441 26364
rect 19024 26324 19030 26336
rect 19429 26333 19441 26336
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 15304 26268 16160 26296
rect 17328 26268 17724 26296
rect 13688 26200 13860 26228
rect 13909 26231 13967 26237
rect 13688 26188 13694 26200
rect 13909 26197 13921 26231
rect 13955 26228 13967 26231
rect 13998 26228 14004 26240
rect 13955 26200 14004 26228
rect 13955 26197 13967 26200
rect 13909 26191 13967 26197
rect 13998 26188 14004 26200
rect 14056 26228 14062 26240
rect 14458 26228 14464 26240
rect 14056 26200 14464 26228
rect 14056 26188 14062 26200
rect 14458 26188 14464 26200
rect 14516 26188 14522 26240
rect 14734 26188 14740 26240
rect 14792 26188 14798 26240
rect 15286 26188 15292 26240
rect 15344 26188 15350 26240
rect 16132 26237 16160 26268
rect 16117 26231 16175 26237
rect 16117 26197 16129 26231
rect 16163 26228 16175 26231
rect 16206 26228 16212 26240
rect 16163 26200 16212 26228
rect 16163 26197 16175 26200
rect 16117 26191 16175 26197
rect 16206 26188 16212 26200
rect 16264 26188 16270 26240
rect 16482 26188 16488 26240
rect 16540 26188 16546 26240
rect 17494 26188 17500 26240
rect 17552 26228 17558 26240
rect 17972 26228 18000 26324
rect 18156 26296 18184 26324
rect 19058 26296 19064 26308
rect 18156 26268 19064 26296
rect 19058 26256 19064 26268
rect 19116 26256 19122 26308
rect 19536 26296 19564 26395
rect 19978 26392 19984 26444
rect 20036 26432 20042 26444
rect 20257 26435 20315 26441
rect 20257 26432 20269 26435
rect 20036 26404 20269 26432
rect 20036 26392 20042 26404
rect 20257 26401 20269 26404
rect 20303 26401 20315 26435
rect 20257 26395 20315 26401
rect 19610 26324 19616 26376
rect 19668 26364 19674 26376
rect 20364 26373 20392 26472
rect 20456 26441 20484 26528
rect 20717 26503 20775 26509
rect 20717 26469 20729 26503
rect 20763 26500 20775 26503
rect 21634 26500 21640 26512
rect 20763 26472 21640 26500
rect 20763 26469 20775 26472
rect 20717 26463 20775 26469
rect 21634 26460 21640 26472
rect 21692 26460 21698 26512
rect 24578 26460 24584 26512
rect 24636 26500 24642 26512
rect 24636 26472 24992 26500
rect 24636 26460 24642 26472
rect 20441 26435 20499 26441
rect 20441 26401 20453 26435
rect 20487 26401 20499 26435
rect 20441 26395 20499 26401
rect 19889 26367 19947 26373
rect 19889 26364 19901 26367
rect 19668 26336 19901 26364
rect 19668 26324 19674 26336
rect 19889 26333 19901 26336
rect 19935 26364 19947 26367
rect 20349 26367 20407 26373
rect 19935 26336 20300 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 20073 26299 20131 26305
rect 20073 26296 20085 26299
rect 19536 26268 20085 26296
rect 20073 26265 20085 26268
rect 20119 26265 20131 26299
rect 20272 26296 20300 26336
rect 20349 26333 20361 26367
rect 20395 26333 20407 26367
rect 20349 26327 20407 26333
rect 20809 26367 20867 26373
rect 20809 26333 20821 26367
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 20824 26296 20852 26327
rect 24118 26324 24124 26376
rect 24176 26364 24182 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 24176 26336 24593 26364
rect 24176 26324 24182 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 24762 26324 24768 26376
rect 24820 26324 24826 26376
rect 24854 26324 24860 26376
rect 24912 26324 24918 26376
rect 24964 26373 24992 26472
rect 27798 26460 27804 26512
rect 27856 26500 27862 26512
rect 28810 26500 28816 26512
rect 27856 26472 28816 26500
rect 27856 26460 27862 26472
rect 28810 26460 28816 26472
rect 28868 26500 28874 26512
rect 31202 26500 31208 26512
rect 28868 26472 29776 26500
rect 28868 26460 28874 26472
rect 27249 26435 27307 26441
rect 27249 26401 27261 26435
rect 27295 26432 27307 26435
rect 27614 26432 27620 26444
rect 27295 26404 27620 26432
rect 27295 26401 27307 26404
rect 27249 26395 27307 26401
rect 27614 26392 27620 26404
rect 27672 26392 27678 26444
rect 27890 26392 27896 26444
rect 27948 26392 27954 26444
rect 28460 26404 29316 26432
rect 24949 26367 25007 26373
rect 24949 26333 24961 26367
rect 24995 26333 25007 26367
rect 24949 26327 25007 26333
rect 25133 26367 25191 26373
rect 25133 26333 25145 26367
rect 25179 26333 25191 26367
rect 25133 26327 25191 26333
rect 20272 26268 20852 26296
rect 23845 26299 23903 26305
rect 20073 26259 20131 26265
rect 23845 26265 23857 26299
rect 23891 26265 23903 26299
rect 23845 26259 23903 26265
rect 17552 26200 18000 26228
rect 18509 26231 18567 26237
rect 17552 26188 17558 26200
rect 18509 26197 18521 26231
rect 18555 26228 18567 26231
rect 18598 26228 18604 26240
rect 18555 26200 18604 26228
rect 18555 26197 18567 26200
rect 18509 26191 18567 26197
rect 18598 26188 18604 26200
rect 18656 26188 18662 26240
rect 18690 26188 18696 26240
rect 18748 26188 18754 26240
rect 19797 26231 19855 26237
rect 19797 26197 19809 26231
rect 19843 26228 19855 26231
rect 20622 26228 20628 26240
rect 19843 26200 20628 26228
rect 19843 26197 19855 26200
rect 19797 26191 19855 26197
rect 20622 26188 20628 26200
rect 20680 26188 20686 26240
rect 20806 26188 20812 26240
rect 20864 26228 20870 26240
rect 20901 26231 20959 26237
rect 20901 26228 20913 26231
rect 20864 26200 20913 26228
rect 20864 26188 20870 26200
rect 20901 26197 20913 26200
rect 20947 26197 20959 26231
rect 23860 26228 23888 26259
rect 24026 26256 24032 26308
rect 24084 26256 24090 26308
rect 24213 26299 24271 26305
rect 24213 26265 24225 26299
rect 24259 26296 24271 26299
rect 25148 26296 25176 26327
rect 28258 26324 28264 26376
rect 28316 26324 28322 26376
rect 28460 26373 28488 26404
rect 28445 26367 28503 26373
rect 28445 26333 28457 26367
rect 28491 26333 28503 26367
rect 28445 26327 28503 26333
rect 29086 26324 29092 26376
rect 29144 26324 29150 26376
rect 29288 26373 29316 26404
rect 29748 26373 29776 26472
rect 29932 26472 31208 26500
rect 29822 26392 29828 26444
rect 29880 26432 29886 26444
rect 29932 26441 29960 26472
rect 31202 26460 31208 26472
rect 31260 26460 31266 26512
rect 37366 26460 37372 26512
rect 37424 26500 37430 26512
rect 38010 26500 38016 26512
rect 37424 26472 38016 26500
rect 37424 26460 37430 26472
rect 38010 26460 38016 26472
rect 38068 26460 38074 26512
rect 29917 26435 29975 26441
rect 29917 26432 29929 26435
rect 29880 26404 29929 26432
rect 29880 26392 29886 26404
rect 29917 26401 29929 26404
rect 29963 26401 29975 26435
rect 29917 26395 29975 26401
rect 30098 26392 30104 26444
rect 30156 26432 30162 26444
rect 30561 26435 30619 26441
rect 30561 26432 30573 26435
rect 30156 26404 30573 26432
rect 30156 26392 30162 26404
rect 30561 26401 30573 26404
rect 30607 26401 30619 26435
rect 30561 26395 30619 26401
rect 37458 26392 37464 26444
rect 37516 26432 37522 26444
rect 37645 26435 37703 26441
rect 37645 26432 37657 26435
rect 37516 26404 37657 26432
rect 37516 26392 37522 26404
rect 37645 26401 37657 26404
rect 37691 26401 37703 26435
rect 37645 26395 37703 26401
rect 29273 26367 29331 26373
rect 29273 26333 29285 26367
rect 29319 26364 29331 26367
rect 29549 26367 29607 26373
rect 29549 26364 29561 26367
rect 29319 26336 29561 26364
rect 29319 26333 29331 26336
rect 29273 26327 29331 26333
rect 29549 26333 29561 26336
rect 29595 26333 29607 26367
rect 29549 26327 29607 26333
rect 29733 26367 29791 26373
rect 29733 26333 29745 26367
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 29840 26336 30512 26364
rect 24259 26268 25176 26296
rect 24259 26265 24271 26268
rect 24213 26259 24271 26265
rect 25590 26256 25596 26308
rect 25648 26296 25654 26308
rect 26973 26299 27031 26305
rect 25648 26268 25806 26296
rect 25648 26256 25654 26268
rect 26973 26265 26985 26299
rect 27019 26296 27031 26299
rect 27341 26299 27399 26305
rect 27341 26296 27353 26299
rect 27019 26268 27353 26296
rect 27019 26265 27031 26268
rect 26973 26259 27031 26265
rect 27341 26265 27353 26268
rect 27387 26265 27399 26299
rect 27341 26259 27399 26265
rect 28534 26256 28540 26308
rect 28592 26296 28598 26308
rect 29840 26296 29868 26336
rect 28592 26268 29868 26296
rect 28592 26256 28598 26268
rect 30098 26256 30104 26308
rect 30156 26256 30162 26308
rect 30484 26305 30512 26336
rect 31018 26324 31024 26376
rect 31076 26324 31082 26376
rect 31202 26324 31208 26376
rect 31260 26324 31266 26376
rect 33778 26324 33784 26376
rect 33836 26364 33842 26376
rect 35069 26367 35127 26373
rect 35069 26364 35081 26367
rect 33836 26336 35081 26364
rect 33836 26324 33842 26336
rect 35069 26333 35081 26336
rect 35115 26364 35127 26367
rect 35345 26367 35403 26373
rect 35345 26364 35357 26367
rect 35115 26336 35357 26364
rect 35115 26333 35127 26336
rect 35069 26327 35127 26333
rect 35345 26333 35357 26336
rect 35391 26333 35403 26367
rect 35345 26327 35403 26333
rect 35529 26367 35587 26373
rect 35529 26333 35541 26367
rect 35575 26333 35587 26367
rect 35529 26327 35587 26333
rect 35897 26367 35955 26373
rect 35897 26333 35909 26367
rect 35943 26364 35955 26367
rect 35986 26364 35992 26376
rect 35943 26336 35992 26364
rect 35943 26333 35955 26336
rect 35897 26327 35955 26333
rect 30469 26299 30527 26305
rect 30469 26265 30481 26299
rect 30515 26296 30527 26299
rect 31662 26296 31668 26308
rect 30515 26268 31668 26296
rect 30515 26265 30527 26268
rect 30469 26259 30527 26265
rect 31662 26256 31668 26268
rect 31720 26256 31726 26308
rect 32674 26256 32680 26308
rect 32732 26296 32738 26308
rect 34885 26299 34943 26305
rect 34885 26296 34897 26299
rect 32732 26268 34897 26296
rect 32732 26256 32738 26268
rect 34885 26265 34897 26268
rect 34931 26296 34943 26299
rect 35544 26296 35572 26327
rect 35986 26324 35992 26336
rect 36044 26324 36050 26376
rect 36078 26324 36084 26376
rect 36136 26324 36142 26376
rect 36170 26324 36176 26376
rect 36228 26324 36234 26376
rect 36265 26367 36323 26373
rect 36265 26333 36277 26367
rect 36311 26364 36323 26367
rect 36722 26364 36728 26376
rect 36311 26336 36728 26364
rect 36311 26333 36323 26336
rect 36265 26327 36323 26333
rect 36722 26324 36728 26336
rect 36780 26324 36786 26376
rect 37366 26324 37372 26376
rect 37424 26364 37430 26376
rect 37737 26367 37795 26373
rect 37737 26364 37749 26367
rect 37424 26336 37749 26364
rect 37424 26324 37430 26336
rect 37737 26333 37749 26336
rect 37783 26333 37795 26367
rect 37737 26327 37795 26333
rect 34931 26268 35572 26296
rect 34931 26265 34943 26268
rect 34885 26259 34943 26265
rect 37642 26256 37648 26308
rect 37700 26296 37706 26308
rect 38105 26299 38163 26305
rect 38105 26296 38117 26299
rect 37700 26268 38117 26296
rect 37700 26256 37706 26268
rect 38105 26265 38117 26268
rect 38151 26265 38163 26299
rect 38105 26259 38163 26265
rect 24302 26228 24308 26240
rect 23860 26200 24308 26228
rect 20901 26191 20959 26197
rect 24302 26188 24308 26200
rect 24360 26188 24366 26240
rect 29178 26188 29184 26240
rect 29236 26188 29242 26240
rect 30926 26188 30932 26240
rect 30984 26228 30990 26240
rect 31021 26231 31079 26237
rect 31021 26228 31033 26231
rect 30984 26200 31033 26228
rect 30984 26188 30990 26200
rect 31021 26197 31033 26200
rect 31067 26197 31079 26231
rect 31021 26191 31079 26197
rect 1104 26138 38824 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 38824 26138
rect 1104 26064 38824 26086
rect 8478 25984 8484 26036
rect 8536 26024 8542 26036
rect 8757 26027 8815 26033
rect 8757 26024 8769 26027
rect 8536 25996 8769 26024
rect 8536 25984 8542 25996
rect 8757 25993 8769 25996
rect 8803 25993 8815 26027
rect 9490 26024 9496 26036
rect 8757 25987 8815 25993
rect 9324 25996 9496 26024
rect 5626 25916 5632 25968
rect 5684 25916 5690 25968
rect 5997 25959 6055 25965
rect 5997 25925 6009 25959
rect 6043 25956 6055 25959
rect 6365 25959 6423 25965
rect 6365 25956 6377 25959
rect 6043 25928 6377 25956
rect 6043 25925 6055 25928
rect 5997 25919 6055 25925
rect 6365 25925 6377 25928
rect 6411 25925 6423 25959
rect 8570 25956 8576 25968
rect 6365 25919 6423 25925
rect 7208 25928 7512 25956
rect 3234 25848 3240 25900
rect 3292 25848 3298 25900
rect 3326 25848 3332 25900
rect 3384 25888 3390 25900
rect 3421 25891 3479 25897
rect 3421 25888 3433 25891
rect 3384 25860 3433 25888
rect 3384 25848 3390 25860
rect 3421 25857 3433 25860
rect 3467 25857 3479 25891
rect 3421 25851 3479 25857
rect 5810 25848 5816 25900
rect 5868 25848 5874 25900
rect 6086 25848 6092 25900
rect 6144 25848 6150 25900
rect 7208 25897 7236 25928
rect 7193 25891 7251 25897
rect 7193 25857 7205 25891
rect 7239 25857 7251 25891
rect 7193 25851 7251 25857
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25857 7435 25891
rect 7377 25851 7435 25857
rect 5721 25823 5779 25829
rect 5721 25789 5733 25823
rect 5767 25820 5779 25823
rect 5994 25820 6000 25832
rect 5767 25792 6000 25820
rect 5767 25789 5779 25792
rect 5721 25783 5779 25789
rect 5994 25780 6000 25792
rect 6052 25780 6058 25832
rect 6104 25752 6132 25848
rect 6362 25780 6368 25832
rect 6420 25820 6426 25832
rect 6917 25823 6975 25829
rect 6917 25820 6929 25823
rect 6420 25792 6929 25820
rect 6420 25780 6426 25792
rect 6917 25789 6929 25792
rect 6963 25789 6975 25823
rect 6917 25783 6975 25789
rect 6822 25752 6828 25764
rect 6104 25724 6828 25752
rect 6822 25712 6828 25724
rect 6880 25752 6886 25764
rect 7392 25752 7420 25851
rect 7484 25829 7512 25928
rect 7668 25928 8576 25956
rect 7668 25897 7696 25928
rect 8570 25916 8576 25928
rect 8628 25956 8634 25968
rect 9324 25965 9352 25996
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 9582 25984 9588 26036
rect 9640 25984 9646 26036
rect 11514 26024 11520 26036
rect 9784 25996 11520 26024
rect 9784 25965 9812 25996
rect 11514 25984 11520 25996
rect 11572 25984 11578 26036
rect 13170 25984 13176 26036
rect 13228 26024 13234 26036
rect 13265 26027 13323 26033
rect 13265 26024 13277 26027
rect 13228 25996 13277 26024
rect 13228 25984 13234 25996
rect 13265 25993 13277 25996
rect 13311 25993 13323 26027
rect 13265 25987 13323 25993
rect 13633 26027 13691 26033
rect 13633 25993 13645 26027
rect 13679 25993 13691 26027
rect 13633 25987 13691 25993
rect 9093 25959 9151 25965
rect 9093 25956 9105 25959
rect 8628 25928 9105 25956
rect 8628 25916 8634 25928
rect 9093 25925 9105 25928
rect 9139 25925 9151 25959
rect 9093 25919 9151 25925
rect 9309 25959 9367 25965
rect 9309 25925 9321 25959
rect 9355 25925 9367 25959
rect 9309 25919 9367 25925
rect 9769 25959 9827 25965
rect 9769 25925 9781 25959
rect 9815 25925 9827 25959
rect 9769 25919 9827 25925
rect 10134 25916 10140 25968
rect 10192 25956 10198 25968
rect 10657 25959 10715 25965
rect 10657 25956 10669 25959
rect 10192 25928 10669 25956
rect 10192 25916 10198 25928
rect 10657 25925 10669 25928
rect 10703 25925 10715 25959
rect 10657 25919 10715 25925
rect 10873 25959 10931 25965
rect 10873 25925 10885 25959
rect 10919 25956 10931 25959
rect 10919 25928 12020 25956
rect 10919 25925 10931 25928
rect 10873 25919 10931 25925
rect 11992 25900 12020 25928
rect 7653 25891 7711 25897
rect 7653 25857 7665 25891
rect 7699 25857 7711 25891
rect 8665 25891 8723 25897
rect 8665 25888 8677 25891
rect 7653 25851 7711 25857
rect 7760 25860 8677 25888
rect 7469 25823 7527 25829
rect 7469 25789 7481 25823
rect 7515 25820 7527 25823
rect 7760 25820 7788 25860
rect 8665 25857 8677 25860
rect 8711 25857 8723 25891
rect 8665 25851 8723 25857
rect 8846 25848 8852 25900
rect 8904 25848 8910 25900
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25857 9551 25891
rect 9493 25851 9551 25857
rect 10045 25891 10103 25897
rect 10045 25857 10057 25891
rect 10091 25888 10103 25891
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 10091 25886 10640 25888
rect 10796 25886 11529 25888
rect 10091 25860 11529 25886
rect 10091 25857 10103 25860
rect 10612 25858 10824 25860
rect 10045 25851 10103 25857
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 7515 25792 7788 25820
rect 7837 25823 7895 25829
rect 7515 25789 7527 25792
rect 7469 25783 7527 25789
rect 7837 25789 7849 25823
rect 7883 25820 7895 25823
rect 8386 25820 8392 25832
rect 7883 25792 8392 25820
rect 7883 25789 7895 25792
rect 7837 25783 7895 25789
rect 8386 25780 8392 25792
rect 8444 25780 8450 25832
rect 8481 25823 8539 25829
rect 8481 25789 8493 25823
rect 8527 25789 8539 25823
rect 9508 25820 9536 25851
rect 11974 25848 11980 25900
rect 12032 25888 12038 25900
rect 12069 25891 12127 25897
rect 12069 25888 12081 25891
rect 12032 25860 12081 25888
rect 12032 25848 12038 25860
rect 12069 25857 12081 25860
rect 12115 25857 12127 25891
rect 12069 25851 12127 25857
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25857 12587 25891
rect 12529 25851 12587 25857
rect 10134 25820 10140 25832
rect 9508 25792 10140 25820
rect 8481 25783 8539 25789
rect 7929 25755 7987 25761
rect 7929 25752 7941 25755
rect 6880 25724 7328 25752
rect 7392 25724 7941 25752
rect 6880 25712 6886 25724
rect 3421 25687 3479 25693
rect 3421 25653 3433 25687
rect 3467 25684 3479 25687
rect 4062 25684 4068 25696
rect 3467 25656 4068 25684
rect 3467 25653 3479 25656
rect 3421 25647 3479 25653
rect 4062 25644 4068 25656
rect 4120 25644 4126 25696
rect 7098 25644 7104 25696
rect 7156 25684 7162 25696
rect 7193 25687 7251 25693
rect 7193 25684 7205 25687
rect 7156 25656 7205 25684
rect 7156 25644 7162 25656
rect 7193 25653 7205 25656
rect 7239 25653 7251 25687
rect 7300 25684 7328 25724
rect 7929 25721 7941 25724
rect 7975 25721 7987 25755
rect 7929 25715 7987 25721
rect 8110 25712 8116 25764
rect 8168 25752 8174 25764
rect 8496 25752 8524 25783
rect 10134 25780 10140 25792
rect 10192 25780 10198 25832
rect 10413 25823 10471 25829
rect 10413 25789 10425 25823
rect 10459 25820 10471 25823
rect 10502 25820 10508 25832
rect 10459 25792 10508 25820
rect 10459 25789 10471 25792
rect 10413 25783 10471 25789
rect 10502 25780 10508 25792
rect 10560 25780 10566 25832
rect 8168 25724 9168 25752
rect 8168 25712 8174 25724
rect 9140 25693 9168 25724
rect 9766 25712 9772 25764
rect 9824 25712 9830 25764
rect 12544 25752 12572 25851
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 12805 25891 12863 25897
rect 12805 25857 12817 25891
rect 12851 25888 12863 25891
rect 13188 25888 13216 25984
rect 12851 25860 13216 25888
rect 13648 25888 13676 25987
rect 15838 25984 15844 26036
rect 15896 26024 15902 26036
rect 15933 26027 15991 26033
rect 15933 26024 15945 26027
rect 15896 25996 15945 26024
rect 15896 25984 15902 25996
rect 15933 25993 15945 25996
rect 15979 25993 15991 26027
rect 15933 25987 15991 25993
rect 17954 25984 17960 26036
rect 18012 26024 18018 26036
rect 19150 26024 19156 26036
rect 18012 25996 19156 26024
rect 18012 25984 18018 25996
rect 19150 25984 19156 25996
rect 19208 26024 19214 26036
rect 20806 26024 20812 26036
rect 19208 25996 19748 26024
rect 19208 25984 19214 25996
rect 15197 25959 15255 25965
rect 14384 25928 15056 25956
rect 14384 25900 14412 25928
rect 13949 25891 14007 25897
rect 13949 25888 13961 25891
rect 13648 25860 13961 25888
rect 12851 25857 12863 25860
rect 12805 25851 12863 25857
rect 13949 25857 13961 25860
rect 13995 25857 14007 25891
rect 13949 25851 14007 25857
rect 14090 25848 14096 25900
rect 14148 25848 14154 25900
rect 14185 25891 14243 25897
rect 14185 25857 14197 25891
rect 14231 25888 14243 25891
rect 14274 25888 14280 25900
rect 14231 25860 14280 25888
rect 14231 25857 14243 25860
rect 14185 25851 14243 25857
rect 14274 25848 14280 25860
rect 14332 25848 14338 25900
rect 14366 25848 14372 25900
rect 14424 25848 14430 25900
rect 14918 25848 14924 25900
rect 14976 25848 14982 25900
rect 15028 25888 15056 25928
rect 15197 25925 15209 25959
rect 15243 25956 15255 25959
rect 17310 25956 17316 25968
rect 15243 25928 17316 25956
rect 15243 25925 15255 25928
rect 15197 25919 15255 25925
rect 15289 25891 15347 25897
rect 15289 25888 15301 25891
rect 15028 25860 15301 25888
rect 15289 25857 15301 25860
rect 15335 25857 15347 25891
rect 15289 25851 15347 25857
rect 15473 25891 15531 25897
rect 15473 25857 15485 25891
rect 15519 25888 15531 25891
rect 15654 25888 15660 25900
rect 15519 25860 15660 25888
rect 15519 25857 15531 25860
rect 15473 25851 15531 25857
rect 13078 25780 13084 25832
rect 13136 25780 13142 25832
rect 13173 25823 13231 25829
rect 13173 25789 13185 25823
rect 13219 25820 13231 25823
rect 13814 25820 13820 25832
rect 13219 25792 13820 25820
rect 13219 25789 13231 25792
rect 13173 25783 13231 25789
rect 13814 25780 13820 25792
rect 13872 25780 13878 25832
rect 14458 25780 14464 25832
rect 14516 25820 14522 25832
rect 15013 25823 15071 25829
rect 15013 25820 15025 25823
rect 14516 25792 15025 25820
rect 14516 25780 14522 25792
rect 15013 25789 15025 25792
rect 15059 25789 15071 25823
rect 15013 25783 15071 25789
rect 15194 25780 15200 25832
rect 15252 25780 15258 25832
rect 15304 25820 15332 25851
rect 15654 25848 15660 25860
rect 15712 25848 15718 25900
rect 15764 25897 15792 25928
rect 17310 25916 17316 25928
rect 17368 25916 17374 25968
rect 17862 25956 17868 25968
rect 17604 25928 17868 25956
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25857 15807 25891
rect 15749 25851 15807 25857
rect 16206 25848 16212 25900
rect 16264 25848 16270 25900
rect 17604 25897 17632 25928
rect 17862 25916 17868 25928
rect 17920 25956 17926 25968
rect 17920 25928 18460 25956
rect 17920 25916 17926 25928
rect 17589 25891 17647 25897
rect 17589 25857 17601 25891
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 17770 25848 17776 25900
rect 17828 25848 17834 25900
rect 18138 25848 18144 25900
rect 18196 25888 18202 25900
rect 18432 25897 18460 25928
rect 18708 25928 19656 25956
rect 18708 25900 18736 25928
rect 18233 25891 18291 25897
rect 18233 25888 18245 25891
rect 18196 25860 18245 25888
rect 18196 25848 18202 25860
rect 18233 25857 18245 25860
rect 18279 25857 18291 25891
rect 18233 25851 18291 25857
rect 18417 25891 18475 25897
rect 18417 25857 18429 25891
rect 18463 25857 18475 25891
rect 18417 25851 18475 25857
rect 18506 25848 18512 25900
rect 18564 25848 18570 25900
rect 18690 25848 18696 25900
rect 18748 25848 18754 25900
rect 18874 25848 18880 25900
rect 18932 25848 18938 25900
rect 19058 25848 19064 25900
rect 19116 25848 19122 25900
rect 19337 25891 19395 25897
rect 19337 25888 19349 25891
rect 19168 25860 19349 25888
rect 16117 25823 16175 25829
rect 16117 25820 16129 25823
rect 15304 25792 16129 25820
rect 16117 25789 16129 25792
rect 16163 25789 16175 25823
rect 16117 25783 16175 25789
rect 18322 25780 18328 25832
rect 18380 25820 18386 25832
rect 18785 25823 18843 25829
rect 18785 25820 18797 25823
rect 18380 25792 18797 25820
rect 18380 25780 18386 25792
rect 18785 25789 18797 25792
rect 18831 25789 18843 25823
rect 18785 25783 18843 25789
rect 13630 25752 13636 25764
rect 12544 25724 13636 25752
rect 13630 25712 13636 25724
rect 13688 25712 13694 25764
rect 18598 25712 18604 25764
rect 18656 25752 18662 25764
rect 19168 25752 19196 25860
rect 19337 25857 19349 25860
rect 19383 25857 19395 25891
rect 19337 25851 19395 25857
rect 19518 25848 19524 25900
rect 19576 25848 19582 25900
rect 19628 25897 19656 25928
rect 19720 25897 19748 25996
rect 20180 25996 20812 26024
rect 20180 25965 20208 25996
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 20916 25996 21588 26024
rect 20916 25965 20944 25996
rect 20165 25959 20223 25965
rect 20165 25925 20177 25959
rect 20211 25925 20223 25959
rect 20165 25919 20223 25925
rect 20901 25959 20959 25965
rect 20901 25925 20913 25959
rect 20947 25925 20959 25959
rect 20901 25919 20959 25925
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 19705 25891 19763 25897
rect 19705 25857 19717 25891
rect 19751 25857 19763 25891
rect 19705 25851 19763 25857
rect 20346 25848 20352 25900
rect 20404 25888 20410 25900
rect 20533 25891 20591 25897
rect 20533 25888 20545 25891
rect 20404 25860 20545 25888
rect 20404 25848 20410 25860
rect 20533 25857 20545 25860
rect 20579 25857 20591 25891
rect 20533 25851 20591 25857
rect 20622 25848 20628 25900
rect 20680 25848 20686 25900
rect 20806 25848 20812 25900
rect 20864 25888 20870 25900
rect 20916 25888 20944 25919
rect 21266 25916 21272 25968
rect 21324 25916 21330 25968
rect 21560 25897 21588 25996
rect 24026 25984 24032 26036
rect 24084 26024 24090 26036
rect 24213 26027 24271 26033
rect 24213 26024 24225 26027
rect 24084 25996 24225 26024
rect 24084 25984 24090 25996
rect 24213 25993 24225 25996
rect 24259 25993 24271 26027
rect 24213 25987 24271 25993
rect 25409 26027 25467 26033
rect 25409 25993 25421 26027
rect 25455 26024 25467 26027
rect 26050 26024 26056 26036
rect 25455 25996 26056 26024
rect 25455 25993 25467 25996
rect 25409 25987 25467 25993
rect 21634 25916 21640 25968
rect 21692 25956 21698 25968
rect 21821 25959 21879 25965
rect 21821 25956 21833 25959
rect 21692 25928 21833 25956
rect 21692 25916 21698 25928
rect 21821 25925 21833 25928
rect 21867 25925 21879 25959
rect 21821 25919 21879 25925
rect 21085 25891 21143 25897
rect 21085 25888 21097 25891
rect 20864 25860 20944 25888
rect 21008 25860 21097 25888
rect 20864 25848 20870 25860
rect 19242 25780 19248 25832
rect 19300 25820 19306 25832
rect 20257 25823 20315 25829
rect 20257 25820 20269 25823
rect 19300 25792 20269 25820
rect 19300 25780 19306 25792
rect 20257 25789 20269 25792
rect 20303 25789 20315 25823
rect 20640 25820 20668 25848
rect 21008 25820 21036 25860
rect 21085 25857 21097 25860
rect 21131 25857 21143 25891
rect 21361 25891 21419 25897
rect 21361 25888 21373 25891
rect 21085 25851 21143 25857
rect 21284 25860 21373 25888
rect 20640 25792 21036 25820
rect 20257 25783 20315 25789
rect 18656 25724 19196 25752
rect 20809 25755 20867 25761
rect 18656 25712 18662 25724
rect 20809 25721 20821 25755
rect 20855 25752 20867 25755
rect 20898 25752 20904 25764
rect 20855 25724 20904 25752
rect 20855 25721 20867 25724
rect 20809 25715 20867 25721
rect 20898 25712 20904 25724
rect 20956 25712 20962 25764
rect 8941 25687 8999 25693
rect 8941 25684 8953 25687
rect 7300 25656 8953 25684
rect 7193 25647 7251 25653
rect 8941 25653 8953 25656
rect 8987 25653 8999 25687
rect 8941 25647 8999 25653
rect 9125 25687 9183 25693
rect 9125 25653 9137 25687
rect 9171 25653 9183 25687
rect 9125 25647 9183 25653
rect 10042 25644 10048 25696
rect 10100 25684 10106 25696
rect 10505 25687 10563 25693
rect 10505 25684 10517 25687
rect 10100 25656 10517 25684
rect 10100 25644 10106 25656
rect 10505 25653 10517 25656
rect 10551 25653 10563 25687
rect 10505 25647 10563 25653
rect 10689 25687 10747 25693
rect 10689 25653 10701 25687
rect 10735 25684 10747 25687
rect 11146 25684 11152 25696
rect 10735 25656 11152 25684
rect 10735 25653 10747 25656
rect 10689 25647 10747 25653
rect 11146 25644 11152 25656
rect 11204 25644 11210 25696
rect 12345 25687 12403 25693
rect 12345 25653 12357 25687
rect 12391 25684 12403 25687
rect 13262 25684 13268 25696
rect 12391 25656 13268 25684
rect 12391 25653 12403 25656
rect 12345 25647 12403 25653
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 13538 25644 13544 25696
rect 13596 25684 13602 25696
rect 13817 25687 13875 25693
rect 13817 25684 13829 25687
rect 13596 25656 13829 25684
rect 13596 25644 13602 25656
rect 13817 25653 13829 25656
rect 13863 25684 13875 25687
rect 17589 25687 17647 25693
rect 17589 25684 17601 25687
rect 13863 25656 17601 25684
rect 13863 25653 13875 25656
rect 13817 25647 13875 25653
rect 17589 25653 17601 25656
rect 17635 25684 17647 25687
rect 17678 25684 17684 25696
rect 17635 25656 17684 25684
rect 17635 25653 17647 25656
rect 17589 25647 17647 25653
rect 17678 25644 17684 25656
rect 17736 25644 17742 25696
rect 17957 25687 18015 25693
rect 17957 25653 17969 25687
rect 18003 25684 18015 25687
rect 18230 25684 18236 25696
rect 18003 25656 18236 25684
rect 18003 25653 18015 25656
rect 17957 25647 18015 25653
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 18417 25687 18475 25693
rect 18417 25653 18429 25687
rect 18463 25684 18475 25687
rect 18966 25684 18972 25696
rect 18463 25656 18972 25684
rect 18463 25653 18475 25656
rect 18417 25647 18475 25653
rect 18966 25644 18972 25656
rect 19024 25644 19030 25696
rect 19245 25687 19303 25693
rect 19245 25653 19257 25687
rect 19291 25684 19303 25687
rect 19886 25684 19892 25696
rect 19291 25656 19892 25684
rect 19291 25653 19303 25656
rect 19245 25647 19303 25653
rect 19886 25644 19892 25656
rect 19944 25644 19950 25696
rect 19981 25687 20039 25693
rect 19981 25653 19993 25687
rect 20027 25684 20039 25687
rect 21284 25684 21312 25860
rect 21361 25857 21373 25860
rect 21407 25857 21419 25891
rect 21361 25851 21419 25857
rect 21545 25891 21603 25897
rect 21545 25857 21557 25891
rect 21591 25857 21603 25891
rect 21545 25851 21603 25857
rect 22278 25848 22284 25900
rect 22336 25848 22342 25900
rect 22554 25848 22560 25900
rect 22612 25888 22618 25900
rect 23106 25897 23112 25900
rect 22833 25891 22891 25897
rect 22833 25888 22845 25891
rect 22612 25860 22845 25888
rect 22612 25848 22618 25860
rect 22833 25857 22845 25860
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23100 25851 23112 25897
rect 23106 25848 23112 25851
rect 23164 25848 23170 25900
rect 24228 25888 24256 25987
rect 26050 25984 26056 25996
rect 26108 25984 26114 26036
rect 29178 26024 29184 26036
rect 28368 25996 29184 26024
rect 24302 25916 24308 25968
rect 24360 25956 24366 25968
rect 28368 25965 28396 25996
rect 29178 25984 29184 25996
rect 29236 25984 29242 26036
rect 29822 25984 29828 26036
rect 29880 26024 29886 26036
rect 30282 26024 30288 26036
rect 29880 25996 30288 26024
rect 29880 25984 29886 25996
rect 30282 25984 30288 25996
rect 30340 25984 30346 26036
rect 31481 26027 31539 26033
rect 31481 25993 31493 26027
rect 31527 26024 31539 26027
rect 31662 26024 31668 26036
rect 31527 25996 31668 26024
rect 31527 25993 31539 25996
rect 31481 25987 31539 25993
rect 31662 25984 31668 25996
rect 31720 26024 31726 26036
rect 31849 26027 31907 26033
rect 31849 26024 31861 26027
rect 31720 25996 31861 26024
rect 31720 25984 31726 25996
rect 31849 25993 31861 25996
rect 31895 25993 31907 26027
rect 33505 26027 33563 26033
rect 31849 25987 31907 25993
rect 32416 25996 33364 26024
rect 32416 25968 32444 25996
rect 25041 25959 25099 25965
rect 25041 25956 25053 25959
rect 24360 25928 25053 25956
rect 24360 25916 24366 25928
rect 25041 25925 25053 25928
rect 25087 25925 25099 25959
rect 25041 25919 25099 25925
rect 28353 25959 28411 25965
rect 28353 25925 28365 25959
rect 28399 25925 28411 25959
rect 29638 25956 29644 25968
rect 29578 25928 29644 25956
rect 28353 25919 28411 25925
rect 29638 25916 29644 25928
rect 29696 25916 29702 25968
rect 32398 25916 32404 25968
rect 32456 25916 32462 25968
rect 32784 25928 33272 25956
rect 24857 25891 24915 25897
rect 24857 25888 24869 25891
rect 24228 25860 24869 25888
rect 24857 25857 24869 25860
rect 24903 25857 24915 25891
rect 24857 25851 24915 25857
rect 25222 25848 25228 25900
rect 25280 25848 25286 25900
rect 26326 25848 26332 25900
rect 26384 25888 26390 25900
rect 27798 25888 27804 25900
rect 26384 25860 27804 25888
rect 26384 25848 26390 25860
rect 27798 25848 27804 25860
rect 27856 25848 27862 25900
rect 27890 25848 27896 25900
rect 27948 25848 27954 25900
rect 29822 25848 29828 25900
rect 29880 25888 29886 25900
rect 30009 25891 30067 25897
rect 30009 25888 30021 25891
rect 29880 25860 30021 25888
rect 29880 25848 29886 25860
rect 30009 25857 30021 25860
rect 30055 25857 30067 25891
rect 30009 25851 30067 25857
rect 31110 25848 31116 25900
rect 31168 25888 31174 25900
rect 31570 25888 31576 25900
rect 31168 25860 31576 25888
rect 31168 25848 31174 25860
rect 31570 25848 31576 25860
rect 31628 25888 31634 25900
rect 32125 25891 32183 25897
rect 32125 25888 32137 25891
rect 31628 25860 32137 25888
rect 31628 25848 31634 25860
rect 32125 25857 32137 25860
rect 32171 25857 32183 25891
rect 32125 25851 32183 25857
rect 32306 25848 32312 25900
rect 32364 25848 32370 25900
rect 32784 25897 32812 25928
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25888 32551 25891
rect 32769 25891 32827 25897
rect 32539 25860 32628 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 22186 25780 22192 25832
rect 22244 25780 22250 25832
rect 25866 25780 25872 25832
rect 25924 25820 25930 25832
rect 27617 25823 27675 25829
rect 27617 25820 27629 25823
rect 25924 25792 27629 25820
rect 25924 25780 25930 25792
rect 27617 25789 27629 25792
rect 27663 25820 27675 25823
rect 27706 25820 27712 25832
rect 27663 25792 27712 25820
rect 27663 25789 27675 25792
rect 27617 25783 27675 25789
rect 27706 25780 27712 25792
rect 27764 25780 27770 25832
rect 28074 25780 28080 25832
rect 28132 25780 28138 25832
rect 26878 25752 26884 25764
rect 23768 25724 26884 25752
rect 20027 25656 21312 25684
rect 20027 25653 20039 25656
rect 19981 25647 20039 25653
rect 21358 25644 21364 25696
rect 21416 25644 21422 25696
rect 22094 25644 22100 25696
rect 22152 25644 22158 25696
rect 22465 25687 22523 25693
rect 22465 25653 22477 25687
rect 22511 25684 22523 25687
rect 22646 25684 22652 25696
rect 22511 25656 22652 25684
rect 22511 25653 22523 25656
rect 22465 25647 22523 25653
rect 22646 25644 22652 25656
rect 22704 25644 22710 25696
rect 22830 25644 22836 25696
rect 22888 25684 22894 25696
rect 23768 25684 23796 25724
rect 26878 25712 26884 25724
rect 26936 25712 26942 25764
rect 27522 25712 27528 25764
rect 27580 25752 27586 25764
rect 28092 25752 28120 25780
rect 27580 25724 28120 25752
rect 27580 25712 27586 25724
rect 22888 25656 23796 25684
rect 22888 25644 22894 25656
rect 24302 25644 24308 25696
rect 24360 25644 24366 25696
rect 27709 25687 27767 25693
rect 27709 25653 27721 25687
rect 27755 25684 27767 25687
rect 29086 25684 29092 25696
rect 27755 25656 29092 25684
rect 27755 25653 27767 25656
rect 27709 25647 27767 25653
rect 29086 25644 29092 25656
rect 29144 25644 29150 25696
rect 32600 25684 32628 25860
rect 32769 25857 32781 25891
rect 32815 25857 32827 25891
rect 32769 25851 32827 25857
rect 32950 25848 32956 25900
rect 33008 25848 33014 25900
rect 33045 25823 33103 25829
rect 33045 25789 33057 25823
rect 33091 25789 33103 25823
rect 33045 25783 33103 25789
rect 32677 25755 32735 25761
rect 32677 25721 32689 25755
rect 32723 25752 32735 25755
rect 33060 25752 33088 25783
rect 33134 25780 33140 25832
rect 33192 25780 33198 25832
rect 32723 25724 33088 25752
rect 33244 25752 33272 25928
rect 33336 25897 33364 25996
rect 33505 25993 33517 26027
rect 33551 26024 33563 26027
rect 35713 26027 35771 26033
rect 33551 25996 34468 26024
rect 33551 25993 33563 25996
rect 33505 25987 33563 25993
rect 33796 25928 34376 25956
rect 33321 25891 33379 25897
rect 33321 25857 33333 25891
rect 33367 25857 33379 25891
rect 33321 25851 33379 25857
rect 33594 25848 33600 25900
rect 33652 25848 33658 25900
rect 33796 25897 33824 25928
rect 34348 25900 34376 25928
rect 33781 25891 33839 25897
rect 33781 25857 33793 25891
rect 33827 25857 33839 25891
rect 33781 25851 33839 25857
rect 34149 25891 34207 25897
rect 34149 25857 34161 25891
rect 34195 25857 34207 25891
rect 34149 25851 34207 25857
rect 33612 25820 33640 25848
rect 34164 25820 34192 25851
rect 34330 25848 34336 25900
rect 34388 25848 34394 25900
rect 34440 25888 34468 25996
rect 35713 25993 35725 26027
rect 35759 26024 35771 26027
rect 35986 26024 35992 26036
rect 35759 25996 35992 26024
rect 35759 25993 35771 25996
rect 35713 25987 35771 25993
rect 35986 25984 35992 25996
rect 36044 25984 36050 26036
rect 36078 25984 36084 26036
rect 36136 26024 36142 26036
rect 36265 26027 36323 26033
rect 36265 26024 36277 26027
rect 36136 25996 36277 26024
rect 36136 25984 36142 25996
rect 36265 25993 36277 25996
rect 36311 25993 36323 26027
rect 36265 25987 36323 25993
rect 34790 25916 34796 25968
rect 34848 25956 34854 25968
rect 34848 25928 36124 25956
rect 34848 25916 34854 25928
rect 35069 25891 35127 25897
rect 35069 25888 35081 25891
rect 34440 25860 35081 25888
rect 35069 25857 35081 25860
rect 35115 25857 35127 25891
rect 35069 25851 35127 25857
rect 35161 25891 35219 25897
rect 35161 25857 35173 25891
rect 35207 25857 35219 25891
rect 35161 25851 35219 25857
rect 35345 25891 35403 25897
rect 35345 25857 35357 25891
rect 35391 25857 35403 25891
rect 35345 25851 35403 25857
rect 33612 25792 34192 25820
rect 34241 25823 34299 25829
rect 34241 25789 34253 25823
rect 34287 25820 34299 25823
rect 35176 25820 35204 25851
rect 34287 25792 35204 25820
rect 34287 25789 34299 25792
rect 34241 25783 34299 25789
rect 33689 25755 33747 25761
rect 33689 25752 33701 25755
rect 33244 25724 33701 25752
rect 32723 25721 32735 25724
rect 32677 25715 32735 25721
rect 33689 25721 33701 25724
rect 33735 25721 33747 25755
rect 35360 25752 35388 25851
rect 35434 25848 35440 25900
rect 35492 25848 35498 25900
rect 35544 25897 35572 25928
rect 36096 25897 36124 25928
rect 37458 25916 37464 25968
rect 37516 25956 37522 25968
rect 37645 25959 37703 25965
rect 37645 25956 37657 25959
rect 37516 25928 37657 25956
rect 37516 25916 37522 25928
rect 37645 25925 37657 25928
rect 37691 25925 37703 25959
rect 37645 25919 37703 25925
rect 35529 25891 35587 25897
rect 35529 25857 35541 25891
rect 35575 25857 35587 25891
rect 35529 25851 35587 25857
rect 35805 25891 35863 25897
rect 35805 25857 35817 25891
rect 35851 25857 35863 25891
rect 35805 25851 35863 25857
rect 35897 25891 35955 25897
rect 35897 25857 35909 25891
rect 35943 25857 35955 25891
rect 35897 25851 35955 25857
rect 36081 25891 36139 25897
rect 36081 25857 36093 25891
rect 36127 25857 36139 25891
rect 36081 25851 36139 25857
rect 35452 25820 35480 25848
rect 35820 25820 35848 25851
rect 35452 25792 35848 25820
rect 35912 25752 35940 25851
rect 37826 25848 37832 25900
rect 37884 25848 37890 25900
rect 37461 25823 37519 25829
rect 37461 25789 37473 25823
rect 37507 25820 37519 25823
rect 37550 25820 37556 25832
rect 37507 25792 37556 25820
rect 37507 25789 37519 25792
rect 37461 25783 37519 25789
rect 37550 25780 37556 25792
rect 37608 25780 37614 25832
rect 35986 25752 35992 25764
rect 35360 25724 35992 25752
rect 33689 25715 33747 25721
rect 35986 25712 35992 25724
rect 36044 25712 36050 25764
rect 33134 25684 33140 25696
rect 32600 25656 33140 25684
rect 33134 25644 33140 25656
rect 33192 25644 33198 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 3237 25483 3295 25489
rect 3237 25449 3249 25483
rect 3283 25480 3295 25483
rect 3326 25480 3332 25492
rect 3283 25452 3332 25480
rect 3283 25449 3295 25452
rect 3237 25443 3295 25449
rect 3326 25440 3332 25452
rect 3384 25440 3390 25492
rect 3421 25483 3479 25489
rect 3421 25449 3433 25483
rect 3467 25449 3479 25483
rect 3421 25443 3479 25449
rect 3142 25372 3148 25424
rect 3200 25412 3206 25424
rect 3436 25412 3464 25443
rect 6086 25440 6092 25492
rect 6144 25440 6150 25492
rect 7006 25440 7012 25492
rect 7064 25480 7070 25492
rect 7101 25483 7159 25489
rect 7101 25480 7113 25483
rect 7064 25452 7113 25480
rect 7064 25440 7070 25452
rect 7101 25449 7113 25452
rect 7147 25449 7159 25483
rect 7101 25443 7159 25449
rect 8110 25440 8116 25492
rect 8168 25480 8174 25492
rect 8297 25483 8355 25489
rect 8297 25480 8309 25483
rect 8168 25452 8309 25480
rect 8168 25440 8174 25452
rect 8297 25449 8309 25452
rect 8343 25449 8355 25483
rect 8297 25443 8355 25449
rect 9214 25440 9220 25492
rect 9272 25480 9278 25492
rect 11146 25480 11152 25492
rect 9272 25452 11152 25480
rect 9272 25440 9278 25452
rect 11146 25440 11152 25452
rect 11204 25440 11210 25492
rect 12805 25483 12863 25489
rect 12805 25449 12817 25483
rect 12851 25480 12863 25483
rect 13170 25480 13176 25492
rect 12851 25452 13176 25480
rect 12851 25449 12863 25452
rect 12805 25443 12863 25449
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 13633 25483 13691 25489
rect 13633 25449 13645 25483
rect 13679 25480 13691 25483
rect 14090 25480 14096 25492
rect 13679 25452 14096 25480
rect 13679 25449 13691 25452
rect 13633 25443 13691 25449
rect 3200 25384 3464 25412
rect 3200 25372 3206 25384
rect 5994 25372 6000 25424
rect 6052 25412 6058 25424
rect 8846 25412 8852 25424
rect 6052 25384 8852 25412
rect 6052 25372 6058 25384
rect 8846 25372 8852 25384
rect 8904 25412 8910 25424
rect 9861 25415 9919 25421
rect 9861 25412 9873 25415
rect 8904 25384 9873 25412
rect 8904 25372 8910 25384
rect 9861 25381 9873 25384
rect 9907 25381 9919 25415
rect 13648 25412 13676 25443
rect 14090 25440 14096 25452
rect 14148 25440 14154 25492
rect 14826 25440 14832 25492
rect 14884 25480 14890 25492
rect 15197 25483 15255 25489
rect 15197 25480 15209 25483
rect 14884 25452 15209 25480
rect 14884 25440 14890 25452
rect 15197 25449 15209 25452
rect 15243 25480 15255 25483
rect 15378 25480 15384 25492
rect 15243 25452 15384 25480
rect 15243 25449 15255 25452
rect 15197 25443 15255 25449
rect 15378 25440 15384 25452
rect 15436 25440 15442 25492
rect 15562 25440 15568 25492
rect 15620 25440 15626 25492
rect 15654 25440 15660 25492
rect 15712 25440 15718 25492
rect 18233 25483 18291 25489
rect 18233 25449 18245 25483
rect 18279 25480 18291 25483
rect 18506 25480 18512 25492
rect 18279 25452 18512 25480
rect 18279 25449 18291 25452
rect 18233 25443 18291 25449
rect 18506 25440 18512 25452
rect 18564 25440 18570 25492
rect 20070 25440 20076 25492
rect 20128 25440 20134 25492
rect 20533 25483 20591 25489
rect 20533 25449 20545 25483
rect 20579 25480 20591 25483
rect 21450 25480 21456 25492
rect 20579 25452 21456 25480
rect 20579 25449 20591 25452
rect 20533 25443 20591 25449
rect 21450 25440 21456 25452
rect 21508 25440 21514 25492
rect 21818 25440 21824 25492
rect 21876 25480 21882 25492
rect 21913 25483 21971 25489
rect 21913 25480 21925 25483
rect 21876 25452 21925 25480
rect 21876 25440 21882 25452
rect 21913 25449 21925 25452
rect 21959 25449 21971 25483
rect 21913 25443 21971 25449
rect 23106 25440 23112 25492
rect 23164 25480 23170 25492
rect 23293 25483 23351 25489
rect 23293 25480 23305 25483
rect 23164 25452 23305 25480
rect 23164 25440 23170 25452
rect 23293 25449 23305 25452
rect 23339 25449 23351 25483
rect 23293 25443 23351 25449
rect 24949 25483 25007 25489
rect 24949 25449 24961 25483
rect 24995 25480 25007 25483
rect 25682 25480 25688 25492
rect 24995 25452 25688 25480
rect 24995 25449 25007 25452
rect 24949 25443 25007 25449
rect 25682 25440 25688 25452
rect 25740 25440 25746 25492
rect 25869 25483 25927 25489
rect 25869 25449 25881 25483
rect 25915 25480 25927 25483
rect 26970 25480 26976 25492
rect 25915 25452 26976 25480
rect 25915 25449 25927 25452
rect 25869 25443 25927 25449
rect 26970 25440 26976 25452
rect 27028 25440 27034 25492
rect 31113 25483 31171 25489
rect 31113 25449 31125 25483
rect 31159 25480 31171 25483
rect 31159 25452 31524 25480
rect 31159 25449 31171 25452
rect 31113 25443 31171 25449
rect 9861 25375 9919 25381
rect 13464 25384 13676 25412
rect 1394 25304 1400 25356
rect 1452 25344 1458 25356
rect 2682 25344 2688 25356
rect 1452 25316 2688 25344
rect 1452 25304 1458 25316
rect 2682 25304 2688 25316
rect 2740 25344 2746 25356
rect 3789 25347 3847 25353
rect 3789 25344 3801 25347
rect 2740 25316 3801 25344
rect 2740 25304 2746 25316
rect 3789 25313 3801 25316
rect 3835 25313 3847 25347
rect 3789 25307 3847 25313
rect 4062 25304 4068 25356
rect 4120 25304 4126 25356
rect 8386 25344 8392 25356
rect 7944 25316 8392 25344
rect 3050 25276 3056 25288
rect 2806 25248 3056 25276
rect 3050 25236 3056 25248
rect 3108 25276 3114 25288
rect 3108 25248 3740 25276
rect 3108 25236 3114 25248
rect 1673 25211 1731 25217
rect 1673 25177 1685 25211
rect 1719 25208 1731 25211
rect 1762 25208 1768 25220
rect 1719 25180 1768 25208
rect 1719 25177 1731 25180
rect 1673 25171 1731 25177
rect 1762 25168 1768 25180
rect 1820 25168 1826 25220
rect 2958 25168 2964 25220
rect 3016 25208 3022 25220
rect 3389 25211 3447 25217
rect 3389 25208 3401 25211
rect 3016 25180 3401 25208
rect 3016 25168 3022 25180
rect 3389 25177 3401 25180
rect 3435 25177 3447 25211
rect 3389 25171 3447 25177
rect 3605 25211 3663 25217
rect 3605 25177 3617 25211
rect 3651 25177 3663 25211
rect 3712 25208 3740 25248
rect 5626 25236 5632 25288
rect 5684 25236 5690 25288
rect 5813 25279 5871 25285
rect 5813 25245 5825 25279
rect 5859 25276 5871 25279
rect 6822 25276 6828 25288
rect 5859 25248 5948 25276
rect 5859 25245 5871 25248
rect 5813 25239 5871 25245
rect 3712 25180 4554 25208
rect 3605 25171 3663 25177
rect 3142 25100 3148 25152
rect 3200 25100 3206 25152
rect 3620 25140 3648 25171
rect 5920 25152 5948 25248
rect 6196 25248 6828 25276
rect 6196 25220 6224 25248
rect 6822 25236 6828 25248
rect 6880 25276 6886 25288
rect 6917 25279 6975 25285
rect 6917 25276 6929 25279
rect 6880 25248 6929 25276
rect 6880 25236 6886 25248
rect 6917 25245 6929 25248
rect 6963 25245 6975 25279
rect 6917 25239 6975 25245
rect 7098 25236 7104 25288
rect 7156 25236 7162 25288
rect 7944 25285 7972 25316
rect 8386 25304 8392 25316
rect 8444 25344 8450 25356
rect 13464 25353 13492 25384
rect 14918 25372 14924 25424
rect 14976 25412 14982 25424
rect 16025 25415 16083 25421
rect 16025 25412 16037 25415
rect 14976 25384 16037 25412
rect 14976 25372 14982 25384
rect 16025 25381 16037 25384
rect 16071 25381 16083 25415
rect 16025 25375 16083 25381
rect 18138 25372 18144 25424
rect 18196 25412 18202 25424
rect 21358 25412 21364 25424
rect 18196 25384 18552 25412
rect 18196 25372 18202 25384
rect 13449 25347 13507 25353
rect 8444 25316 9536 25344
rect 8444 25304 8450 25316
rect 9508 25288 9536 25316
rect 13449 25313 13461 25347
rect 13495 25313 13507 25347
rect 15286 25344 15292 25356
rect 13449 25307 13507 25313
rect 14752 25316 15292 25344
rect 7837 25279 7895 25285
rect 7837 25245 7849 25279
rect 7883 25245 7895 25279
rect 7837 25239 7895 25245
rect 7929 25279 7987 25285
rect 7929 25245 7941 25279
rect 7975 25245 7987 25279
rect 7929 25239 7987 25245
rect 8297 25279 8355 25285
rect 8297 25245 8309 25279
rect 8343 25276 8355 25279
rect 9214 25276 9220 25288
rect 8343 25248 9220 25276
rect 8343 25245 8355 25248
rect 8297 25239 8355 25245
rect 6073 25211 6131 25217
rect 6073 25177 6085 25211
rect 6119 25208 6131 25211
rect 6178 25208 6184 25220
rect 6119 25180 6184 25208
rect 6119 25177 6131 25180
rect 6073 25171 6131 25177
rect 6178 25168 6184 25180
rect 6236 25168 6242 25220
rect 6273 25211 6331 25217
rect 6273 25177 6285 25211
rect 6319 25208 6331 25211
rect 6362 25208 6368 25220
rect 6319 25180 6368 25208
rect 6319 25177 6331 25180
rect 6273 25171 6331 25177
rect 6362 25168 6368 25180
rect 6420 25208 6426 25220
rect 7852 25208 7880 25239
rect 9214 25236 9220 25248
rect 9272 25236 9278 25288
rect 9490 25236 9496 25288
rect 9548 25276 9554 25288
rect 10229 25279 10287 25285
rect 10229 25276 10241 25279
rect 9548 25248 10241 25276
rect 9548 25236 9554 25248
rect 10229 25245 10241 25248
rect 10275 25245 10287 25279
rect 10229 25239 10287 25245
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25276 10471 25279
rect 12066 25276 12072 25288
rect 10459 25248 12072 25276
rect 10459 25245 10471 25248
rect 10413 25239 10471 25245
rect 12066 25236 12072 25248
rect 12124 25236 12130 25288
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25276 12403 25279
rect 12529 25279 12587 25285
rect 12529 25276 12541 25279
rect 12391 25248 12541 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 12529 25245 12541 25248
rect 12575 25276 12587 25279
rect 12802 25276 12808 25288
rect 12575 25248 12808 25276
rect 12575 25245 12587 25248
rect 12529 25239 12587 25245
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 12986 25236 12992 25288
rect 13044 25236 13050 25288
rect 13262 25236 13268 25288
rect 13320 25285 13326 25288
rect 13320 25279 13349 25285
rect 13337 25245 13349 25279
rect 13320 25239 13349 25245
rect 13725 25279 13783 25285
rect 13725 25245 13737 25279
rect 13771 25276 13783 25279
rect 14752 25276 14780 25316
rect 15286 25304 15292 25316
rect 15344 25304 15350 25356
rect 15562 25304 15568 25356
rect 15620 25344 15626 25356
rect 15620 25316 15976 25344
rect 15620 25304 15626 25316
rect 13771 25248 14780 25276
rect 15105 25279 15163 25285
rect 13771 25245 13783 25248
rect 13725 25239 13783 25245
rect 15105 25245 15117 25279
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 13320 25236 13326 25239
rect 6420 25180 7880 25208
rect 6420 25168 6426 25180
rect 9030 25168 9036 25220
rect 9088 25208 9094 25220
rect 10045 25211 10103 25217
rect 10045 25208 10057 25211
rect 9088 25180 10057 25208
rect 9088 25168 9094 25180
rect 10045 25177 10057 25180
rect 10091 25208 10103 25211
rect 11146 25208 11152 25220
rect 10091 25180 11152 25208
rect 10091 25177 10103 25180
rect 10045 25171 10103 25177
rect 11146 25168 11152 25180
rect 11204 25168 11210 25220
rect 13081 25211 13139 25217
rect 13081 25177 13093 25211
rect 13127 25177 13139 25211
rect 13081 25171 13139 25177
rect 13173 25211 13231 25217
rect 13173 25177 13185 25211
rect 13219 25208 13231 25211
rect 14366 25208 14372 25220
rect 13219 25180 14372 25208
rect 13219 25177 13231 25180
rect 13173 25171 13231 25177
rect 4706 25140 4712 25152
rect 3620 25112 4712 25140
rect 4706 25100 4712 25112
rect 4764 25140 4770 25152
rect 5537 25143 5595 25149
rect 5537 25140 5549 25143
rect 4764 25112 5549 25140
rect 4764 25100 4770 25112
rect 5537 25109 5549 25112
rect 5583 25109 5595 25143
rect 5537 25103 5595 25109
rect 5718 25100 5724 25152
rect 5776 25100 5782 25152
rect 5902 25100 5908 25152
rect 5960 25100 5966 25152
rect 8478 25100 8484 25152
rect 8536 25100 8542 25152
rect 10318 25100 10324 25152
rect 10376 25100 10382 25152
rect 11054 25100 11060 25152
rect 11112 25140 11118 25152
rect 12618 25140 12624 25152
rect 11112 25112 12624 25140
rect 11112 25100 11118 25112
rect 12618 25100 12624 25112
rect 12676 25100 12682 25152
rect 13096 25140 13124 25171
rect 14366 25168 14372 25180
rect 14424 25168 14430 25220
rect 14734 25140 14740 25152
rect 13096 25112 14740 25140
rect 14734 25100 14740 25112
rect 14792 25100 14798 25152
rect 15120 25140 15148 25239
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 15657 25279 15715 25285
rect 15657 25276 15669 25279
rect 15436 25248 15669 25276
rect 15436 25236 15442 25248
rect 15657 25245 15669 25248
rect 15703 25245 15715 25279
rect 15657 25239 15715 25245
rect 15746 25236 15752 25288
rect 15804 25276 15810 25288
rect 15948 25285 15976 25316
rect 18322 25304 18328 25356
rect 18380 25304 18386 25356
rect 15841 25279 15899 25285
rect 15841 25276 15853 25279
rect 15804 25248 15853 25276
rect 15804 25236 15810 25248
rect 15841 25245 15853 25248
rect 15887 25245 15899 25279
rect 15841 25239 15899 25245
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25245 15991 25279
rect 15933 25239 15991 25245
rect 16298 25236 16304 25288
rect 16356 25236 16362 25288
rect 17954 25236 17960 25288
rect 18012 25276 18018 25288
rect 18049 25279 18107 25285
rect 18049 25276 18061 25279
rect 18012 25248 18061 25276
rect 18012 25236 18018 25248
rect 18049 25245 18061 25248
rect 18095 25245 18107 25279
rect 18049 25239 18107 25245
rect 18138 25236 18144 25288
rect 18196 25236 18202 25288
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 18417 25279 18475 25285
rect 18417 25276 18429 25279
rect 18288 25248 18429 25276
rect 18288 25236 18294 25248
rect 18417 25245 18429 25248
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 15470 25168 15476 25220
rect 15528 25208 15534 25220
rect 16025 25211 16083 25217
rect 16025 25208 16037 25211
rect 15528 25180 16037 25208
rect 15528 25168 15534 25180
rect 16025 25177 16037 25180
rect 16071 25177 16083 25211
rect 16025 25171 16083 25177
rect 16209 25211 16267 25217
rect 16209 25177 16221 25211
rect 16255 25208 16267 25211
rect 16390 25208 16396 25220
rect 16255 25180 16396 25208
rect 16255 25177 16267 25180
rect 16209 25171 16267 25177
rect 16390 25168 16396 25180
rect 16448 25168 16454 25220
rect 18524 25208 18552 25384
rect 20272 25384 21364 25412
rect 20272 25353 20300 25384
rect 21358 25372 21364 25384
rect 21416 25372 21422 25424
rect 27522 25372 27528 25424
rect 27580 25372 27586 25424
rect 28629 25415 28687 25421
rect 28629 25381 28641 25415
rect 28675 25412 28687 25415
rect 28675 25384 31432 25412
rect 28675 25381 28687 25384
rect 28629 25375 28687 25381
rect 20257 25347 20315 25353
rect 20257 25313 20269 25347
rect 20303 25313 20315 25347
rect 20257 25307 20315 25313
rect 20993 25347 21051 25353
rect 20993 25313 21005 25347
rect 21039 25344 21051 25347
rect 21634 25344 21640 25356
rect 21039 25316 21640 25344
rect 21039 25313 21051 25316
rect 20993 25307 21051 25313
rect 21634 25304 21640 25316
rect 21692 25304 21698 25356
rect 22738 25304 22744 25356
rect 22796 25344 22802 25356
rect 26145 25347 26203 25353
rect 22796 25316 22968 25344
rect 22796 25304 22802 25316
rect 18598 25236 18604 25288
rect 18656 25236 18662 25288
rect 19886 25236 19892 25288
rect 19944 25236 19950 25288
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25276 20407 25279
rect 20530 25276 20536 25288
rect 20395 25248 20536 25276
rect 20395 25245 20407 25248
rect 20349 25239 20407 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 20806 25276 20812 25288
rect 20640 25248 20812 25276
rect 20640 25208 20668 25248
rect 20806 25236 20812 25248
rect 20864 25236 20870 25288
rect 20898 25236 20904 25288
rect 20956 25236 20962 25288
rect 21085 25279 21143 25285
rect 21085 25245 21097 25279
rect 21131 25245 21143 25279
rect 21085 25239 21143 25245
rect 21177 25279 21235 25285
rect 21177 25245 21189 25279
rect 21223 25245 21235 25279
rect 21177 25239 21235 25245
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25276 21327 25279
rect 21358 25276 21364 25285
rect 21315 25248 21364 25276
rect 21315 25245 21327 25248
rect 21269 25239 21327 25245
rect 18524 25180 20668 25208
rect 20714 25168 20720 25220
rect 20772 25208 20778 25220
rect 21100 25208 21128 25239
rect 20772 25180 21128 25208
rect 20772 25168 20778 25180
rect 21192 25152 21220 25239
rect 21358 25233 21364 25248
rect 21416 25233 21422 25285
rect 22002 25236 22008 25288
rect 22060 25236 22066 25288
rect 22189 25279 22247 25285
rect 22189 25245 22201 25279
rect 22235 25276 22247 25279
rect 22278 25276 22284 25288
rect 22235 25248 22284 25276
rect 22235 25245 22247 25248
rect 22189 25239 22247 25245
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 22646 25236 22652 25288
rect 22704 25236 22710 25288
rect 22830 25236 22836 25288
rect 22888 25236 22894 25288
rect 22940 25285 22968 25316
rect 26145 25313 26157 25347
rect 26191 25344 26203 25347
rect 27540 25344 27568 25372
rect 26191 25316 27568 25344
rect 26191 25313 26203 25316
rect 26145 25307 26203 25313
rect 27890 25304 27896 25356
rect 27948 25344 27954 25356
rect 30282 25344 30288 25356
rect 27948 25316 30288 25344
rect 27948 25304 27954 25316
rect 22925 25279 22983 25285
rect 22925 25245 22937 25279
rect 22971 25245 22983 25279
rect 22925 25239 22983 25245
rect 23017 25279 23075 25285
rect 23017 25245 23029 25279
rect 23063 25276 23075 25279
rect 24302 25276 24308 25288
rect 23063 25248 24308 25276
rect 23063 25245 23075 25248
rect 23017 25239 23075 25245
rect 24302 25236 24308 25248
rect 24360 25236 24366 25288
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25245 25559 25279
rect 25501 25239 25559 25245
rect 21545 25211 21603 25217
rect 21545 25177 21557 25211
rect 21591 25208 21603 25211
rect 22097 25211 22155 25217
rect 22097 25208 22109 25211
rect 21591 25180 22109 25208
rect 21591 25177 21603 25180
rect 21545 25171 21603 25177
rect 22097 25177 22109 25180
rect 22143 25177 22155 25211
rect 22097 25171 22155 25177
rect 25133 25211 25191 25217
rect 25133 25177 25145 25211
rect 25179 25177 25191 25211
rect 25516 25208 25544 25239
rect 27982 25236 27988 25288
rect 28040 25236 28046 25288
rect 28166 25236 28172 25288
rect 28224 25236 28230 25288
rect 28368 25285 28396 25316
rect 30282 25304 30288 25316
rect 30340 25344 30346 25356
rect 30469 25347 30527 25353
rect 30469 25344 30481 25347
rect 30340 25316 30481 25344
rect 30340 25304 30346 25316
rect 30469 25313 30481 25316
rect 30515 25313 30527 25347
rect 30469 25307 30527 25313
rect 28261 25279 28319 25285
rect 28261 25245 28273 25279
rect 28307 25245 28319 25279
rect 28261 25239 28319 25245
rect 28353 25279 28411 25285
rect 28353 25245 28365 25279
rect 28399 25245 28411 25279
rect 28353 25239 28411 25245
rect 26326 25208 26332 25220
rect 25516 25180 26332 25208
rect 25133 25171 25191 25177
rect 15746 25140 15752 25152
rect 15120 25112 15752 25140
rect 15746 25100 15752 25112
rect 15804 25100 15810 25152
rect 18601 25143 18659 25149
rect 18601 25109 18613 25143
rect 18647 25140 18659 25143
rect 18782 25140 18788 25152
rect 18647 25112 18788 25140
rect 18647 25109 18659 25112
rect 18601 25103 18659 25109
rect 18782 25100 18788 25112
rect 18840 25100 18846 25152
rect 18874 25100 18880 25152
rect 18932 25140 18938 25152
rect 21174 25140 21180 25152
rect 18932 25112 21180 25140
rect 18932 25100 18938 25112
rect 21174 25100 21180 25112
rect 21232 25100 21238 25152
rect 21266 25100 21272 25152
rect 21324 25140 21330 25152
rect 21634 25149 21640 25152
rect 21453 25143 21511 25149
rect 21453 25140 21465 25143
rect 21324 25112 21465 25140
rect 21324 25100 21330 25112
rect 21453 25109 21465 25112
rect 21499 25109 21511 25143
rect 21631 25140 21640 25149
rect 21595 25112 21640 25140
rect 21453 25103 21511 25109
rect 21631 25103 21640 25112
rect 21634 25100 21640 25103
rect 21692 25100 21698 25152
rect 24762 25100 24768 25152
rect 24820 25100 24826 25152
rect 24933 25143 24991 25149
rect 24933 25109 24945 25143
rect 24979 25140 24991 25143
rect 25038 25140 25044 25152
rect 24979 25112 25044 25140
rect 24979 25109 24991 25112
rect 24933 25103 24991 25109
rect 25038 25100 25044 25112
rect 25096 25100 25102 25152
rect 25148 25140 25176 25171
rect 26326 25168 26332 25180
rect 26384 25168 26390 25220
rect 26421 25211 26479 25217
rect 26421 25177 26433 25211
rect 26467 25177 26479 25211
rect 26421 25171 26479 25177
rect 25314 25140 25320 25152
rect 25148 25112 25320 25140
rect 25314 25100 25320 25112
rect 25372 25140 25378 25152
rect 25866 25140 25872 25152
rect 25372 25112 25872 25140
rect 25372 25100 25378 25112
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 26053 25143 26111 25149
rect 26053 25109 26065 25143
rect 26099 25140 26111 25143
rect 26436 25140 26464 25171
rect 26878 25168 26884 25220
rect 26936 25168 26942 25220
rect 28276 25208 28304 25239
rect 30926 25236 30932 25288
rect 30984 25236 30990 25288
rect 31202 25236 31208 25288
rect 31260 25236 31266 25288
rect 31404 25285 31432 25384
rect 31496 25353 31524 25452
rect 32306 25440 32312 25492
rect 32364 25480 32370 25492
rect 32493 25483 32551 25489
rect 32493 25480 32505 25483
rect 32364 25452 32505 25480
rect 32364 25440 32370 25452
rect 32493 25449 32505 25452
rect 32539 25449 32551 25483
rect 32493 25443 32551 25449
rect 33134 25440 33140 25492
rect 33192 25480 33198 25492
rect 33229 25483 33287 25489
rect 33229 25480 33241 25483
rect 33192 25452 33241 25480
rect 33192 25440 33198 25452
rect 33229 25449 33241 25452
rect 33275 25449 33287 25483
rect 33229 25443 33287 25449
rect 34330 25440 34336 25492
rect 34388 25480 34394 25492
rect 35069 25483 35127 25489
rect 35069 25480 35081 25483
rect 34388 25452 35081 25480
rect 34388 25440 34394 25452
rect 35069 25449 35081 25452
rect 35115 25449 35127 25483
rect 35069 25443 35127 25449
rect 36722 25440 36728 25492
rect 36780 25440 36786 25492
rect 37001 25483 37059 25489
rect 37001 25449 37013 25483
rect 37047 25449 37059 25483
rect 37001 25443 37059 25449
rect 31481 25347 31539 25353
rect 31481 25313 31493 25347
rect 31527 25313 31539 25347
rect 31481 25307 31539 25313
rect 31570 25304 31576 25356
rect 31628 25304 31634 25356
rect 32324 25344 32352 25440
rect 35986 25372 35992 25424
rect 36044 25412 36050 25424
rect 37016 25412 37044 25443
rect 37458 25440 37464 25492
rect 37516 25480 37522 25492
rect 37737 25483 37795 25489
rect 37737 25480 37749 25483
rect 37516 25452 37749 25480
rect 37516 25440 37522 25452
rect 37737 25449 37749 25452
rect 37783 25449 37795 25483
rect 37737 25443 37795 25449
rect 37826 25440 37832 25492
rect 37884 25440 37890 25492
rect 36044 25384 37044 25412
rect 36044 25372 36050 25384
rect 37090 25344 37096 25356
rect 31772 25316 32352 25344
rect 36556 25316 37096 25344
rect 31772 25285 31800 25316
rect 31389 25279 31447 25285
rect 31389 25245 31401 25279
rect 31435 25245 31447 25279
rect 31389 25239 31447 25245
rect 31757 25279 31815 25285
rect 31757 25245 31769 25279
rect 31803 25245 31815 25279
rect 31757 25239 31815 25245
rect 32214 25236 32220 25288
rect 32272 25236 32278 25288
rect 32309 25279 32367 25285
rect 32309 25245 32321 25279
rect 32355 25245 32367 25279
rect 32309 25239 32367 25245
rect 29086 25208 29092 25220
rect 28276 25180 29092 25208
rect 29086 25168 29092 25180
rect 29144 25208 29150 25220
rect 30607 25211 30665 25217
rect 30607 25208 30619 25211
rect 29144 25180 30619 25208
rect 29144 25168 29150 25180
rect 30607 25177 30619 25180
rect 30653 25177 30665 25211
rect 30607 25171 30665 25177
rect 30742 25168 30748 25220
rect 30800 25168 30806 25220
rect 30837 25211 30895 25217
rect 30837 25177 30849 25211
rect 30883 25208 30895 25211
rect 31110 25208 31116 25220
rect 30883 25180 31116 25208
rect 30883 25177 30895 25180
rect 30837 25171 30895 25177
rect 31110 25168 31116 25180
rect 31168 25208 31174 25220
rect 32033 25211 32091 25217
rect 32033 25208 32045 25211
rect 31168 25180 32045 25208
rect 31168 25168 31174 25180
rect 32033 25177 32045 25180
rect 32079 25177 32091 25211
rect 32033 25171 32091 25177
rect 32122 25168 32128 25220
rect 32180 25208 32186 25220
rect 32324 25208 32352 25239
rect 32674 25236 32680 25288
rect 32732 25236 32738 25288
rect 32769 25279 32827 25285
rect 32769 25245 32781 25279
rect 32815 25245 32827 25279
rect 32769 25239 32827 25245
rect 32180 25180 32352 25208
rect 32180 25168 32186 25180
rect 32582 25168 32588 25220
rect 32640 25208 32646 25220
rect 32784 25208 32812 25239
rect 33410 25236 33416 25288
rect 33468 25236 33474 25288
rect 33594 25236 33600 25288
rect 33652 25236 33658 25288
rect 36556 25285 36584 25316
rect 37090 25304 37096 25316
rect 37148 25304 37154 25356
rect 37277 25347 37335 25353
rect 37277 25313 37289 25347
rect 37323 25344 37335 25347
rect 37323 25316 37964 25344
rect 37323 25313 37335 25316
rect 37277 25307 37335 25313
rect 37936 25288 37964 25316
rect 36541 25279 36599 25285
rect 36541 25245 36553 25279
rect 36587 25245 36599 25279
rect 36541 25239 36599 25245
rect 36725 25279 36783 25285
rect 36725 25245 36737 25279
rect 36771 25276 36783 25279
rect 36771 25248 36860 25276
rect 36771 25245 36783 25248
rect 36725 25239 36783 25245
rect 32640 25180 32812 25208
rect 32640 25168 32646 25180
rect 34698 25168 34704 25220
rect 34756 25168 34762 25220
rect 34882 25168 34888 25220
rect 34940 25168 34946 25220
rect 26099 25112 26464 25140
rect 26099 25109 26111 25112
rect 26053 25103 26111 25109
rect 27430 25100 27436 25152
rect 27488 25140 27494 25152
rect 27893 25143 27951 25149
rect 27893 25140 27905 25143
rect 27488 25112 27905 25140
rect 27488 25100 27494 25112
rect 27893 25109 27905 25112
rect 27939 25109 27951 25143
rect 27893 25103 27951 25109
rect 29822 25100 29828 25152
rect 29880 25100 29886 25152
rect 31941 25143 31999 25149
rect 31941 25109 31953 25143
rect 31987 25140 31999 25143
rect 32950 25140 32956 25152
rect 31987 25112 32956 25140
rect 31987 25109 31999 25112
rect 31941 25103 31999 25109
rect 32950 25100 32956 25112
rect 33008 25100 33014 25152
rect 36832 25149 36860 25248
rect 36906 25236 36912 25288
rect 36964 25276 36970 25288
rect 37369 25279 37427 25285
rect 36964 25248 37228 25276
rect 36964 25236 36970 25248
rect 37200 25217 37228 25248
rect 37369 25245 37381 25279
rect 37415 25245 37427 25279
rect 37369 25239 37427 25245
rect 37553 25279 37611 25285
rect 37553 25245 37565 25279
rect 37599 25276 37611 25279
rect 37734 25276 37740 25288
rect 37599 25248 37740 25276
rect 37599 25245 37611 25248
rect 37553 25239 37611 25245
rect 37185 25211 37243 25217
rect 37185 25177 37197 25211
rect 37231 25177 37243 25211
rect 37185 25171 37243 25177
rect 37384 25208 37412 25239
rect 37734 25236 37740 25248
rect 37792 25236 37798 25288
rect 37829 25279 37887 25285
rect 37829 25245 37841 25279
rect 37875 25245 37887 25279
rect 37829 25239 37887 25245
rect 37844 25208 37872 25239
rect 37918 25236 37924 25288
rect 37976 25236 37982 25288
rect 37384 25180 37872 25208
rect 38105 25211 38163 25217
rect 36998 25149 37004 25152
rect 36817 25143 36875 25149
rect 36817 25109 36829 25143
rect 36863 25109 36875 25143
rect 36817 25103 36875 25109
rect 36985 25143 37004 25149
rect 36985 25109 36997 25143
rect 36985 25103 37004 25109
rect 36998 25100 37004 25103
rect 37056 25100 37062 25152
rect 37090 25100 37096 25152
rect 37148 25140 37154 25152
rect 37384 25140 37412 25180
rect 38105 25177 38117 25211
rect 38151 25177 38163 25211
rect 38105 25171 38163 25177
rect 37148 25112 37412 25140
rect 37148 25100 37154 25112
rect 37826 25100 37832 25152
rect 37884 25140 37890 25152
rect 38120 25140 38148 25171
rect 37884 25112 38148 25140
rect 37884 25100 37890 25112
rect 1104 25050 38824 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 38824 25050
rect 1104 24976 38824 24998
rect 6086 24896 6092 24948
rect 6144 24936 6150 24948
rect 6181 24939 6239 24945
rect 6181 24936 6193 24939
rect 6144 24908 6193 24936
rect 6144 24896 6150 24908
rect 6181 24905 6193 24908
rect 6227 24905 6239 24939
rect 8018 24936 8024 24948
rect 6181 24899 6239 24905
rect 6748 24908 8024 24936
rect 4706 24868 4712 24880
rect 4172 24840 4712 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24769 1731 24803
rect 1673 24763 1731 24769
rect 2133 24803 2191 24809
rect 2133 24769 2145 24803
rect 2179 24769 2191 24803
rect 2133 24763 2191 24769
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24800 2651 24803
rect 2866 24800 2872 24812
rect 2639 24772 2872 24800
rect 2639 24769 2651 24772
rect 2593 24763 2651 24769
rect 1302 24624 1308 24676
rect 1360 24664 1366 24676
rect 1489 24667 1547 24673
rect 1489 24664 1501 24667
rect 1360 24636 1501 24664
rect 1360 24624 1366 24636
rect 1489 24633 1501 24636
rect 1535 24633 1547 24667
rect 1688 24664 1716 24763
rect 1762 24692 1768 24744
rect 1820 24692 1826 24744
rect 2038 24692 2044 24744
rect 2096 24692 2102 24744
rect 2148 24732 2176 24763
rect 2866 24760 2872 24772
rect 2924 24760 2930 24812
rect 4172 24809 4200 24840
rect 4706 24828 4712 24840
rect 4764 24828 4770 24880
rect 6270 24868 6276 24880
rect 5934 24840 6276 24868
rect 6270 24828 6276 24840
rect 6328 24868 6334 24880
rect 6748 24868 6776 24908
rect 8018 24896 8024 24908
rect 8076 24896 8082 24948
rect 9582 24896 9588 24948
rect 9640 24896 9646 24948
rect 12986 24896 12992 24948
rect 13044 24936 13050 24948
rect 13725 24939 13783 24945
rect 13725 24936 13737 24939
rect 13044 24908 13737 24936
rect 13044 24896 13050 24908
rect 13725 24905 13737 24908
rect 13771 24905 13783 24939
rect 13725 24899 13783 24905
rect 15194 24896 15200 24948
rect 15252 24936 15258 24948
rect 15289 24939 15347 24945
rect 15289 24936 15301 24939
rect 15252 24908 15301 24936
rect 15252 24896 15258 24908
rect 15289 24905 15301 24908
rect 15335 24905 15347 24939
rect 15838 24936 15844 24948
rect 15289 24899 15347 24905
rect 15396 24908 15844 24936
rect 8110 24868 8116 24880
rect 6328 24840 6776 24868
rect 6932 24840 8116 24868
rect 6328 24828 6334 24840
rect 4157 24803 4215 24809
rect 4157 24769 4169 24803
rect 4203 24769 4215 24803
rect 4157 24763 4215 24769
rect 6362 24760 6368 24812
rect 6420 24800 6426 24812
rect 6932 24809 6960 24840
rect 8110 24828 8116 24840
rect 8168 24828 8174 24880
rect 9030 24828 9036 24880
rect 9088 24828 9094 24880
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 6420 24772 6561 24800
rect 6420 24760 6426 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24769 6975 24803
rect 7193 24803 7251 24809
rect 7193 24800 7205 24803
rect 6917 24763 6975 24769
rect 7116 24772 7205 24800
rect 2685 24735 2743 24741
rect 2685 24732 2697 24735
rect 2148 24704 2697 24732
rect 2685 24701 2697 24704
rect 2731 24701 2743 24735
rect 2685 24695 2743 24701
rect 3142 24692 3148 24744
rect 3200 24732 3206 24744
rect 3237 24735 3295 24741
rect 3237 24732 3249 24735
rect 3200 24704 3249 24732
rect 3200 24692 3206 24704
rect 3237 24701 3249 24704
rect 3283 24701 3295 24735
rect 3237 24695 3295 24701
rect 3878 24692 3884 24744
rect 3936 24732 3942 24744
rect 4433 24735 4491 24741
rect 4433 24732 4445 24735
rect 3936 24704 4445 24732
rect 3936 24692 3942 24704
rect 4433 24701 4445 24704
rect 4479 24701 4491 24735
rect 4433 24695 4491 24701
rect 4709 24735 4767 24741
rect 4709 24701 4721 24735
rect 4755 24732 4767 24735
rect 5718 24732 5724 24744
rect 4755 24704 5724 24732
rect 4755 24701 4767 24704
rect 4709 24695 4767 24701
rect 5718 24692 5724 24704
rect 5776 24692 5782 24744
rect 6457 24735 6515 24741
rect 6457 24701 6469 24735
rect 6503 24732 6515 24735
rect 7006 24732 7012 24744
rect 6503 24704 7012 24732
rect 6503 24701 6515 24704
rect 6457 24695 6515 24701
rect 7006 24692 7012 24704
rect 7064 24692 7070 24744
rect 7116 24673 7144 24772
rect 7193 24769 7205 24772
rect 7239 24769 7251 24803
rect 7193 24763 7251 24769
rect 7469 24803 7527 24809
rect 7469 24769 7481 24803
rect 7515 24800 7527 24803
rect 7650 24800 7656 24812
rect 7515 24772 7656 24800
rect 7515 24769 7527 24772
rect 7469 24763 7527 24769
rect 7650 24760 7656 24772
rect 7708 24760 7714 24812
rect 8202 24760 8208 24812
rect 8260 24760 8266 24812
rect 8478 24760 8484 24812
rect 8536 24760 8542 24812
rect 8754 24760 8760 24812
rect 8812 24760 8818 24812
rect 8849 24803 8907 24809
rect 8849 24769 8861 24803
rect 8895 24769 8907 24803
rect 8849 24763 8907 24769
rect 7282 24692 7288 24744
rect 7340 24692 7346 24744
rect 7834 24692 7840 24744
rect 7892 24732 7898 24744
rect 8864 24732 8892 24763
rect 9122 24760 9128 24812
rect 9180 24760 9186 24812
rect 9600 24809 9628 24896
rect 14553 24871 14611 24877
rect 10152 24840 10364 24868
rect 9585 24803 9643 24809
rect 9585 24769 9597 24803
rect 9631 24769 9643 24803
rect 9585 24763 9643 24769
rect 9674 24760 9680 24812
rect 9732 24800 9738 24812
rect 10152 24800 10180 24840
rect 9732 24772 10180 24800
rect 9732 24760 9738 24772
rect 10226 24760 10232 24812
rect 10284 24760 10290 24812
rect 10336 24800 10364 24840
rect 13004 24840 14412 24868
rect 10505 24803 10563 24809
rect 10505 24800 10517 24803
rect 10336 24772 10517 24800
rect 10505 24769 10517 24772
rect 10551 24769 10563 24803
rect 10505 24763 10563 24769
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 7892 24704 8892 24732
rect 9493 24735 9551 24741
rect 7892 24692 7898 24704
rect 9493 24701 9505 24735
rect 9539 24732 9551 24735
rect 10318 24732 10324 24744
rect 9539 24704 10324 24732
rect 9539 24701 9551 24704
rect 9493 24695 9551 24701
rect 10318 24692 10324 24704
rect 10376 24692 10382 24744
rect 10612 24732 10640 24763
rect 10778 24760 10784 24812
rect 10836 24760 10842 24812
rect 11057 24803 11115 24809
rect 11057 24769 11069 24803
rect 11103 24800 11115 24803
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 11103 24772 11529 24800
rect 11103 24769 11115 24772
rect 11057 24763 11115 24769
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 12066 24760 12072 24812
rect 12124 24760 12130 24812
rect 12710 24760 12716 24812
rect 12768 24800 12774 24812
rect 13004 24809 13032 24840
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12768 24772 13001 24800
rect 12768 24760 12774 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13078 24760 13084 24812
rect 13136 24800 13142 24812
rect 13173 24803 13231 24809
rect 13173 24800 13185 24803
rect 13136 24772 13185 24800
rect 13136 24760 13142 24772
rect 13173 24769 13185 24772
rect 13219 24769 13231 24803
rect 13173 24763 13231 24769
rect 13357 24803 13415 24809
rect 13357 24769 13369 24803
rect 13403 24800 13415 24803
rect 13446 24800 13452 24812
rect 13403 24772 13452 24800
rect 13403 24769 13415 24772
rect 13357 24763 13415 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 13906 24760 13912 24812
rect 13964 24760 13970 24812
rect 14384 24809 14412 24840
rect 14553 24837 14565 24871
rect 14599 24868 14611 24871
rect 14826 24868 14832 24880
rect 14599 24840 14832 24868
rect 14599 24837 14611 24840
rect 14553 24831 14611 24837
rect 14826 24828 14832 24840
rect 14884 24868 14890 24880
rect 15396 24868 15424 24908
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 16209 24939 16267 24945
rect 16209 24905 16221 24939
rect 16255 24936 16267 24939
rect 16298 24936 16304 24948
rect 16255 24908 16304 24936
rect 16255 24905 16267 24908
rect 16209 24899 16267 24905
rect 16298 24896 16304 24908
rect 16356 24896 16362 24948
rect 18138 24896 18144 24948
rect 18196 24936 18202 24948
rect 18509 24939 18567 24945
rect 18509 24936 18521 24939
rect 18196 24908 18521 24936
rect 18196 24896 18202 24908
rect 18509 24905 18521 24908
rect 18555 24936 18567 24939
rect 19058 24936 19064 24948
rect 18555 24908 19064 24936
rect 18555 24905 18567 24908
rect 18509 24899 18567 24905
rect 19058 24896 19064 24908
rect 19116 24896 19122 24948
rect 19153 24939 19211 24945
rect 19153 24905 19165 24939
rect 19199 24905 19211 24939
rect 19153 24899 19211 24905
rect 14884 24840 15424 24868
rect 15488 24840 16252 24868
rect 14884 24828 14890 24840
rect 14001 24803 14059 24809
rect 14001 24769 14013 24803
rect 14047 24769 14059 24803
rect 14001 24763 14059 24769
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24769 14243 24803
rect 14185 24763 14243 24769
rect 14277 24803 14335 24809
rect 14277 24769 14289 24803
rect 14323 24769 14335 24803
rect 14277 24763 14335 24769
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 10965 24735 11023 24741
rect 10965 24732 10977 24735
rect 10612 24704 10977 24732
rect 2409 24667 2467 24673
rect 2409 24664 2421 24667
rect 1688 24636 2421 24664
rect 1489 24627 1547 24633
rect 2409 24633 2421 24636
rect 2455 24633 2467 24667
rect 2409 24627 2467 24633
rect 7101 24667 7159 24673
rect 7101 24633 7113 24667
rect 7147 24633 7159 24667
rect 7101 24627 7159 24633
rect 9858 24624 9864 24676
rect 9916 24664 9922 24676
rect 10612 24664 10640 24704
rect 10965 24701 10977 24704
rect 11011 24701 11023 24735
rect 13464 24732 13492 24760
rect 14016 24732 14044 24763
rect 13464 24704 14044 24732
rect 10965 24695 11023 24701
rect 9916 24636 10640 24664
rect 14200 24664 14228 24763
rect 14292 24732 14320 24763
rect 15194 24760 15200 24812
rect 15252 24760 15258 24812
rect 15488 24809 15516 24840
rect 16224 24812 16252 24840
rect 18782 24828 18788 24880
rect 18840 24828 18846 24880
rect 19168 24868 19196 24899
rect 19978 24896 19984 24948
rect 20036 24936 20042 24948
rect 20254 24936 20260 24948
rect 20036 24908 20260 24936
rect 20036 24896 20042 24908
rect 20254 24896 20260 24908
rect 20312 24896 20318 24948
rect 21545 24939 21603 24945
rect 21545 24905 21557 24939
rect 21591 24936 21603 24939
rect 21818 24936 21824 24948
rect 21591 24908 21824 24936
rect 21591 24905 21603 24908
rect 21545 24899 21603 24905
rect 21818 24896 21824 24908
rect 21876 24896 21882 24948
rect 22186 24896 22192 24948
rect 22244 24936 22250 24948
rect 22833 24939 22891 24945
rect 22833 24936 22845 24939
rect 22244 24908 22845 24936
rect 22244 24896 22250 24908
rect 22833 24905 22845 24908
rect 22879 24905 22891 24939
rect 22833 24899 22891 24905
rect 30742 24896 30748 24948
rect 30800 24936 30806 24948
rect 30929 24939 30987 24945
rect 30929 24936 30941 24939
rect 30800 24908 30941 24936
rect 30800 24896 30806 24908
rect 30929 24905 30941 24908
rect 30975 24905 30987 24939
rect 30929 24899 30987 24905
rect 31202 24896 31208 24948
rect 31260 24936 31266 24948
rect 31297 24939 31355 24945
rect 31297 24936 31309 24939
rect 31260 24908 31309 24936
rect 31260 24896 31266 24908
rect 31297 24905 31309 24908
rect 31343 24905 31355 24939
rect 31297 24899 31355 24905
rect 32582 24896 32588 24948
rect 32640 24896 32646 24948
rect 32674 24896 32680 24948
rect 32732 24896 32738 24948
rect 33410 24896 33416 24948
rect 33468 24936 33474 24948
rect 33781 24939 33839 24945
rect 33781 24936 33793 24939
rect 33468 24908 33793 24936
rect 33468 24896 33474 24908
rect 33781 24905 33793 24908
rect 33827 24905 33839 24939
rect 34517 24939 34575 24945
rect 33781 24899 33839 24905
rect 34164 24908 34468 24936
rect 20438 24868 20444 24880
rect 19168 24840 20444 24868
rect 20438 24828 20444 24840
rect 20496 24868 20502 24880
rect 22002 24868 22008 24880
rect 20496 24840 22008 24868
rect 20496 24828 20502 24840
rect 15473 24803 15531 24809
rect 15473 24769 15485 24803
rect 15519 24769 15531 24803
rect 15473 24763 15531 24769
rect 15565 24803 15623 24809
rect 15565 24769 15577 24803
rect 15611 24800 15623 24803
rect 15654 24800 15660 24812
rect 15611 24772 15660 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 15746 24760 15752 24812
rect 15804 24760 15810 24812
rect 15838 24760 15844 24812
rect 15896 24760 15902 24812
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 16117 24763 16175 24769
rect 15105 24735 15163 24741
rect 15105 24732 15117 24735
rect 14292 24704 15117 24732
rect 15105 24701 15117 24704
rect 15151 24732 15163 24735
rect 15378 24732 15384 24744
rect 15151 24704 15384 24732
rect 15151 24701 15163 24704
rect 15105 24695 15163 24701
rect 15378 24692 15384 24704
rect 15436 24692 15442 24744
rect 15672 24732 15700 24760
rect 16132 24732 16160 24763
rect 16206 24760 16212 24812
rect 16264 24800 16270 24812
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 16264 24772 16313 24800
rect 16264 24760 16270 24772
rect 16301 24769 16313 24772
rect 16347 24769 16359 24803
rect 16301 24763 16359 24769
rect 17770 24760 17776 24812
rect 17828 24800 17834 24812
rect 18141 24803 18199 24809
rect 18141 24800 18153 24803
rect 17828 24772 18153 24800
rect 17828 24760 17834 24772
rect 18141 24769 18153 24772
rect 18187 24769 18199 24803
rect 18141 24763 18199 24769
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 18601 24803 18659 24809
rect 18601 24769 18613 24803
rect 18647 24800 18659 24803
rect 18690 24800 18696 24812
rect 18647 24772 18696 24800
rect 18647 24769 18659 24772
rect 18601 24763 18659 24769
rect 15672 24704 16160 24732
rect 18340 24732 18368 24763
rect 18690 24760 18696 24772
rect 18748 24760 18754 24812
rect 18877 24803 18935 24809
rect 18877 24769 18889 24803
rect 18923 24769 18935 24803
rect 18877 24763 18935 24769
rect 18414 24732 18420 24744
rect 18340 24704 18420 24732
rect 18414 24692 18420 24704
rect 18472 24732 18478 24744
rect 18892 24732 18920 24763
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19978 24800 19984 24812
rect 19024 24772 19984 24800
rect 19024 24760 19030 24772
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20530 24760 20536 24812
rect 20588 24800 20594 24812
rect 21376 24809 21404 24840
rect 22002 24828 22008 24840
rect 22060 24828 22066 24880
rect 24762 24828 24768 24880
rect 24820 24828 24826 24880
rect 25498 24828 25504 24880
rect 25556 24828 25562 24880
rect 30668 24840 31248 24868
rect 21177 24803 21235 24809
rect 21177 24800 21189 24803
rect 20588 24772 21189 24800
rect 20588 24760 20594 24772
rect 21177 24769 21189 24772
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 21361 24803 21419 24809
rect 21361 24769 21373 24803
rect 21407 24769 21419 24803
rect 21361 24763 21419 24769
rect 21818 24760 21824 24812
rect 21876 24760 21882 24812
rect 22094 24760 22100 24812
rect 22152 24760 22158 24812
rect 22373 24803 22431 24809
rect 22373 24769 22385 24803
rect 22419 24769 22431 24803
rect 22373 24763 22431 24769
rect 18472 24704 18920 24732
rect 18472 24692 18478 24704
rect 19334 24692 19340 24744
rect 19392 24732 19398 24744
rect 20898 24732 20904 24744
rect 19392 24704 20904 24732
rect 19392 24692 19398 24704
rect 20898 24692 20904 24704
rect 20956 24732 20962 24744
rect 20956 24704 21772 24732
rect 20956 24692 20962 24704
rect 15746 24664 15752 24676
rect 14200 24636 15752 24664
rect 9916 24624 9922 24636
rect 15746 24624 15752 24636
rect 15804 24624 15810 24676
rect 2038 24556 2044 24608
rect 2096 24596 2102 24608
rect 2958 24596 2964 24608
rect 2096 24568 2964 24596
rect 2096 24556 2102 24568
rect 2958 24556 2964 24568
rect 3016 24556 3022 24608
rect 3418 24556 3424 24608
rect 3476 24596 3482 24608
rect 3513 24599 3571 24605
rect 3513 24596 3525 24599
rect 3476 24568 3525 24596
rect 3476 24556 3482 24568
rect 3513 24565 3525 24568
rect 3559 24565 3571 24599
rect 3513 24559 3571 24565
rect 6086 24556 6092 24608
rect 6144 24596 6150 24608
rect 6546 24596 6552 24608
rect 6144 24568 6552 24596
rect 6144 24556 6150 24568
rect 6546 24556 6552 24568
rect 6604 24596 6610 24608
rect 6825 24599 6883 24605
rect 6825 24596 6837 24599
rect 6604 24568 6837 24596
rect 6604 24556 6610 24568
rect 6825 24565 6837 24568
rect 6871 24565 6883 24599
rect 6825 24559 6883 24565
rect 6914 24556 6920 24608
rect 6972 24596 6978 24608
rect 7193 24599 7251 24605
rect 7193 24596 7205 24599
rect 6972 24568 7205 24596
rect 6972 24556 6978 24568
rect 7193 24565 7205 24568
rect 7239 24596 7251 24599
rect 7466 24596 7472 24608
rect 7239 24568 7472 24596
rect 7239 24565 7251 24568
rect 7193 24559 7251 24565
rect 7466 24556 7472 24568
rect 7524 24556 7530 24608
rect 7653 24599 7711 24605
rect 7653 24565 7665 24599
rect 7699 24596 7711 24599
rect 8110 24596 8116 24608
rect 7699 24568 8116 24596
rect 7699 24565 7711 24568
rect 7653 24559 7711 24565
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 9214 24556 9220 24608
rect 9272 24556 9278 24608
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 9769 24599 9827 24605
rect 9769 24596 9781 24599
rect 9364 24568 9781 24596
rect 9364 24556 9370 24568
rect 9769 24565 9781 24568
rect 9815 24565 9827 24599
rect 9769 24559 9827 24565
rect 10502 24556 10508 24608
rect 10560 24596 10566 24608
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 10560 24568 10793 24596
rect 10560 24556 10566 24568
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 10781 24559 10839 24565
rect 14737 24599 14795 24605
rect 14737 24565 14749 24599
rect 14783 24596 14795 24599
rect 15562 24596 15568 24608
rect 14783 24568 15568 24596
rect 14783 24565 14795 24568
rect 14737 24559 14795 24565
rect 15562 24556 15568 24568
rect 15620 24556 15626 24608
rect 21266 24556 21272 24608
rect 21324 24556 21330 24608
rect 21744 24596 21772 24704
rect 22002 24692 22008 24744
rect 22060 24732 22066 24744
rect 22388 24732 22416 24763
rect 22646 24760 22652 24812
rect 22704 24760 22710 24812
rect 23290 24809 23296 24812
rect 23284 24763 23296 24809
rect 23290 24760 23296 24763
rect 23348 24760 23354 24812
rect 24210 24760 24216 24812
rect 24268 24800 24274 24812
rect 24489 24803 24547 24809
rect 24489 24800 24501 24803
rect 24268 24772 24501 24800
rect 24268 24760 24274 24772
rect 24489 24769 24501 24772
rect 24535 24769 24547 24803
rect 24489 24763 24547 24769
rect 26418 24760 26424 24812
rect 26476 24800 26482 24812
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 26476 24772 27169 24800
rect 26476 24760 26482 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 27430 24760 27436 24812
rect 27488 24760 27494 24812
rect 28626 24760 28632 24812
rect 28684 24800 28690 24812
rect 30561 24803 30619 24809
rect 30561 24800 30573 24803
rect 28684 24772 30573 24800
rect 28684 24760 28690 24772
rect 30561 24769 30573 24772
rect 30607 24800 30619 24803
rect 30668 24800 30696 24840
rect 30607 24772 30696 24800
rect 30745 24803 30803 24809
rect 30607 24769 30619 24772
rect 30561 24763 30619 24769
rect 30745 24769 30757 24803
rect 30791 24769 30803 24803
rect 30745 24763 30803 24769
rect 22060 24704 22416 24732
rect 22060 24692 22066 24704
rect 22462 24692 22468 24744
rect 22520 24692 22526 24744
rect 22922 24692 22928 24744
rect 22980 24732 22986 24744
rect 23017 24735 23075 24741
rect 23017 24732 23029 24735
rect 22980 24704 23029 24732
rect 22980 24692 22986 24704
rect 23017 24701 23029 24704
rect 23063 24701 23075 24735
rect 23017 24695 23075 24701
rect 26970 24692 26976 24744
rect 27028 24692 27034 24744
rect 27249 24735 27307 24741
rect 27249 24732 27261 24735
rect 27080 24704 27261 24732
rect 26694 24624 26700 24676
rect 26752 24664 26758 24676
rect 27080 24664 27108 24704
rect 27249 24701 27261 24704
rect 27295 24701 27307 24735
rect 27249 24695 27307 24701
rect 27341 24735 27399 24741
rect 27341 24701 27353 24735
rect 27387 24701 27399 24735
rect 27341 24695 27399 24701
rect 26752 24636 27108 24664
rect 26752 24624 26758 24636
rect 27154 24624 27160 24676
rect 27212 24664 27218 24676
rect 27356 24664 27384 24695
rect 29086 24692 29092 24744
rect 29144 24692 29150 24744
rect 29546 24692 29552 24744
rect 29604 24692 29610 24744
rect 30760 24732 30788 24763
rect 30834 24760 30840 24812
rect 30892 24760 30898 24812
rect 31110 24760 31116 24812
rect 31168 24760 31174 24812
rect 31220 24800 31248 24840
rect 31570 24828 31576 24880
rect 31628 24828 31634 24880
rect 32600 24868 32628 24896
rect 32600 24840 33548 24868
rect 31389 24803 31447 24809
rect 31389 24800 31401 24803
rect 31220 24772 31401 24800
rect 31389 24769 31401 24772
rect 31435 24769 31447 24803
rect 31389 24763 31447 24769
rect 31757 24803 31815 24809
rect 31757 24769 31769 24803
rect 31803 24800 31815 24803
rect 32122 24800 32128 24812
rect 31803 24772 32128 24800
rect 31803 24769 31815 24772
rect 31757 24763 31815 24769
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 32217 24803 32275 24809
rect 32217 24769 32229 24803
rect 32263 24800 32275 24803
rect 32401 24803 32459 24809
rect 32263 24772 32352 24800
rect 32263 24769 32275 24772
rect 32217 24763 32275 24769
rect 31570 24732 31576 24744
rect 30760 24704 31576 24732
rect 31570 24692 31576 24704
rect 31628 24692 31634 24744
rect 32324 24676 32352 24772
rect 32401 24769 32413 24803
rect 32447 24800 32459 24803
rect 32674 24800 32680 24812
rect 32447 24772 32680 24800
rect 32447 24769 32459 24772
rect 32401 24763 32459 24769
rect 32674 24760 32680 24772
rect 32732 24760 32738 24812
rect 32769 24803 32827 24809
rect 32769 24769 32781 24803
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 32953 24803 33011 24809
rect 32953 24769 32965 24803
rect 32999 24769 33011 24803
rect 33060 24800 33088 24840
rect 33137 24803 33195 24809
rect 33137 24800 33149 24803
rect 33060 24772 33149 24800
rect 32953 24763 33011 24769
rect 33137 24769 33149 24772
rect 33183 24769 33195 24803
rect 33137 24763 33195 24769
rect 33229 24803 33287 24809
rect 33229 24769 33241 24803
rect 33275 24800 33287 24803
rect 33413 24803 33471 24809
rect 33275 24772 33364 24800
rect 33275 24769 33287 24772
rect 33229 24763 33287 24769
rect 27212 24636 27384 24664
rect 27212 24624 27218 24636
rect 28994 24624 29000 24676
rect 29052 24664 29058 24676
rect 29181 24667 29239 24673
rect 29181 24664 29193 24667
rect 29052 24636 29193 24664
rect 29052 24624 29058 24636
rect 29181 24633 29193 24636
rect 29227 24633 29239 24667
rect 29181 24627 29239 24633
rect 30653 24667 30711 24673
rect 30653 24633 30665 24667
rect 30699 24664 30711 24667
rect 32214 24664 32220 24676
rect 30699 24636 32220 24664
rect 30699 24633 30711 24636
rect 30653 24627 30711 24633
rect 32214 24624 32220 24636
rect 32272 24624 32278 24676
rect 32306 24624 32312 24676
rect 32364 24664 32370 24676
rect 32784 24664 32812 24763
rect 32364 24636 32812 24664
rect 32364 24624 32370 24636
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21744 24568 21833 24596
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 21821 24559 21879 24565
rect 22278 24556 22284 24608
rect 22336 24556 22342 24608
rect 22370 24556 22376 24608
rect 22428 24556 22434 24608
rect 24397 24599 24455 24605
rect 24397 24565 24409 24599
rect 24443 24596 24455 24599
rect 25222 24596 25228 24608
rect 24443 24568 25228 24596
rect 24443 24565 24455 24568
rect 24397 24559 24455 24565
rect 25222 24556 25228 24568
rect 25280 24556 25286 24608
rect 26234 24556 26240 24608
rect 26292 24596 26298 24608
rect 27172 24596 27200 24624
rect 26292 24568 27200 24596
rect 26292 24556 26298 24568
rect 32122 24556 32128 24608
rect 32180 24596 32186 24608
rect 32968 24596 32996 24763
rect 33336 24664 33364 24772
rect 33413 24769 33425 24803
rect 33459 24769 33471 24803
rect 33520 24800 33548 24840
rect 33594 24828 33600 24880
rect 33652 24868 33658 24880
rect 34164 24877 34192 24908
rect 34149 24871 34207 24877
rect 33652 24840 34100 24868
rect 33652 24828 33658 24840
rect 33689 24803 33747 24809
rect 33689 24800 33701 24803
rect 33520 24772 33701 24800
rect 33413 24763 33471 24769
rect 33689 24769 33701 24772
rect 33735 24769 33747 24803
rect 33689 24763 33747 24769
rect 33428 24732 33456 24763
rect 33778 24760 33784 24812
rect 33836 24800 33842 24812
rect 33873 24803 33931 24809
rect 33873 24800 33885 24803
rect 33836 24772 33885 24800
rect 33836 24760 33842 24772
rect 33873 24769 33885 24772
rect 33919 24769 33931 24803
rect 33873 24763 33931 24769
rect 33965 24803 34023 24809
rect 33965 24769 33977 24803
rect 34011 24769 34023 24803
rect 34072 24800 34100 24840
rect 34149 24837 34161 24871
rect 34195 24837 34207 24871
rect 34349 24871 34407 24877
rect 34349 24868 34361 24871
rect 34149 24831 34207 24837
rect 34348 24837 34361 24868
rect 34395 24837 34407 24871
rect 34440 24868 34468 24908
rect 34517 24905 34529 24939
rect 34563 24936 34575 24939
rect 34698 24936 34704 24948
rect 34563 24908 34704 24936
rect 34563 24905 34575 24908
rect 34517 24899 34575 24905
rect 34698 24896 34704 24908
rect 34756 24896 34762 24948
rect 35434 24896 35440 24948
rect 35492 24936 35498 24948
rect 35621 24939 35679 24945
rect 35621 24936 35633 24939
rect 35492 24908 35633 24936
rect 35492 24896 35498 24908
rect 35621 24905 35633 24908
rect 35667 24905 35679 24939
rect 35621 24899 35679 24905
rect 35986 24896 35992 24948
rect 36044 24896 36050 24948
rect 34440 24840 34836 24868
rect 34348 24831 34407 24837
rect 34348 24800 34376 24831
rect 34808 24812 34836 24840
rect 34609 24803 34667 24809
rect 34609 24800 34621 24803
rect 34072 24772 34621 24800
rect 33965 24763 34023 24769
rect 34609 24769 34621 24772
rect 34655 24769 34667 24803
rect 34609 24763 34667 24769
rect 34701 24803 34759 24809
rect 34701 24769 34713 24803
rect 34747 24769 34759 24803
rect 34701 24763 34759 24769
rect 33980 24732 34008 24763
rect 33428 24704 34008 24732
rect 33888 24676 33916 24704
rect 33686 24664 33692 24676
rect 33336 24636 33692 24664
rect 33686 24624 33692 24636
rect 33744 24624 33750 24676
rect 33870 24624 33876 24676
rect 33928 24624 33934 24676
rect 32180 24568 32996 24596
rect 32180 24556 32186 24568
rect 33778 24556 33784 24608
rect 33836 24596 33842 24608
rect 34333 24599 34391 24605
rect 34333 24596 34345 24599
rect 33836 24568 34345 24596
rect 33836 24556 33842 24568
rect 34333 24565 34345 24568
rect 34379 24596 34391 24599
rect 34716 24596 34744 24763
rect 34790 24760 34796 24812
rect 34848 24800 34854 24812
rect 34885 24803 34943 24809
rect 34885 24800 34897 24803
rect 34848 24772 34897 24800
rect 34848 24760 34854 24772
rect 34885 24769 34897 24772
rect 34931 24769 34943 24803
rect 34885 24763 34943 24769
rect 35253 24803 35311 24809
rect 35253 24769 35265 24803
rect 35299 24769 35311 24803
rect 35253 24763 35311 24769
rect 35268 24732 35296 24763
rect 35434 24760 35440 24812
rect 35492 24800 35498 24812
rect 35713 24803 35771 24809
rect 35713 24800 35725 24803
rect 35492 24772 35725 24800
rect 35492 24760 35498 24772
rect 35713 24769 35725 24772
rect 35759 24769 35771 24803
rect 36004 24800 36032 24896
rect 36725 24803 36783 24809
rect 36725 24800 36737 24803
rect 36004 24772 36737 24800
rect 35713 24763 35771 24769
rect 36725 24769 36737 24772
rect 36771 24769 36783 24803
rect 36725 24763 36783 24769
rect 36814 24760 36820 24812
rect 36872 24760 36878 24812
rect 36998 24760 37004 24812
rect 37056 24760 37062 24812
rect 34900 24704 35296 24732
rect 34900 24676 34928 24704
rect 34882 24624 34888 24676
rect 34940 24624 34946 24676
rect 35268 24664 35296 24704
rect 35345 24735 35403 24741
rect 35345 24701 35357 24735
rect 35391 24732 35403 24735
rect 35526 24732 35532 24744
rect 35391 24704 35532 24732
rect 35391 24701 35403 24704
rect 35345 24695 35403 24701
rect 35526 24692 35532 24704
rect 35584 24732 35590 24744
rect 35989 24735 36047 24741
rect 35989 24732 36001 24735
rect 35584 24704 36001 24732
rect 35584 24692 35590 24704
rect 35989 24701 36001 24704
rect 36035 24701 36047 24735
rect 35989 24695 36047 24701
rect 35805 24667 35863 24673
rect 35805 24664 35817 24667
rect 35268 24636 35817 24664
rect 35805 24633 35817 24636
rect 35851 24633 35863 24667
rect 35805 24627 35863 24633
rect 37001 24667 37059 24673
rect 37001 24633 37013 24667
rect 37047 24664 37059 24667
rect 37090 24664 37096 24676
rect 37047 24636 37096 24664
rect 37047 24633 37059 24636
rect 37001 24627 37059 24633
rect 37090 24624 37096 24636
rect 37148 24624 37154 24676
rect 34379 24568 34744 24596
rect 34379 24565 34391 24568
rect 34333 24559 34391 24565
rect 35434 24556 35440 24608
rect 35492 24556 35498 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 3234 24352 3240 24404
rect 3292 24352 3298 24404
rect 3970 24352 3976 24404
rect 4028 24392 4034 24404
rect 4525 24395 4583 24401
rect 4525 24392 4537 24395
rect 4028 24364 4537 24392
rect 4028 24352 4034 24364
rect 4525 24361 4537 24364
rect 4571 24361 4583 24395
rect 4525 24355 4583 24361
rect 5626 24352 5632 24404
rect 5684 24352 5690 24404
rect 7282 24352 7288 24404
rect 7340 24352 7346 24404
rect 7374 24352 7380 24404
rect 7432 24352 7438 24404
rect 7834 24352 7840 24404
rect 7892 24352 7898 24404
rect 8205 24395 8263 24401
rect 8205 24361 8217 24395
rect 8251 24392 8263 24395
rect 9306 24392 9312 24404
rect 8251 24364 9312 24392
rect 8251 24361 8263 24364
rect 8205 24355 8263 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 9490 24352 9496 24404
rect 9548 24392 9554 24404
rect 9585 24395 9643 24401
rect 9585 24392 9597 24395
rect 9548 24364 9597 24392
rect 9548 24352 9554 24364
rect 9585 24361 9597 24364
rect 9631 24361 9643 24395
rect 9585 24355 9643 24361
rect 11977 24395 12035 24401
rect 11977 24361 11989 24395
rect 12023 24392 12035 24395
rect 12066 24392 12072 24404
rect 12023 24364 12072 24392
rect 12023 24361 12035 24364
rect 11977 24355 12035 24361
rect 12066 24352 12072 24364
rect 12124 24352 12130 24404
rect 13265 24395 13323 24401
rect 13265 24392 13277 24395
rect 13096 24364 13277 24392
rect 4982 24284 4988 24336
rect 5040 24284 5046 24336
rect 7300 24324 7328 24352
rect 7208 24296 7328 24324
rect 3418 24256 3424 24268
rect 3252 24228 3424 24256
rect 2958 24148 2964 24200
rect 3016 24148 3022 24200
rect 3252 24197 3280 24228
rect 3418 24216 3424 24228
rect 3476 24216 3482 24268
rect 4706 24216 4712 24268
rect 4764 24216 4770 24268
rect 6546 24216 6552 24268
rect 6604 24216 6610 24268
rect 3237 24191 3295 24197
rect 3237 24157 3249 24191
rect 3283 24157 3295 24191
rect 3237 24151 3295 24157
rect 3326 24148 3332 24200
rect 3384 24148 3390 24200
rect 3513 24191 3571 24197
rect 3513 24157 3525 24191
rect 3559 24188 3571 24191
rect 3789 24191 3847 24197
rect 3789 24188 3801 24191
rect 3559 24160 3801 24188
rect 3559 24157 3571 24160
rect 3513 24151 3571 24157
rect 3789 24157 3801 24160
rect 3835 24157 3847 24191
rect 3789 24151 3847 24157
rect 4341 24191 4399 24197
rect 4341 24157 4353 24191
rect 4387 24188 4399 24191
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 4387 24160 4813 24188
rect 4387 24157 4399 24160
rect 4341 24151 4399 24157
rect 4801 24157 4813 24160
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 5905 24191 5963 24197
rect 5905 24157 5917 24191
rect 5951 24188 5963 24191
rect 6178 24188 6184 24200
rect 5951 24160 6184 24188
rect 5951 24157 5963 24160
rect 5905 24151 5963 24157
rect 3053 24123 3111 24129
rect 3053 24089 3065 24123
rect 3099 24120 3111 24123
rect 3142 24120 3148 24132
rect 3099 24092 3148 24120
rect 3099 24089 3111 24092
rect 3053 24083 3111 24089
rect 3142 24080 3148 24092
rect 3200 24120 3206 24132
rect 3200 24092 3556 24120
rect 3200 24080 3206 24092
rect 3418 24012 3424 24064
rect 3476 24012 3482 24064
rect 3528 24052 3556 24092
rect 3602 24080 3608 24132
rect 3660 24120 3666 24132
rect 4356 24120 4384 24151
rect 6178 24148 6184 24160
rect 6236 24148 6242 24200
rect 6564 24188 6592 24216
rect 6825 24191 6883 24197
rect 6825 24188 6837 24191
rect 6564 24160 6837 24188
rect 6825 24157 6837 24160
rect 6871 24157 6883 24191
rect 6825 24151 6883 24157
rect 6914 24148 6920 24200
rect 6972 24148 6978 24200
rect 7208 24188 7236 24296
rect 8754 24284 8760 24336
rect 8812 24324 8818 24336
rect 9401 24327 9459 24333
rect 9401 24324 9413 24327
rect 8812 24296 9413 24324
rect 8812 24284 8818 24296
rect 9401 24293 9413 24296
rect 9447 24293 9459 24327
rect 9401 24287 9459 24293
rect 7282 24216 7288 24268
rect 7340 24216 7346 24268
rect 7466 24216 7472 24268
rect 7524 24216 7530 24268
rect 8202 24216 8208 24268
rect 8260 24216 8266 24268
rect 9769 24259 9827 24265
rect 9769 24225 9781 24259
rect 9815 24256 9827 24259
rect 9858 24256 9864 24268
rect 9815 24228 9864 24256
rect 9815 24225 9827 24228
rect 9769 24219 9827 24225
rect 9858 24216 9864 24228
rect 9916 24216 9922 24268
rect 10226 24216 10232 24268
rect 10284 24216 10290 24268
rect 10502 24216 10508 24268
rect 10560 24216 10566 24268
rect 12897 24259 12955 24265
rect 12897 24225 12909 24259
rect 12943 24256 12955 24259
rect 13096 24256 13124 24364
rect 13265 24361 13277 24364
rect 13311 24392 13323 24395
rect 13906 24392 13912 24404
rect 13311 24364 13912 24392
rect 13311 24361 13323 24364
rect 13265 24355 13323 24361
rect 13906 24352 13912 24364
rect 13964 24352 13970 24404
rect 14093 24395 14151 24401
rect 14093 24361 14105 24395
rect 14139 24392 14151 24395
rect 14274 24392 14280 24404
rect 14139 24364 14280 24392
rect 14139 24361 14151 24364
rect 14093 24355 14151 24361
rect 14274 24352 14280 24364
rect 14332 24352 14338 24404
rect 14366 24352 14372 24404
rect 14424 24392 14430 24404
rect 14921 24395 14979 24401
rect 14921 24392 14933 24395
rect 14424 24364 14933 24392
rect 14424 24352 14430 24364
rect 14921 24361 14933 24364
rect 14967 24361 14979 24395
rect 15746 24392 15752 24404
rect 14921 24355 14979 24361
rect 15120 24364 15752 24392
rect 13173 24327 13231 24333
rect 13173 24293 13185 24327
rect 13219 24324 13231 24327
rect 13219 24296 14688 24324
rect 13219 24293 13231 24296
rect 13173 24287 13231 24293
rect 14660 24265 14688 24296
rect 15120 24268 15148 24364
rect 15746 24352 15752 24364
rect 15804 24352 15810 24404
rect 18049 24395 18107 24401
rect 18049 24361 18061 24395
rect 18095 24392 18107 24395
rect 19141 24392 19147 24404
rect 18095 24364 19147 24392
rect 18095 24361 18107 24364
rect 18049 24355 18107 24361
rect 19141 24352 19147 24364
rect 19199 24352 19205 24404
rect 19242 24352 19248 24404
rect 19300 24392 19306 24404
rect 19334 24392 19340 24404
rect 19300 24364 19340 24392
rect 19300 24352 19306 24364
rect 19334 24352 19340 24364
rect 19392 24352 19398 24404
rect 19429 24395 19487 24401
rect 19429 24361 19441 24395
rect 19475 24392 19487 24395
rect 19794 24392 19800 24404
rect 19475 24364 19800 24392
rect 19475 24361 19487 24364
rect 19429 24355 19487 24361
rect 19794 24352 19800 24364
rect 19852 24352 19858 24404
rect 19886 24352 19892 24404
rect 19944 24352 19950 24404
rect 21082 24352 21088 24404
rect 21140 24392 21146 24404
rect 21361 24395 21419 24401
rect 21361 24392 21373 24395
rect 21140 24364 21373 24392
rect 21140 24352 21146 24364
rect 21361 24361 21373 24364
rect 21407 24361 21419 24395
rect 21361 24355 21419 24361
rect 21821 24395 21879 24401
rect 21821 24361 21833 24395
rect 21867 24392 21879 24395
rect 21910 24392 21916 24404
rect 21867 24364 21916 24392
rect 21867 24361 21879 24364
rect 21821 24355 21879 24361
rect 21910 24352 21916 24364
rect 21968 24352 21974 24404
rect 23290 24352 23296 24404
rect 23348 24392 23354 24404
rect 23477 24395 23535 24401
rect 23477 24392 23489 24395
rect 23348 24364 23489 24392
rect 23348 24352 23354 24364
rect 23477 24361 23489 24364
rect 23523 24361 23535 24395
rect 23477 24355 23535 24361
rect 25038 24352 25044 24404
rect 25096 24392 25102 24404
rect 25133 24395 25191 24401
rect 25133 24392 25145 24395
rect 25096 24364 25145 24392
rect 25096 24352 25102 24364
rect 25133 24361 25145 24364
rect 25179 24361 25191 24395
rect 25133 24355 25191 24361
rect 25682 24352 25688 24404
rect 25740 24352 25746 24404
rect 26326 24352 26332 24404
rect 26384 24392 26390 24404
rect 26421 24395 26479 24401
rect 26421 24392 26433 24395
rect 26384 24364 26433 24392
rect 26384 24352 26390 24364
rect 26421 24361 26433 24364
rect 26467 24361 26479 24395
rect 26421 24355 26479 24361
rect 27709 24395 27767 24401
rect 27709 24361 27721 24395
rect 27755 24392 27767 24395
rect 27982 24392 27988 24404
rect 27755 24364 27988 24392
rect 27755 24361 27767 24364
rect 27709 24355 27767 24361
rect 27982 24352 27988 24364
rect 28040 24352 28046 24404
rect 28626 24352 28632 24404
rect 28684 24352 28690 24404
rect 29546 24392 29552 24404
rect 28736 24364 29552 24392
rect 15657 24327 15715 24333
rect 15657 24293 15669 24327
rect 15703 24293 15715 24327
rect 15657 24287 15715 24293
rect 12943 24228 13124 24256
rect 13725 24259 13783 24265
rect 12943 24225 12955 24228
rect 12897 24219 12955 24225
rect 13725 24225 13737 24259
rect 13771 24225 13783 24259
rect 13725 24219 13783 24225
rect 14645 24259 14703 24265
rect 14645 24225 14657 24259
rect 14691 24225 14703 24259
rect 14645 24219 14703 24225
rect 7377 24191 7435 24197
rect 7208 24182 7328 24188
rect 7377 24182 7389 24191
rect 7208 24160 7389 24182
rect 7300 24157 7389 24160
rect 7423 24157 7435 24191
rect 7300 24154 7435 24157
rect 7377 24151 7435 24154
rect 7650 24148 7656 24200
rect 7708 24148 7714 24200
rect 8110 24148 8116 24200
rect 8168 24148 8174 24200
rect 9214 24148 9220 24200
rect 9272 24188 9278 24200
rect 9585 24191 9643 24197
rect 9585 24188 9597 24191
rect 9272 24160 9597 24188
rect 9272 24148 9278 24160
rect 9585 24157 9597 24160
rect 9631 24157 9643 24191
rect 9585 24151 9643 24157
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24188 12863 24191
rect 12986 24188 12992 24200
rect 12851 24160 12992 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 12986 24148 12992 24160
rect 13044 24148 13050 24200
rect 13630 24148 13636 24200
rect 13688 24148 13694 24200
rect 13740 24188 13768 24219
rect 15102 24216 15108 24268
rect 15160 24216 15166 24268
rect 15562 24216 15568 24268
rect 15620 24216 15626 24268
rect 15672 24256 15700 24287
rect 16298 24284 16304 24336
rect 16356 24324 16362 24336
rect 16945 24327 17003 24333
rect 16356 24296 16804 24324
rect 16356 24284 16362 24296
rect 15672 24228 16712 24256
rect 14826 24188 14832 24200
rect 13740 24160 14832 24188
rect 14826 24148 14832 24160
rect 14884 24188 14890 24200
rect 15197 24191 15255 24197
rect 15197 24188 15209 24191
rect 14884 24160 15209 24188
rect 14884 24148 14890 24160
rect 15197 24157 15209 24160
rect 15243 24157 15255 24191
rect 15580 24188 15608 24216
rect 16132 24197 16160 24228
rect 15933 24191 15991 24197
rect 15933 24188 15945 24191
rect 15580 24160 15945 24188
rect 15197 24151 15255 24157
rect 15933 24157 15945 24160
rect 15979 24157 15991 24191
rect 15933 24151 15991 24157
rect 16117 24191 16175 24197
rect 16117 24157 16129 24191
rect 16163 24157 16175 24191
rect 16117 24151 16175 24157
rect 16209 24191 16267 24197
rect 16209 24157 16221 24191
rect 16255 24188 16267 24191
rect 16298 24188 16304 24200
rect 16255 24160 16304 24188
rect 16255 24157 16267 24160
rect 16209 24151 16267 24157
rect 16298 24148 16304 24160
rect 16356 24148 16362 24200
rect 16393 24191 16451 24197
rect 16393 24157 16405 24191
rect 16439 24188 16451 24191
rect 16482 24188 16488 24200
rect 16439 24160 16488 24188
rect 16439 24157 16451 24160
rect 16393 24151 16451 24157
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 16684 24197 16712 24228
rect 16776 24197 16804 24296
rect 16945 24293 16957 24327
rect 16991 24324 17003 24327
rect 17494 24324 17500 24336
rect 16991 24296 17500 24324
rect 16991 24293 17003 24296
rect 16945 24287 17003 24293
rect 17494 24284 17500 24296
rect 17552 24324 17558 24336
rect 18325 24327 18383 24333
rect 17552 24296 17908 24324
rect 17552 24284 17558 24296
rect 17880 24256 17908 24296
rect 18325 24293 18337 24327
rect 18371 24324 18383 24327
rect 19518 24324 19524 24336
rect 18371 24296 19524 24324
rect 18371 24293 18383 24296
rect 18325 24287 18383 24293
rect 19518 24284 19524 24296
rect 19576 24284 19582 24336
rect 19705 24327 19763 24333
rect 19705 24293 19717 24327
rect 19751 24324 19763 24327
rect 20070 24324 20076 24336
rect 19751 24296 20076 24324
rect 19751 24293 19763 24296
rect 19705 24287 19763 24293
rect 20070 24284 20076 24296
rect 20128 24324 20134 24336
rect 21634 24324 21640 24336
rect 20128 24296 21640 24324
rect 20128 24284 20134 24296
rect 21634 24284 21640 24296
rect 21692 24284 21698 24336
rect 22002 24284 22008 24336
rect 22060 24324 22066 24336
rect 22370 24324 22376 24336
rect 22060 24296 22376 24324
rect 22060 24284 22066 24296
rect 22370 24284 22376 24296
rect 22428 24284 22434 24336
rect 26234 24324 26240 24336
rect 25700 24296 26240 24324
rect 17880 24228 18276 24256
rect 17880 24197 17908 24228
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 16761 24191 16819 24197
rect 16761 24157 16773 24191
rect 16807 24157 16819 24191
rect 16761 24151 16819 24157
rect 17865 24191 17923 24197
rect 17865 24157 17877 24191
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 18138 24188 18144 24200
rect 18095 24160 18144 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18248 24197 18276 24228
rect 18414 24216 18420 24268
rect 18472 24216 18478 24268
rect 18506 24216 18512 24268
rect 18564 24216 18570 24268
rect 19797 24259 19855 24265
rect 19797 24225 19809 24259
rect 19843 24256 19855 24259
rect 20438 24256 20444 24268
rect 19843 24228 20444 24256
rect 19843 24225 19855 24228
rect 19797 24219 19855 24225
rect 20438 24216 20444 24228
rect 20496 24216 20502 24268
rect 21729 24259 21787 24265
rect 21729 24256 21741 24259
rect 21468 24228 21741 24256
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24157 18291 24191
rect 18432 24188 18460 24216
rect 18601 24191 18659 24197
rect 18601 24188 18613 24191
rect 18233 24151 18291 24157
rect 18340 24160 18613 24188
rect 3660 24092 4384 24120
rect 4525 24123 4583 24129
rect 3660 24080 3666 24092
rect 4525 24089 4537 24123
rect 4571 24089 4583 24123
rect 4525 24083 4583 24089
rect 5629 24123 5687 24129
rect 5629 24089 5641 24123
rect 5675 24120 5687 24123
rect 5997 24123 6055 24129
rect 5997 24120 6009 24123
rect 5675 24092 6009 24120
rect 5675 24089 5687 24092
rect 5629 24083 5687 24089
rect 5997 24089 6009 24092
rect 6043 24089 6055 24123
rect 5997 24083 6055 24089
rect 4540 24052 4568 24083
rect 7006 24080 7012 24132
rect 7064 24080 7070 24132
rect 7101 24123 7159 24129
rect 7101 24089 7113 24123
rect 7147 24120 7159 24123
rect 7466 24120 7472 24132
rect 7147 24092 7472 24120
rect 7147 24089 7159 24092
rect 7101 24083 7159 24089
rect 7466 24080 7472 24092
rect 7524 24120 7530 24132
rect 8294 24120 8300 24132
rect 7524 24092 8300 24120
rect 7524 24080 7530 24092
rect 8294 24080 8300 24092
rect 8352 24080 8358 24132
rect 9030 24080 9036 24132
rect 9088 24120 9094 24132
rect 10045 24123 10103 24129
rect 10045 24120 10057 24123
rect 9088 24092 10057 24120
rect 9088 24080 9094 24092
rect 10045 24089 10057 24092
rect 10091 24089 10103 24123
rect 11790 24120 11796 24132
rect 11730 24092 11796 24120
rect 10045 24083 10103 24089
rect 11790 24080 11796 24092
rect 11848 24080 11854 24132
rect 14553 24123 14611 24129
rect 14553 24089 14565 24123
rect 14599 24120 14611 24123
rect 15010 24120 15016 24132
rect 14599 24092 15016 24120
rect 14599 24089 14611 24092
rect 14553 24083 14611 24089
rect 15010 24080 15016 24092
rect 15068 24120 15074 24132
rect 15657 24123 15715 24129
rect 15657 24120 15669 24123
rect 15068 24092 15669 24120
rect 15068 24080 15074 24092
rect 15657 24089 15669 24092
rect 15703 24089 15715 24123
rect 16500 24120 16528 24148
rect 16945 24123 17003 24129
rect 16945 24120 16957 24123
rect 16500 24092 16957 24120
rect 15657 24083 15715 24089
rect 16945 24089 16957 24092
rect 16991 24089 17003 24123
rect 16945 24083 17003 24089
rect 17770 24080 17776 24132
rect 17828 24120 17834 24132
rect 18340 24120 18368 24160
rect 18601 24157 18613 24160
rect 18647 24157 18659 24191
rect 18779 24191 18837 24197
rect 18779 24188 18791 24191
rect 18601 24151 18659 24157
rect 18708 24160 18791 24188
rect 17828 24092 18368 24120
rect 17828 24080 17834 24092
rect 18414 24080 18420 24132
rect 18472 24120 18478 24132
rect 18509 24123 18567 24129
rect 18509 24120 18521 24123
rect 18472 24092 18521 24120
rect 18472 24080 18478 24092
rect 18509 24089 18521 24092
rect 18555 24089 18567 24123
rect 18708 24120 18736 24160
rect 18779 24157 18791 24160
rect 18825 24157 18837 24191
rect 18779 24151 18837 24157
rect 18874 24148 18880 24200
rect 18932 24190 18938 24200
rect 18932 24162 18975 24190
rect 18932 24148 18938 24162
rect 19058 24148 19064 24200
rect 19116 24148 19122 24200
rect 19150 24148 19156 24200
rect 19208 24190 19214 24200
rect 19981 24191 20039 24197
rect 19208 24188 19334 24190
rect 19981 24188 19993 24191
rect 19208 24162 19993 24188
rect 19208 24148 19214 24162
rect 19306 24160 19993 24162
rect 19981 24157 19993 24160
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20162 24148 20168 24200
rect 20220 24148 20226 24200
rect 20806 24148 20812 24200
rect 20864 24188 20870 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 20864 24160 21373 24188
rect 20864 24148 20870 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 18509 24083 18567 24089
rect 18616 24092 18736 24120
rect 18616 24064 18644 24092
rect 19242 24080 19248 24132
rect 19300 24120 19306 24132
rect 20070 24120 20076 24132
rect 19300 24092 20076 24120
rect 19300 24080 19306 24092
rect 20070 24080 20076 24092
rect 20128 24080 20134 24132
rect 21468 24120 21496 24228
rect 21729 24225 21741 24228
rect 21775 24225 21787 24259
rect 21729 24219 21787 24225
rect 21910 24216 21916 24268
rect 21968 24256 21974 24268
rect 25041 24259 25099 24265
rect 21968 24228 23152 24256
rect 21968 24216 21974 24228
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24157 21603 24191
rect 21545 24151 21603 24157
rect 21637 24191 21695 24197
rect 21637 24157 21649 24191
rect 21683 24188 21695 24191
rect 21818 24188 21824 24200
rect 21683 24160 21824 24188
rect 21683 24157 21695 24160
rect 21637 24151 21695 24157
rect 21376 24092 21496 24120
rect 21560 24120 21588 24151
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22278 24148 22284 24200
rect 22336 24188 22342 24200
rect 23124 24197 23152 24228
rect 25041 24225 25053 24259
rect 25087 24256 25099 24259
rect 25222 24256 25228 24268
rect 25087 24228 25228 24256
rect 25087 24225 25099 24228
rect 25041 24219 25099 24225
rect 25222 24216 25228 24228
rect 25280 24216 25286 24268
rect 25700 24256 25728 24296
rect 26234 24284 26240 24296
rect 26292 24284 26298 24336
rect 27157 24327 27215 24333
rect 27157 24293 27169 24327
rect 27203 24324 27215 24327
rect 28258 24324 28264 24336
rect 27203 24296 28264 24324
rect 27203 24293 27215 24296
rect 27157 24287 27215 24293
rect 28258 24284 28264 24296
rect 28316 24284 28322 24336
rect 28736 24324 28764 24364
rect 29546 24352 29552 24364
rect 29604 24352 29610 24404
rect 31570 24352 31576 24404
rect 31628 24392 31634 24404
rect 31849 24395 31907 24401
rect 31849 24392 31861 24395
rect 31628 24364 31861 24392
rect 31628 24352 31634 24364
rect 31849 24361 31861 24364
rect 31895 24361 31907 24395
rect 31849 24355 31907 24361
rect 32674 24352 32680 24404
rect 32732 24352 32738 24404
rect 33870 24352 33876 24404
rect 33928 24352 33934 24404
rect 35526 24352 35532 24404
rect 35584 24352 35590 24404
rect 36998 24352 37004 24404
rect 37056 24392 37062 24404
rect 37645 24395 37703 24401
rect 37645 24392 37657 24395
rect 37056 24364 37657 24392
rect 37056 24352 37062 24364
rect 37645 24361 37657 24364
rect 37691 24361 37703 24395
rect 37645 24355 37703 24361
rect 30193 24327 30251 24333
rect 30193 24324 30205 24327
rect 28644 24296 28764 24324
rect 28920 24296 30205 24324
rect 25332 24228 25728 24256
rect 25332 24197 25360 24228
rect 22833 24191 22891 24197
rect 22833 24188 22845 24191
rect 22336 24160 22845 24188
rect 22336 24148 22342 24160
rect 22833 24157 22845 24160
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24157 23075 24191
rect 23017 24151 23075 24157
rect 23109 24191 23167 24197
rect 23109 24157 23121 24191
rect 23155 24157 23167 24191
rect 23109 24151 23167 24157
rect 23201 24191 23259 24197
rect 23201 24157 23213 24191
rect 23247 24188 23259 24191
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 23247 24160 24409 24188
rect 23247 24157 23259 24160
rect 23201 24151 23259 24157
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24397 24151 24455 24157
rect 25317 24191 25375 24197
rect 25317 24157 25329 24191
rect 25363 24157 25375 24191
rect 25317 24151 25375 24157
rect 22094 24120 22100 24132
rect 21560 24092 22100 24120
rect 21376 24064 21404 24092
rect 22094 24080 22100 24092
rect 22152 24080 22158 24132
rect 23032 24120 23060 24151
rect 25590 24148 25596 24200
rect 25648 24148 25654 24200
rect 25700 24197 25728 24228
rect 27065 24259 27123 24265
rect 27065 24225 27077 24259
rect 27111 24256 27123 24259
rect 27246 24256 27252 24268
rect 27111 24228 27252 24256
rect 27111 24225 27123 24228
rect 27065 24219 27123 24225
rect 27246 24216 27252 24228
rect 27304 24216 27310 24268
rect 25685 24191 25743 24197
rect 25685 24157 25697 24191
rect 25731 24157 25743 24191
rect 25685 24151 25743 24157
rect 25777 24191 25835 24197
rect 25777 24157 25789 24191
rect 25823 24188 25835 24191
rect 26694 24188 26700 24200
rect 25823 24160 26700 24188
rect 25823 24157 25835 24160
rect 25777 24151 25835 24157
rect 23658 24120 23664 24132
rect 22848 24092 23664 24120
rect 22848 24064 22876 24092
rect 23658 24080 23664 24092
rect 23716 24080 23722 24132
rect 24762 24080 24768 24132
rect 24820 24120 24826 24132
rect 25501 24123 25559 24129
rect 25501 24120 25513 24123
rect 24820 24092 25513 24120
rect 24820 24080 24826 24092
rect 25501 24089 25513 24092
rect 25547 24120 25559 24123
rect 25792 24120 25820 24151
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 26789 24191 26847 24197
rect 26789 24157 26801 24191
rect 26835 24188 26847 24191
rect 27430 24188 27436 24200
rect 26835 24160 27436 24188
rect 26835 24157 26847 24160
rect 26789 24151 26847 24157
rect 27430 24148 27436 24160
rect 27488 24188 27494 24200
rect 28644 24197 28672 24296
rect 28810 24216 28816 24268
rect 28868 24216 28874 24268
rect 28920 24197 28948 24296
rect 30193 24293 30205 24296
rect 30239 24293 30251 24327
rect 36170 24324 36176 24336
rect 30193 24287 30251 24293
rect 35912 24296 36176 24324
rect 29273 24259 29331 24265
rect 29273 24225 29285 24259
rect 29319 24256 29331 24259
rect 29454 24256 29460 24268
rect 29319 24228 29460 24256
rect 29319 24225 29331 24228
rect 29273 24219 29331 24225
rect 29454 24216 29460 24228
rect 29512 24256 29518 24268
rect 31389 24259 31447 24265
rect 29512 24228 29776 24256
rect 29512 24216 29518 24228
rect 29748 24197 29776 24228
rect 31389 24225 31401 24259
rect 31435 24256 31447 24259
rect 33686 24256 33692 24268
rect 31435 24228 31800 24256
rect 31435 24225 31447 24228
rect 31389 24219 31447 24225
rect 27528 24191 27586 24197
rect 27528 24188 27540 24191
rect 27488 24160 27540 24188
rect 27488 24148 27494 24160
rect 27528 24157 27540 24160
rect 27574 24157 27586 24191
rect 27528 24151 27586 24157
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 28629 24191 28687 24197
rect 28629 24157 28641 24191
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 28905 24191 28963 24197
rect 28905 24157 28917 24191
rect 28951 24157 28963 24191
rect 28905 24151 28963 24157
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 25547 24092 25820 24120
rect 25961 24123 26019 24129
rect 25547 24089 25559 24092
rect 25501 24083 25559 24089
rect 25961 24089 25973 24123
rect 26007 24089 26019 24123
rect 25961 24083 26019 24089
rect 26973 24123 27031 24129
rect 26973 24089 26985 24123
rect 27019 24120 27031 24123
rect 27154 24120 27160 24132
rect 27019 24092 27160 24120
rect 27019 24089 27031 24092
rect 26973 24083 27031 24089
rect 3528 24024 4568 24052
rect 5813 24055 5871 24061
rect 5813 24021 5825 24055
rect 5859 24052 5871 24055
rect 6362 24052 6368 24064
rect 5859 24024 6368 24052
rect 5859 24021 5871 24024
rect 5813 24015 5871 24021
rect 6362 24012 6368 24024
rect 6420 24012 6426 24064
rect 8481 24055 8539 24061
rect 8481 24021 8493 24055
rect 8527 24052 8539 24055
rect 8754 24052 8760 24064
rect 8527 24024 8760 24052
rect 8527 24021 8539 24024
rect 8481 24015 8539 24021
rect 8754 24012 8760 24024
rect 8812 24012 8818 24064
rect 14461 24055 14519 24061
rect 14461 24021 14473 24055
rect 14507 24052 14519 24055
rect 14734 24052 14740 24064
rect 14507 24024 14740 24052
rect 14507 24021 14519 24024
rect 14461 24015 14519 24021
rect 14734 24012 14740 24024
rect 14792 24052 14798 24064
rect 15194 24052 15200 24064
rect 14792 24024 15200 24052
rect 14792 24012 14798 24024
rect 15194 24012 15200 24024
rect 15252 24052 15258 24064
rect 15841 24055 15899 24061
rect 15841 24052 15853 24055
rect 15252 24024 15853 24052
rect 15252 24012 15258 24024
rect 15841 24021 15853 24024
rect 15887 24052 15899 24055
rect 16390 24052 16396 24064
rect 15887 24024 16396 24052
rect 15887 24021 15899 24024
rect 15841 24015 15899 24021
rect 16390 24012 16396 24024
rect 16448 24012 16454 24064
rect 16574 24012 16580 24064
rect 16632 24012 16638 24064
rect 18598 24012 18604 24064
rect 18656 24012 18662 24064
rect 18693 24055 18751 24061
rect 18693 24021 18705 24055
rect 18739 24052 18751 24055
rect 18874 24052 18880 24064
rect 18739 24024 18880 24052
rect 18739 24021 18751 24024
rect 18693 24015 18751 24021
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 18969 24055 19027 24061
rect 18969 24021 18981 24055
rect 19015 24052 19027 24055
rect 21358 24052 21364 24064
rect 19015 24024 21364 24052
rect 19015 24021 19027 24024
rect 18969 24015 19027 24021
rect 21358 24012 21364 24024
rect 21416 24012 21422 24064
rect 21634 24012 21640 24064
rect 21692 24052 21698 24064
rect 22462 24052 22468 24064
rect 21692 24024 22468 24052
rect 21692 24012 21698 24024
rect 22462 24012 22468 24024
rect 22520 24012 22526 24064
rect 22830 24012 22836 24064
rect 22888 24012 22894 24064
rect 25590 24012 25596 24064
rect 25648 24052 25654 24064
rect 25976 24052 26004 24083
rect 27154 24080 27160 24092
rect 27212 24080 27218 24132
rect 26418 24052 26424 24064
rect 25648 24024 26424 24052
rect 25648 24012 25654 24024
rect 26418 24012 26424 24024
rect 26476 24052 26482 24064
rect 26605 24055 26663 24061
rect 26605 24052 26617 24055
rect 26476 24024 26617 24052
rect 26476 24012 26482 24024
rect 26605 24021 26617 24024
rect 26651 24021 26663 24055
rect 26605 24015 26663 24021
rect 26694 24012 26700 24064
rect 26752 24012 26758 24064
rect 27525 24055 27583 24061
rect 27525 24021 27537 24055
rect 27571 24052 27583 24055
rect 27706 24052 27712 24064
rect 27571 24024 27712 24052
rect 27571 24021 27583 24024
rect 27525 24015 27583 24021
rect 27706 24012 27712 24024
rect 27764 24012 27770 24064
rect 28368 24052 28396 24151
rect 28445 24123 28503 24129
rect 28445 24089 28457 24123
rect 28491 24120 28503 24123
rect 28920 24120 28948 24151
rect 30190 24148 30196 24200
rect 30248 24148 30254 24200
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 31772 24197 31800 24228
rect 32600 24228 33692 24256
rect 31021 24191 31079 24197
rect 31021 24188 31033 24191
rect 30432 24160 31033 24188
rect 30432 24148 30438 24160
rect 31021 24157 31033 24160
rect 31067 24188 31079 24191
rect 31481 24191 31539 24197
rect 31481 24188 31493 24191
rect 31067 24160 31493 24188
rect 31067 24157 31079 24160
rect 31021 24151 31079 24157
rect 31481 24157 31493 24160
rect 31527 24157 31539 24191
rect 31481 24151 31539 24157
rect 31665 24191 31723 24197
rect 31665 24157 31677 24191
rect 31711 24157 31723 24191
rect 31665 24151 31723 24157
rect 31757 24191 31815 24197
rect 31757 24157 31769 24191
rect 31803 24157 31815 24191
rect 31757 24151 31815 24157
rect 31941 24191 31999 24197
rect 31941 24157 31953 24191
rect 31987 24188 31999 24191
rect 32306 24188 32312 24200
rect 31987 24160 32312 24188
rect 31987 24157 31999 24160
rect 31941 24151 31999 24157
rect 28491 24092 28948 24120
rect 28491 24089 28503 24092
rect 28445 24083 28503 24089
rect 29362 24080 29368 24132
rect 29420 24120 29426 24132
rect 30101 24123 30159 24129
rect 30101 24120 30113 24123
rect 29420 24092 30113 24120
rect 29420 24080 29426 24092
rect 30101 24089 30113 24092
rect 30147 24089 30159 24123
rect 30101 24083 30159 24089
rect 31205 24123 31263 24129
rect 31205 24089 31217 24123
rect 31251 24120 31263 24123
rect 31570 24120 31576 24132
rect 31251 24092 31576 24120
rect 31251 24089 31263 24092
rect 31205 24083 31263 24089
rect 31570 24080 31576 24092
rect 31628 24120 31634 24132
rect 31680 24120 31708 24151
rect 31628 24092 31708 24120
rect 31628 24080 31634 24092
rect 28810 24052 28816 24064
rect 28368 24024 28816 24052
rect 28810 24012 28816 24024
rect 28868 24012 28874 24064
rect 28902 24012 28908 24064
rect 28960 24052 28966 24064
rect 29825 24055 29883 24061
rect 29825 24052 29837 24055
rect 28960 24024 29837 24052
rect 28960 24012 28966 24024
rect 29825 24021 29837 24024
rect 29871 24021 29883 24055
rect 29825 24015 29883 24021
rect 29917 24055 29975 24061
rect 29917 24021 29929 24055
rect 29963 24052 29975 24055
rect 30006 24052 30012 24064
rect 29963 24024 30012 24052
rect 29963 24021 29975 24024
rect 29917 24015 29975 24021
rect 30006 24012 30012 24024
rect 30064 24012 30070 24064
rect 31665 24055 31723 24061
rect 31665 24021 31677 24055
rect 31711 24052 31723 24055
rect 31956 24052 31984 24151
rect 32306 24148 32312 24160
rect 32364 24148 32370 24200
rect 32600 24197 32628 24228
rect 33686 24216 33692 24228
rect 33744 24216 33750 24268
rect 35912 24265 35940 24296
rect 36170 24284 36176 24296
rect 36228 24284 36234 24336
rect 36449 24327 36507 24333
rect 36449 24293 36461 24327
rect 36495 24324 36507 24327
rect 36814 24324 36820 24336
rect 36495 24296 36820 24324
rect 36495 24293 36507 24296
rect 36449 24287 36507 24293
rect 36814 24284 36820 24296
rect 36872 24284 36878 24336
rect 35897 24259 35955 24265
rect 35897 24225 35909 24259
rect 35943 24256 35955 24259
rect 35943 24228 36032 24256
rect 35943 24225 35955 24228
rect 35897 24219 35955 24225
rect 32585 24191 32643 24197
rect 32585 24157 32597 24191
rect 32631 24157 32643 24191
rect 32585 24151 32643 24157
rect 32769 24191 32827 24197
rect 32769 24157 32781 24191
rect 32815 24188 32827 24191
rect 32858 24188 32864 24200
rect 32815 24160 32864 24188
rect 32815 24157 32827 24160
rect 32769 24151 32827 24157
rect 32858 24148 32864 24160
rect 32916 24148 32922 24200
rect 33778 24148 33784 24200
rect 33836 24148 33842 24200
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 34514 24188 34520 24200
rect 34011 24160 34520 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 34514 24148 34520 24160
rect 34572 24148 34578 24200
rect 35805 24191 35863 24197
rect 35805 24157 35817 24191
rect 35851 24157 35863 24191
rect 36004 24188 36032 24228
rect 36070 24191 36128 24197
rect 36070 24188 36082 24191
rect 36004 24160 36082 24188
rect 35805 24151 35863 24157
rect 36070 24157 36082 24160
rect 36116 24157 36128 24191
rect 36070 24151 36128 24157
rect 36235 24191 36293 24197
rect 36235 24157 36247 24191
rect 36281 24188 36293 24191
rect 36354 24188 36360 24200
rect 36281 24160 36360 24188
rect 36281 24157 36308 24160
rect 36235 24151 36308 24157
rect 35820 24120 35848 24151
rect 36280 24120 36308 24151
rect 36354 24148 36360 24160
rect 36412 24148 36418 24200
rect 35820 24092 36308 24120
rect 36630 24080 36636 24132
rect 36688 24120 36694 24132
rect 37277 24123 37335 24129
rect 37277 24120 37289 24123
rect 36688 24092 37289 24120
rect 36688 24080 36694 24092
rect 37277 24089 37289 24092
rect 37323 24089 37335 24123
rect 37277 24083 37335 24089
rect 37461 24123 37519 24129
rect 37461 24089 37473 24123
rect 37507 24120 37519 24123
rect 37918 24120 37924 24132
rect 37507 24092 37924 24120
rect 37507 24089 37519 24092
rect 37461 24083 37519 24089
rect 37918 24080 37924 24092
rect 37976 24080 37982 24132
rect 31711 24024 31984 24052
rect 31711 24021 31723 24024
rect 31665 24015 31723 24021
rect 1104 23962 38824 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 38824 23962
rect 1104 23888 38824 23910
rect 2958 23808 2964 23860
rect 3016 23848 3022 23860
rect 3237 23851 3295 23857
rect 3237 23848 3249 23851
rect 3016 23820 3249 23848
rect 3016 23808 3022 23820
rect 3237 23817 3249 23820
rect 3283 23817 3295 23851
rect 3237 23811 3295 23817
rect 3957 23851 4015 23857
rect 3957 23817 3969 23851
rect 4003 23848 4015 23851
rect 5166 23848 5172 23860
rect 4003 23820 5172 23848
rect 4003 23817 4015 23820
rect 3957 23811 4015 23817
rect 5166 23808 5172 23820
rect 5224 23808 5230 23860
rect 8021 23851 8079 23857
rect 8021 23817 8033 23851
rect 8067 23848 8079 23851
rect 8202 23848 8208 23860
rect 8067 23820 8208 23848
rect 8067 23817 8079 23820
rect 8021 23811 8079 23817
rect 8202 23808 8208 23820
rect 8260 23808 8266 23860
rect 8294 23808 8300 23860
rect 8352 23848 8358 23860
rect 8481 23851 8539 23857
rect 8481 23848 8493 23851
rect 8352 23820 8493 23848
rect 8352 23808 8358 23820
rect 8481 23817 8493 23820
rect 8527 23817 8539 23851
rect 8481 23811 8539 23817
rect 8570 23808 8576 23860
rect 8628 23848 8634 23860
rect 9030 23848 9036 23860
rect 8628 23820 9036 23848
rect 8628 23808 8634 23820
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 9217 23851 9275 23857
rect 9217 23817 9229 23851
rect 9263 23848 9275 23851
rect 9582 23848 9588 23860
rect 9263 23820 9588 23848
rect 9263 23817 9275 23820
rect 9217 23811 9275 23817
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 9876 23820 11652 23848
rect 3050 23780 3056 23792
rect 2898 23752 3056 23780
rect 3050 23740 3056 23752
rect 3108 23740 3114 23792
rect 4157 23783 4215 23789
rect 4157 23749 4169 23783
rect 4203 23749 4215 23783
rect 4157 23743 4215 23749
rect 2958 23672 2964 23724
rect 3016 23712 3022 23724
rect 3326 23712 3332 23724
rect 3016 23684 3332 23712
rect 3016 23672 3022 23684
rect 3326 23672 3332 23684
rect 3384 23712 3390 23724
rect 3421 23715 3479 23721
rect 3421 23712 3433 23715
rect 3384 23684 3433 23712
rect 3384 23672 3390 23684
rect 3421 23681 3433 23684
rect 3467 23712 3479 23715
rect 3467 23684 3832 23712
rect 3467 23681 3479 23684
rect 3421 23675 3479 23681
rect 1394 23604 1400 23656
rect 1452 23604 1458 23656
rect 1670 23604 1676 23656
rect 1728 23604 1734 23656
rect 3145 23647 3203 23653
rect 3145 23613 3157 23647
rect 3191 23644 3203 23647
rect 3602 23644 3608 23656
rect 3191 23616 3608 23644
rect 3191 23613 3203 23616
rect 3145 23607 3203 23613
rect 3602 23604 3608 23616
rect 3660 23604 3666 23656
rect 3804 23585 3832 23684
rect 4172 23644 4200 23743
rect 8846 23740 8852 23792
rect 8904 23780 8910 23792
rect 9876 23789 9904 23820
rect 9861 23783 9919 23789
rect 9861 23780 9873 23783
rect 8904 23752 9873 23780
rect 8904 23740 8910 23752
rect 9861 23749 9873 23752
rect 9907 23749 9919 23783
rect 9861 23743 9919 23749
rect 10226 23740 10232 23792
rect 10284 23780 10290 23792
rect 10597 23783 10655 23789
rect 10597 23780 10609 23783
rect 10284 23752 10609 23780
rect 10284 23740 10290 23752
rect 10597 23749 10609 23752
rect 10643 23749 10655 23783
rect 10597 23743 10655 23749
rect 10778 23740 10784 23792
rect 10836 23780 10842 23792
rect 11241 23783 11299 23789
rect 11241 23780 11253 23783
rect 10836 23752 11253 23780
rect 10836 23740 10842 23752
rect 11241 23749 11253 23752
rect 11287 23749 11299 23783
rect 11241 23743 11299 23749
rect 8386 23721 8392 23724
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23712 7987 23715
rect 8364 23715 8392 23721
rect 7975 23684 8156 23712
rect 7975 23681 7987 23684
rect 7929 23675 7987 23681
rect 5350 23644 5356 23656
rect 4172 23616 5356 23644
rect 5350 23604 5356 23616
rect 5408 23644 5414 23656
rect 5994 23644 6000 23656
rect 5408 23616 6000 23644
rect 5408 23604 5414 23616
rect 5994 23604 6000 23616
rect 6052 23644 6058 23656
rect 7006 23644 7012 23656
rect 6052 23616 7012 23644
rect 6052 23604 6058 23616
rect 7006 23604 7012 23616
rect 7064 23604 7070 23656
rect 3789 23579 3847 23585
rect 3789 23545 3801 23579
rect 3835 23545 3847 23579
rect 3789 23539 3847 23545
rect 3970 23468 3976 23520
rect 4028 23468 4034 23520
rect 8128 23508 8156 23684
rect 8364 23681 8376 23715
rect 8364 23675 8392 23681
rect 8386 23672 8392 23675
rect 8444 23672 8450 23724
rect 8938 23672 8944 23724
rect 8996 23672 9002 23724
rect 9030 23672 9036 23724
rect 9088 23712 9094 23724
rect 9125 23715 9183 23721
rect 9125 23712 9137 23715
rect 9088 23684 9137 23712
rect 9088 23672 9094 23684
rect 9125 23681 9137 23684
rect 9171 23681 9183 23715
rect 9125 23675 9183 23681
rect 9214 23672 9220 23724
rect 9272 23672 9278 23724
rect 9582 23672 9588 23724
rect 9640 23672 9646 23724
rect 9766 23672 9772 23724
rect 9824 23672 9830 23724
rect 10873 23715 10931 23721
rect 10873 23681 10885 23715
rect 10919 23681 10931 23715
rect 10873 23675 10931 23681
rect 11057 23715 11115 23721
rect 11057 23681 11069 23715
rect 11103 23712 11115 23715
rect 11146 23712 11152 23724
rect 11103 23684 11152 23712
rect 11103 23681 11115 23684
rect 11057 23675 11115 23681
rect 8849 23647 8907 23653
rect 8849 23613 8861 23647
rect 8895 23644 8907 23647
rect 9232 23644 9260 23672
rect 8895 23616 9260 23644
rect 9677 23647 9735 23653
rect 8895 23613 8907 23616
rect 8849 23607 8907 23613
rect 9677 23613 9689 23647
rect 9723 23644 9735 23647
rect 10134 23644 10140 23656
rect 9723 23616 10140 23644
rect 9723 23613 9735 23616
rect 9677 23607 9735 23613
rect 10134 23604 10140 23616
rect 10192 23644 10198 23656
rect 10888 23644 10916 23675
rect 11146 23672 11152 23684
rect 11204 23672 11210 23724
rect 11624 23653 11652 23820
rect 13906 23808 13912 23860
rect 13964 23848 13970 23860
rect 14461 23851 14519 23857
rect 14461 23848 14473 23851
rect 13964 23820 14473 23848
rect 13964 23808 13970 23820
rect 14461 23817 14473 23820
rect 14507 23817 14519 23851
rect 14734 23848 14740 23860
rect 14461 23811 14519 23817
rect 14660 23820 14740 23848
rect 13446 23740 13452 23792
rect 13504 23740 13510 23792
rect 14660 23789 14688 23820
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 14826 23808 14832 23860
rect 14884 23808 14890 23860
rect 18506 23808 18512 23860
rect 18564 23808 18570 23860
rect 19242 23808 19248 23860
rect 19300 23808 19306 23860
rect 20070 23848 20076 23860
rect 19352 23820 20076 23848
rect 14645 23783 14703 23789
rect 14645 23749 14657 23783
rect 14691 23749 14703 23783
rect 14645 23743 14703 23749
rect 15013 23783 15071 23789
rect 15013 23749 15025 23783
rect 15059 23780 15071 23783
rect 15194 23780 15200 23792
rect 15059 23752 15200 23780
rect 15059 23749 15071 23752
rect 15013 23743 15071 23749
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 16761 23783 16819 23789
rect 15672 23752 16712 23780
rect 14366 23672 14372 23724
rect 14424 23672 14430 23724
rect 14737 23715 14795 23721
rect 14568 23710 14688 23712
rect 14737 23710 14749 23715
rect 14568 23684 14749 23710
rect 10192 23616 10916 23644
rect 11609 23647 11667 23653
rect 10192 23604 10198 23616
rect 11609 23613 11621 23647
rect 11655 23644 11667 23647
rect 12618 23644 12624 23656
rect 11655 23616 12624 23644
rect 11655 23613 11667 23616
rect 11609 23607 11667 23613
rect 12618 23604 12624 23616
rect 12676 23644 12682 23656
rect 13909 23647 13967 23653
rect 12676 23616 13852 23644
rect 12676 23604 12682 23616
rect 8205 23579 8263 23585
rect 8205 23545 8217 23579
rect 8251 23576 8263 23579
rect 9122 23576 9128 23588
rect 8251 23548 9128 23576
rect 8251 23545 8263 23548
rect 8205 23539 8263 23545
rect 9122 23536 9128 23548
rect 9180 23536 9186 23588
rect 12986 23536 12992 23588
rect 13044 23576 13050 23588
rect 13725 23579 13783 23585
rect 13725 23576 13737 23579
rect 13044 23548 13737 23576
rect 13044 23536 13050 23548
rect 13725 23545 13737 23548
rect 13771 23545 13783 23579
rect 13824 23576 13852 23616
rect 13909 23613 13921 23647
rect 13955 23644 13967 23647
rect 14568 23644 14596 23684
rect 14660 23682 14749 23684
rect 14737 23681 14749 23682
rect 14783 23712 14795 23715
rect 15102 23712 15108 23724
rect 14783 23684 15108 23712
rect 14783 23681 14795 23684
rect 14737 23675 14795 23681
rect 15102 23672 15108 23684
rect 15160 23672 15166 23724
rect 15672 23644 15700 23752
rect 16684 23721 16712 23752
rect 16761 23749 16773 23783
rect 16807 23780 16819 23783
rect 17589 23783 17647 23789
rect 17589 23780 17601 23783
rect 16807 23752 17601 23780
rect 16807 23749 16819 23752
rect 16761 23743 16819 23749
rect 16675 23715 16733 23721
rect 16675 23681 16687 23715
rect 16721 23681 16733 23715
rect 16675 23675 16733 23681
rect 16850 23672 16856 23724
rect 16908 23672 16914 23724
rect 17328 23721 17356 23752
rect 17589 23749 17601 23752
rect 17635 23780 17647 23783
rect 17635 23752 17908 23780
rect 17635 23749 17647 23752
rect 17589 23743 17647 23749
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23681 17371 23715
rect 17313 23675 17371 23681
rect 17494 23672 17500 23724
rect 17552 23672 17558 23724
rect 17773 23715 17831 23721
rect 17773 23681 17785 23715
rect 17819 23681 17831 23715
rect 17880 23712 17908 23752
rect 17954 23740 17960 23792
rect 18012 23740 18018 23792
rect 18141 23783 18199 23789
rect 18141 23749 18153 23783
rect 18187 23780 18199 23783
rect 18690 23780 18696 23792
rect 18187 23752 18696 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 18690 23740 18696 23752
rect 18748 23740 18754 23792
rect 19058 23740 19064 23792
rect 19116 23780 19122 23792
rect 19260 23780 19288 23808
rect 19352 23780 19380 23820
rect 20070 23808 20076 23820
rect 20128 23848 20134 23860
rect 20346 23848 20352 23860
rect 20128 23820 20352 23848
rect 20128 23808 20134 23820
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 20622 23808 20628 23860
rect 20680 23848 20686 23860
rect 22002 23848 22008 23860
rect 20680 23820 22008 23848
rect 20680 23808 20686 23820
rect 22002 23808 22008 23820
rect 22060 23808 22066 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23848 22247 23851
rect 22554 23848 22560 23860
rect 22235 23820 22560 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 22554 23808 22560 23820
rect 22612 23808 22618 23860
rect 28994 23808 29000 23860
rect 29052 23808 29058 23860
rect 30190 23808 30196 23860
rect 30248 23848 30254 23860
rect 30561 23851 30619 23857
rect 30561 23848 30573 23851
rect 30248 23820 30573 23848
rect 30248 23808 30254 23820
rect 30561 23817 30573 23820
rect 30607 23817 30619 23851
rect 30561 23811 30619 23817
rect 31570 23808 31576 23860
rect 31628 23848 31634 23860
rect 31665 23851 31723 23857
rect 31665 23848 31677 23851
rect 31628 23820 31677 23848
rect 31628 23808 31634 23820
rect 31665 23817 31677 23820
rect 31711 23817 31723 23851
rect 31665 23811 31723 23817
rect 32858 23808 32864 23860
rect 32916 23808 32922 23860
rect 33137 23851 33195 23857
rect 33137 23817 33149 23851
rect 33183 23848 33195 23851
rect 33686 23848 33692 23860
rect 33183 23820 33692 23848
rect 33183 23817 33195 23820
rect 33137 23811 33195 23817
rect 33686 23808 33692 23820
rect 33744 23808 33750 23860
rect 33778 23808 33784 23860
rect 33836 23848 33842 23860
rect 33965 23851 34023 23857
rect 33965 23848 33977 23851
rect 33836 23820 33977 23848
rect 33836 23808 33842 23820
rect 33965 23817 33977 23820
rect 34011 23817 34023 23851
rect 33965 23811 34023 23817
rect 34514 23808 34520 23860
rect 34572 23808 34578 23860
rect 34790 23808 34796 23860
rect 34848 23848 34854 23860
rect 35253 23851 35311 23857
rect 35253 23848 35265 23851
rect 34848 23820 35265 23848
rect 34848 23808 34854 23820
rect 35253 23817 35265 23820
rect 35299 23817 35311 23851
rect 35253 23811 35311 23817
rect 36354 23808 36360 23860
rect 36412 23808 36418 23860
rect 37918 23808 37924 23860
rect 37976 23808 37982 23860
rect 19116 23752 19187 23780
rect 19260 23752 19380 23780
rect 19429 23783 19487 23789
rect 19116 23740 19122 23752
rect 18049 23715 18107 23721
rect 18049 23712 18061 23715
rect 17880 23684 18061 23712
rect 17773 23675 17831 23681
rect 18049 23681 18061 23684
rect 18095 23681 18107 23715
rect 18227 23715 18285 23721
rect 18227 23712 18239 23715
rect 18049 23675 18107 23681
rect 18156 23684 18239 23712
rect 13955 23616 14596 23644
rect 14660 23616 15700 23644
rect 13955 23613 13967 23616
rect 13909 23607 13967 23613
rect 14182 23576 14188 23588
rect 13824 23548 14188 23576
rect 13725 23539 13783 23545
rect 14182 23536 14188 23548
rect 14240 23576 14246 23588
rect 14458 23576 14464 23588
rect 14240 23548 14464 23576
rect 14240 23536 14246 23548
rect 14458 23536 14464 23548
rect 14516 23536 14522 23588
rect 14660 23585 14688 23616
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 17788 23644 17816 23675
rect 18156 23656 18184 23684
rect 18227 23681 18239 23684
rect 18273 23681 18285 23715
rect 18227 23675 18285 23681
rect 18874 23672 18880 23724
rect 18932 23712 18938 23724
rect 19159 23712 19187 23752
rect 19429 23749 19441 23783
rect 19475 23780 19487 23783
rect 20162 23780 20168 23792
rect 19475 23752 20168 23780
rect 19475 23749 19487 23752
rect 19429 23743 19487 23749
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 19245 23715 19303 23721
rect 19245 23712 19257 23715
rect 18932 23702 19012 23712
rect 19055 23705 19113 23711
rect 19055 23702 19067 23705
rect 18932 23684 19067 23702
rect 18932 23672 18938 23684
rect 18984 23674 19067 23684
rect 18138 23644 18144 23656
rect 16632 23616 18144 23644
rect 16632 23604 16638 23616
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 18782 23604 18788 23656
rect 18840 23604 18846 23656
rect 14645 23579 14703 23585
rect 14645 23545 14657 23579
rect 14691 23545 14703 23579
rect 14645 23539 14703 23545
rect 15010 23536 15016 23588
rect 15068 23536 15074 23588
rect 18984 23576 19012 23674
rect 19055 23671 19067 23674
rect 19101 23671 19113 23705
rect 19159 23684 19257 23712
rect 19245 23681 19257 23684
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 19334 23672 19340 23724
rect 19392 23712 19398 23724
rect 19521 23715 19579 23721
rect 19521 23712 19533 23715
rect 19392 23684 19533 23712
rect 19392 23672 19398 23684
rect 19521 23681 19533 23684
rect 19567 23681 19579 23715
rect 19521 23675 19579 23681
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23681 19671 23715
rect 19613 23675 19671 23681
rect 19055 23665 19113 23671
rect 19628 23644 19656 23675
rect 19978 23672 19984 23724
rect 20036 23672 20042 23724
rect 20254 23672 20260 23724
rect 20312 23672 20318 23724
rect 20364 23721 20392 23808
rect 22830 23740 22836 23792
rect 22888 23780 22894 23792
rect 26973 23783 27031 23789
rect 26973 23780 26985 23783
rect 22888 23752 26985 23780
rect 22888 23740 22894 23752
rect 26973 23749 26985 23752
rect 27019 23780 27031 23783
rect 28261 23783 28319 23789
rect 28261 23780 28273 23783
rect 27019 23752 28273 23780
rect 27019 23749 27031 23752
rect 26973 23743 27031 23749
rect 28261 23749 28273 23752
rect 28307 23780 28319 23783
rect 28534 23780 28540 23792
rect 28307 23752 28540 23780
rect 28307 23749 28319 23752
rect 28261 23743 28319 23749
rect 28534 23740 28540 23752
rect 28592 23740 28598 23792
rect 30006 23780 30012 23792
rect 29288 23752 30012 23780
rect 29288 23724 29316 23752
rect 30006 23740 30012 23752
rect 30064 23740 30070 23792
rect 30374 23740 30380 23792
rect 30432 23740 30438 23792
rect 32677 23783 32735 23789
rect 32677 23749 32689 23783
rect 32723 23780 32735 23783
rect 33042 23780 33048 23792
rect 32723 23752 33048 23780
rect 32723 23749 32735 23752
rect 32677 23743 32735 23749
rect 33042 23740 33048 23752
rect 33100 23780 33106 23792
rect 34149 23783 34207 23789
rect 33100 23752 33180 23780
rect 33100 23740 33106 23752
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23681 20407 23715
rect 20349 23675 20407 23681
rect 21082 23672 21088 23724
rect 21140 23712 21146 23724
rect 21177 23715 21235 23721
rect 21177 23712 21189 23715
rect 21140 23684 21189 23712
rect 21140 23672 21146 23684
rect 21177 23681 21189 23684
rect 21223 23681 21235 23715
rect 21177 23675 21235 23681
rect 21358 23672 21364 23724
rect 21416 23672 21422 23724
rect 21818 23672 21824 23724
rect 21876 23672 21882 23724
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23712 22063 23715
rect 22462 23712 22468 23724
rect 22051 23684 22468 23712
rect 22051 23681 22063 23684
rect 22005 23675 22063 23681
rect 22462 23672 22468 23684
rect 22520 23672 22526 23724
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23712 24455 23715
rect 24762 23712 24768 23724
rect 24443 23684 24768 23712
rect 24443 23681 24455 23684
rect 24397 23675 24455 23681
rect 24762 23672 24768 23684
rect 24820 23712 24826 23724
rect 25041 23715 25099 23721
rect 25041 23712 25053 23715
rect 24820 23684 25053 23712
rect 24820 23672 24826 23684
rect 25041 23681 25053 23684
rect 25087 23681 25099 23715
rect 25041 23675 25099 23681
rect 25314 23672 25320 23724
rect 25372 23712 25378 23724
rect 25409 23715 25467 23721
rect 25409 23712 25421 23715
rect 25372 23684 25421 23712
rect 25372 23672 25378 23684
rect 25409 23681 25421 23684
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 25498 23672 25504 23724
rect 25556 23672 25562 23724
rect 26697 23715 26755 23721
rect 26697 23681 26709 23715
rect 26743 23681 26755 23715
rect 26697 23675 26755 23681
rect 19889 23647 19947 23653
rect 19889 23644 19901 23647
rect 19266 23616 19656 23644
rect 19720 23616 19901 23644
rect 19266 23576 19294 23616
rect 15120 23548 18828 23576
rect 18984 23548 19294 23576
rect 8478 23508 8484 23520
rect 8128 23480 8484 23508
rect 8478 23468 8484 23480
rect 8536 23508 8542 23520
rect 8938 23508 8944 23520
rect 8536 23480 8944 23508
rect 8536 23468 8542 23480
rect 8938 23468 8944 23480
rect 8996 23468 9002 23520
rect 11146 23468 11152 23520
rect 11204 23508 11210 23520
rect 15120 23508 15148 23548
rect 11204 23480 15148 23508
rect 11204 23468 11210 23480
rect 16114 23468 16120 23520
rect 16172 23508 16178 23520
rect 16850 23508 16856 23520
rect 16172 23480 16856 23508
rect 16172 23468 16178 23480
rect 16850 23468 16856 23480
rect 16908 23468 16914 23520
rect 17405 23511 17463 23517
rect 17405 23477 17417 23511
rect 17451 23508 17463 23511
rect 18046 23508 18052 23520
rect 17451 23480 18052 23508
rect 17451 23477 17463 23480
rect 17405 23471 17463 23477
rect 18046 23468 18052 23480
rect 18104 23508 18110 23520
rect 18690 23508 18696 23520
rect 18104 23480 18696 23508
rect 18104 23468 18110 23480
rect 18690 23468 18696 23480
rect 18748 23468 18754 23520
rect 18800 23508 18828 23548
rect 19334 23536 19340 23588
rect 19392 23576 19398 23588
rect 19720 23576 19748 23616
rect 19889 23613 19901 23616
rect 19935 23613 19947 23647
rect 20806 23644 20812 23656
rect 19889 23607 19947 23613
rect 20387 23616 20812 23644
rect 19392 23548 19748 23576
rect 19797 23579 19855 23585
rect 19392 23536 19398 23548
rect 19797 23545 19809 23579
rect 19843 23576 19855 23579
rect 20387 23576 20415 23616
rect 20806 23604 20812 23616
rect 20864 23604 20870 23656
rect 24121 23647 24179 23653
rect 24121 23613 24133 23647
rect 24167 23644 24179 23647
rect 25332 23644 25360 23672
rect 24167 23616 25360 23644
rect 24167 23613 24179 23616
rect 24121 23607 24179 23613
rect 26234 23604 26240 23656
rect 26292 23644 26298 23656
rect 26712 23644 26740 23675
rect 27154 23672 27160 23724
rect 27212 23712 27218 23724
rect 27985 23715 28043 23721
rect 27985 23712 27997 23715
rect 27212 23684 27997 23712
rect 27212 23672 27218 23684
rect 27985 23681 27997 23684
rect 28031 23681 28043 23715
rect 27985 23675 28043 23681
rect 28169 23715 28227 23721
rect 28169 23681 28181 23715
rect 28215 23681 28227 23715
rect 28169 23675 28227 23681
rect 27522 23644 27528 23656
rect 26292 23616 27528 23644
rect 26292 23604 26298 23616
rect 27522 23604 27528 23616
rect 27580 23644 27586 23656
rect 27709 23647 27767 23653
rect 27709 23644 27721 23647
rect 27580 23616 27721 23644
rect 27580 23604 27586 23616
rect 27709 23613 27721 23616
rect 27755 23613 27767 23647
rect 27709 23607 27767 23613
rect 19843 23548 20415 23576
rect 19843 23545 19855 23548
rect 19797 23539 19855 23545
rect 20438 23508 20444 23520
rect 18800 23480 20444 23508
rect 20438 23468 20444 23480
rect 20496 23468 20502 23520
rect 20533 23511 20591 23517
rect 20533 23477 20545 23511
rect 20579 23508 20591 23511
rect 20622 23508 20628 23520
rect 20579 23480 20628 23508
rect 20579 23477 20591 23480
rect 20533 23471 20591 23477
rect 20622 23468 20628 23480
rect 20680 23468 20686 23520
rect 20824 23508 20852 23604
rect 21177 23579 21235 23585
rect 21177 23545 21189 23579
rect 21223 23576 21235 23579
rect 22094 23576 22100 23588
rect 21223 23548 22100 23576
rect 21223 23545 21235 23548
rect 21177 23539 21235 23545
rect 22094 23536 22100 23548
rect 22152 23536 22158 23588
rect 24302 23536 24308 23588
rect 24360 23576 24366 23588
rect 25590 23576 25596 23588
rect 24360 23548 25596 23576
rect 24360 23536 24366 23548
rect 25590 23536 25596 23548
rect 25648 23536 25654 23588
rect 26878 23536 26884 23588
rect 26936 23576 26942 23588
rect 28184 23576 28212 23675
rect 28902 23672 28908 23724
rect 28960 23712 28966 23724
rect 29181 23715 29239 23721
rect 29181 23712 29193 23715
rect 28960 23684 29193 23712
rect 28960 23672 28966 23684
rect 29181 23681 29193 23684
rect 29227 23681 29239 23715
rect 29181 23675 29239 23681
rect 29270 23672 29276 23724
rect 29328 23672 29334 23724
rect 29362 23672 29368 23724
rect 29420 23672 29426 23724
rect 29454 23672 29460 23724
rect 29512 23672 29518 23724
rect 30190 23672 30196 23724
rect 30248 23712 30254 23724
rect 30469 23715 30527 23721
rect 30469 23712 30481 23715
rect 30248 23684 30481 23712
rect 30248 23672 30254 23684
rect 30469 23681 30481 23684
rect 30515 23681 30527 23715
rect 30469 23675 30527 23681
rect 30653 23715 30711 23721
rect 30653 23681 30665 23715
rect 30699 23681 30711 23715
rect 30653 23675 30711 23681
rect 30009 23647 30067 23653
rect 30009 23613 30021 23647
rect 30055 23644 30067 23647
rect 30098 23644 30104 23656
rect 30055 23616 30104 23644
rect 30055 23613 30067 23616
rect 30009 23607 30067 23613
rect 30098 23604 30104 23616
rect 30156 23644 30162 23656
rect 30668 23644 30696 23675
rect 31570 23672 31576 23724
rect 31628 23672 31634 23724
rect 31757 23715 31815 23721
rect 31757 23681 31769 23715
rect 31803 23712 31815 23715
rect 32122 23712 32128 23724
rect 31803 23684 32128 23712
rect 31803 23681 31815 23684
rect 31757 23675 31815 23681
rect 32122 23672 32128 23684
rect 32180 23712 32186 23724
rect 33152 23721 33180 23752
rect 34149 23749 34161 23783
rect 34195 23780 34207 23783
rect 34195 23752 34652 23780
rect 34195 23749 34207 23752
rect 34149 23743 34207 23749
rect 34624 23724 34652 23752
rect 36630 23740 36636 23792
rect 36688 23740 36694 23792
rect 37001 23783 37059 23789
rect 37001 23749 37013 23783
rect 37047 23780 37059 23783
rect 37047 23752 37504 23780
rect 37047 23749 37059 23752
rect 37001 23743 37059 23749
rect 37476 23724 37504 23752
rect 32493 23715 32551 23721
rect 32493 23712 32505 23715
rect 32180 23684 32505 23712
rect 32180 23672 32186 23684
rect 32493 23681 32505 23684
rect 32539 23712 32551 23715
rect 32953 23715 33011 23721
rect 32953 23712 32965 23715
rect 32539 23684 32965 23712
rect 32539 23681 32551 23684
rect 32493 23675 32551 23681
rect 32953 23681 32965 23684
rect 32999 23681 33011 23715
rect 32953 23675 33011 23681
rect 33137 23715 33195 23721
rect 33137 23681 33149 23715
rect 33183 23681 33195 23715
rect 33137 23675 33195 23681
rect 34330 23672 34336 23724
rect 34388 23712 34394 23724
rect 34425 23715 34483 23721
rect 34425 23712 34437 23715
rect 34388 23684 34437 23712
rect 34388 23672 34394 23684
rect 34425 23681 34437 23684
rect 34471 23681 34483 23715
rect 34425 23675 34483 23681
rect 34606 23672 34612 23724
rect 34664 23672 34670 23724
rect 34790 23672 34796 23724
rect 34848 23712 34854 23724
rect 34885 23715 34943 23721
rect 34885 23712 34897 23715
rect 34848 23684 34897 23712
rect 34848 23672 34854 23684
rect 34885 23681 34897 23684
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 35069 23715 35127 23721
rect 35069 23681 35081 23715
rect 35115 23712 35127 23715
rect 35434 23712 35440 23724
rect 35115 23684 35440 23712
rect 35115 23681 35127 23684
rect 35069 23675 35127 23681
rect 35434 23672 35440 23684
rect 35492 23672 35498 23724
rect 36262 23672 36268 23724
rect 36320 23672 36326 23724
rect 36449 23715 36507 23721
rect 36449 23681 36461 23715
rect 36495 23681 36507 23715
rect 36449 23675 36507 23681
rect 37093 23715 37151 23721
rect 37093 23681 37105 23715
rect 37139 23712 37151 23715
rect 37274 23712 37280 23724
rect 37139 23684 37280 23712
rect 37139 23681 37151 23684
rect 37093 23675 37151 23681
rect 30156 23616 30696 23644
rect 30156 23604 30162 23616
rect 26936 23548 28212 23576
rect 26936 23536 26942 23548
rect 21821 23511 21879 23517
rect 21821 23508 21833 23511
rect 20824 23480 21833 23508
rect 21821 23477 21833 23480
rect 21867 23477 21879 23511
rect 21821 23471 21879 23477
rect 23934 23468 23940 23520
rect 23992 23508 23998 23520
rect 24213 23511 24271 23517
rect 24213 23508 24225 23511
rect 23992 23480 24225 23508
rect 23992 23468 23998 23480
rect 24213 23477 24225 23480
rect 24259 23477 24271 23511
rect 24213 23471 24271 23477
rect 24486 23468 24492 23520
rect 24544 23468 24550 23520
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25225 23511 25283 23517
rect 25225 23508 25237 23511
rect 25004 23480 25237 23508
rect 25004 23468 25010 23480
rect 25225 23477 25237 23480
rect 25271 23477 25283 23511
rect 25225 23471 25283 23477
rect 26602 23468 26608 23520
rect 26660 23508 26666 23520
rect 27798 23508 27804 23520
rect 26660 23480 27804 23508
rect 26660 23468 26666 23480
rect 27798 23468 27804 23480
rect 27856 23508 27862 23520
rect 28077 23511 28135 23517
rect 28077 23508 28089 23511
rect 27856 23480 28089 23508
rect 27856 23468 27862 23480
rect 28077 23477 28089 23480
rect 28123 23477 28135 23511
rect 36464 23508 36492 23675
rect 37274 23672 37280 23684
rect 37332 23672 37338 23724
rect 37458 23672 37464 23724
rect 37516 23672 37522 23724
rect 37553 23715 37611 23721
rect 37553 23681 37565 23715
rect 37599 23681 37611 23715
rect 37553 23675 37611 23681
rect 37645 23715 37703 23721
rect 37645 23681 37657 23715
rect 37691 23681 37703 23715
rect 37645 23675 37703 23681
rect 36630 23604 36636 23656
rect 36688 23644 36694 23656
rect 36725 23647 36783 23653
rect 36725 23644 36737 23647
rect 36688 23616 36737 23644
rect 36688 23604 36694 23616
rect 36725 23613 36737 23616
rect 36771 23613 36783 23647
rect 36725 23607 36783 23613
rect 36740 23576 36768 23607
rect 37568 23576 37596 23675
rect 36740 23548 37596 23576
rect 36817 23511 36875 23517
rect 36817 23508 36829 23511
rect 36464 23480 36829 23508
rect 28077 23471 28135 23477
rect 36817 23477 36829 23480
rect 36863 23508 36875 23511
rect 36906 23508 36912 23520
rect 36863 23480 36912 23508
rect 36863 23477 36875 23480
rect 36817 23471 36875 23477
rect 36906 23468 36912 23480
rect 36964 23508 36970 23520
rect 37660 23508 37688 23675
rect 36964 23480 37688 23508
rect 36964 23468 36970 23480
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1670 23264 1676 23316
rect 1728 23304 1734 23316
rect 2133 23307 2191 23313
rect 2133 23304 2145 23307
rect 1728 23276 2145 23304
rect 1728 23264 1734 23276
rect 2133 23273 2145 23276
rect 2179 23273 2191 23307
rect 2133 23267 2191 23273
rect 5166 23264 5172 23316
rect 5224 23264 5230 23316
rect 5353 23307 5411 23313
rect 5353 23273 5365 23307
rect 5399 23304 5411 23307
rect 6822 23304 6828 23316
rect 5399 23276 6828 23304
rect 5399 23273 5411 23276
rect 5353 23267 5411 23273
rect 3418 23236 3424 23248
rect 2746 23208 3424 23236
rect 2038 23060 2044 23112
rect 2096 23100 2102 23112
rect 2133 23103 2191 23109
rect 2133 23100 2145 23103
rect 2096 23072 2145 23100
rect 2096 23060 2102 23072
rect 2133 23069 2145 23072
rect 2179 23069 2191 23103
rect 2133 23063 2191 23069
rect 2317 23103 2375 23109
rect 2317 23069 2329 23103
rect 2363 23100 2375 23103
rect 2746 23100 2774 23208
rect 3418 23196 3424 23208
rect 3476 23196 3482 23248
rect 4801 23239 4859 23245
rect 4801 23205 4813 23239
rect 4847 23205 4859 23239
rect 4801 23199 4859 23205
rect 4816 23168 4844 23199
rect 5920 23177 5948 23276
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 9214 23304 9220 23316
rect 8864 23276 9220 23304
rect 6454 23196 6460 23248
rect 6512 23236 6518 23248
rect 8754 23236 8760 23248
rect 6512 23208 8760 23236
rect 6512 23196 6518 23208
rect 8754 23196 8760 23208
rect 8812 23196 8818 23248
rect 3160 23140 4844 23168
rect 5905 23171 5963 23177
rect 2363 23072 2774 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 2958 23060 2964 23112
rect 3016 23060 3022 23112
rect 3160 23109 3188 23140
rect 5905 23137 5917 23171
rect 5951 23137 5963 23171
rect 5905 23131 5963 23137
rect 3145 23103 3203 23109
rect 3145 23069 3157 23103
rect 3191 23069 3203 23103
rect 3145 23063 3203 23069
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 4065 23103 4123 23109
rect 4065 23100 4077 23103
rect 4028 23072 4077 23100
rect 4028 23060 4034 23072
rect 4065 23069 4077 23072
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 4890 23060 4896 23112
rect 4948 23100 4954 23112
rect 5077 23103 5135 23109
rect 5077 23100 5089 23103
rect 4948 23072 5089 23100
rect 4948 23060 4954 23072
rect 5077 23069 5089 23072
rect 5123 23100 5135 23103
rect 5166 23100 5172 23112
rect 5123 23072 5172 23100
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 5166 23060 5172 23072
rect 5224 23060 5230 23112
rect 5718 23100 5724 23112
rect 5460 23072 5724 23100
rect 4709 23035 4767 23041
rect 4709 23001 4721 23035
rect 4755 23032 4767 23035
rect 4801 23035 4859 23041
rect 4801 23032 4813 23035
rect 4755 23004 4813 23032
rect 4755 23001 4767 23004
rect 4709 22995 4767 23001
rect 4801 23001 4813 23004
rect 4847 23001 4859 23035
rect 4801 22995 4859 23001
rect 5337 23035 5395 23041
rect 5337 23001 5349 23035
rect 5383 23032 5395 23035
rect 5460 23032 5488 23072
rect 5718 23060 5724 23072
rect 5776 23060 5782 23112
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23069 5871 23103
rect 5813 23063 5871 23069
rect 5383 23004 5488 23032
rect 5537 23035 5595 23041
rect 5383 23001 5395 23004
rect 5337 22995 5395 23001
rect 5537 23001 5549 23035
rect 5583 23032 5595 23035
rect 5828 23032 5856 23063
rect 5994 23060 6000 23112
rect 6052 23060 6058 23112
rect 6086 23060 6092 23112
rect 6144 23100 6150 23112
rect 6362 23100 6368 23112
rect 6144 23072 6368 23100
rect 6144 23060 6150 23072
rect 6362 23060 6368 23072
rect 6420 23060 6426 23112
rect 6454 23060 6460 23112
rect 6512 23060 6518 23112
rect 6638 23060 6644 23112
rect 6696 23060 6702 23112
rect 6733 23103 6791 23109
rect 6733 23069 6745 23103
rect 6779 23069 6791 23103
rect 6733 23063 6791 23069
rect 6178 23032 6184 23044
rect 5583 23004 5764 23032
rect 5828 23004 6184 23032
rect 5583 23001 5595 23004
rect 5537 22995 5595 23001
rect 5736 22976 5764 23004
rect 6178 22992 6184 23004
rect 6236 23032 6242 23044
rect 6748 23032 6776 23063
rect 6822 23060 6828 23112
rect 6880 23060 6886 23112
rect 8297 23103 8355 23109
rect 8297 23069 8309 23103
rect 8343 23100 8355 23103
rect 8478 23100 8484 23112
rect 8343 23072 8484 23100
rect 8343 23069 8355 23072
rect 8297 23063 8355 23069
rect 8478 23060 8484 23072
rect 8536 23060 8542 23112
rect 8573 23103 8631 23109
rect 8573 23069 8585 23103
rect 8619 23100 8631 23103
rect 8864 23100 8892 23276
rect 9214 23264 9220 23276
rect 9272 23304 9278 23316
rect 10689 23307 10747 23313
rect 10689 23304 10701 23307
rect 9272 23276 10701 23304
rect 9272 23264 9278 23276
rect 10689 23273 10701 23276
rect 10735 23273 10747 23307
rect 10689 23267 10747 23273
rect 18598 23264 18604 23316
rect 18656 23304 18662 23316
rect 18693 23307 18751 23313
rect 18693 23304 18705 23307
rect 18656 23276 18705 23304
rect 18656 23264 18662 23276
rect 18693 23273 18705 23276
rect 18739 23273 18751 23307
rect 18693 23267 18751 23273
rect 20530 23264 20536 23316
rect 20588 23264 20594 23316
rect 28077 23307 28135 23313
rect 28077 23273 28089 23307
rect 28123 23304 28135 23307
rect 28166 23304 28172 23316
rect 28123 23276 28172 23304
rect 28123 23273 28135 23276
rect 28077 23267 28135 23273
rect 28166 23264 28172 23276
rect 28224 23264 28230 23316
rect 28258 23264 28264 23316
rect 28316 23264 28322 23316
rect 31481 23307 31539 23313
rect 31481 23273 31493 23307
rect 31527 23304 31539 23307
rect 31570 23304 31576 23316
rect 31527 23276 31576 23304
rect 31527 23273 31539 23276
rect 31481 23267 31539 23273
rect 31570 23264 31576 23276
rect 31628 23264 31634 23316
rect 32122 23264 32128 23316
rect 32180 23264 32186 23316
rect 32953 23307 33011 23313
rect 32953 23273 32965 23307
rect 32999 23304 33011 23307
rect 33042 23304 33048 23316
rect 32999 23276 33048 23304
rect 32999 23273 33011 23276
rect 32953 23267 33011 23273
rect 33042 23264 33048 23276
rect 33100 23264 33106 23316
rect 36262 23264 36268 23316
rect 36320 23304 36326 23316
rect 36357 23307 36415 23313
rect 36357 23304 36369 23307
rect 36320 23276 36369 23304
rect 36320 23264 36326 23276
rect 36357 23273 36369 23276
rect 36403 23273 36415 23307
rect 36357 23267 36415 23273
rect 36906 23264 36912 23316
rect 36964 23264 36970 23316
rect 37274 23264 37280 23316
rect 37332 23304 37338 23316
rect 37645 23307 37703 23313
rect 37645 23304 37657 23307
rect 37332 23276 37657 23304
rect 37332 23264 37338 23276
rect 37645 23273 37657 23276
rect 37691 23273 37703 23307
rect 37645 23267 37703 23273
rect 21910 23236 21916 23248
rect 16776 23208 21916 23236
rect 8941 23171 8999 23177
rect 8941 23137 8953 23171
rect 8987 23168 8999 23171
rect 10226 23168 10232 23180
rect 8987 23140 10232 23168
rect 8987 23137 8999 23140
rect 8941 23131 8999 23137
rect 10226 23128 10232 23140
rect 10284 23168 10290 23180
rect 10502 23168 10508 23180
rect 10284 23140 10508 23168
rect 10284 23128 10290 23140
rect 10502 23128 10508 23140
rect 10560 23128 10566 23180
rect 16393 23171 16451 23177
rect 16393 23137 16405 23171
rect 16439 23168 16451 23171
rect 16776 23168 16804 23208
rect 21910 23196 21916 23208
rect 21968 23196 21974 23248
rect 23198 23196 23204 23248
rect 23256 23236 23262 23248
rect 23937 23239 23995 23245
rect 23937 23236 23949 23239
rect 23256 23208 23949 23236
rect 23256 23196 23262 23208
rect 23937 23205 23949 23208
rect 23983 23205 23995 23239
rect 27890 23236 27896 23248
rect 23937 23199 23995 23205
rect 26988 23208 27896 23236
rect 16439 23140 16804 23168
rect 16439 23137 16451 23140
rect 16393 23131 16451 23137
rect 8619 23072 8892 23100
rect 8619 23069 8631 23072
rect 8573 23063 8631 23069
rect 16022 23060 16028 23112
rect 16080 23100 16086 23112
rect 16408 23100 16436 23131
rect 17678 23128 17684 23180
rect 17736 23168 17742 23180
rect 18601 23171 18659 23177
rect 18601 23168 18613 23171
rect 17736 23140 18613 23168
rect 17736 23128 17742 23140
rect 18601 23137 18613 23140
rect 18647 23168 18659 23171
rect 18782 23168 18788 23180
rect 18647 23140 18788 23168
rect 18647 23137 18659 23140
rect 18601 23131 18659 23137
rect 18782 23128 18788 23140
rect 18840 23128 18846 23180
rect 19797 23171 19855 23177
rect 19797 23137 19809 23171
rect 19843 23168 19855 23171
rect 19843 23140 20392 23168
rect 19843 23137 19855 23140
rect 19797 23131 19855 23137
rect 16080 23072 16436 23100
rect 16080 23060 16086 23072
rect 18874 23060 18880 23112
rect 18932 23060 18938 23112
rect 19334 23060 19340 23112
rect 19392 23060 19398 23112
rect 19610 23060 19616 23112
rect 19668 23060 19674 23112
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 6236 23004 6776 23032
rect 6236 22992 6242 23004
rect 9214 22992 9220 23044
rect 9272 22992 9278 23044
rect 9674 22992 9680 23044
rect 9732 22992 9738 23044
rect 16209 23035 16267 23041
rect 16209 23001 16221 23035
rect 16255 23032 16267 23035
rect 16574 23032 16580 23044
rect 16255 23004 16580 23032
rect 16255 23001 16267 23004
rect 16209 22995 16267 23001
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 19061 23035 19119 23041
rect 19061 23001 19073 23035
rect 19107 23032 19119 23035
rect 19904 23032 19932 23063
rect 19978 23060 19984 23112
rect 20036 23060 20042 23112
rect 20070 23060 20076 23112
rect 20128 23100 20134 23112
rect 20364 23109 20392 23140
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 21269 23171 21327 23177
rect 21269 23168 21281 23171
rect 20864 23140 21281 23168
rect 20864 23128 20870 23140
rect 21269 23137 21281 23140
rect 21315 23137 21327 23171
rect 22830 23168 22836 23180
rect 21269 23131 21327 23137
rect 22112 23140 22836 23168
rect 20165 23103 20223 23109
rect 20165 23100 20177 23103
rect 20128 23072 20177 23100
rect 20128 23060 20134 23072
rect 20165 23069 20177 23072
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 20349 23103 20407 23109
rect 20349 23069 20361 23103
rect 20395 23069 20407 23103
rect 20349 23063 20407 23069
rect 21082 23060 21088 23112
rect 21140 23060 21146 23112
rect 19107 23004 19932 23032
rect 20257 23035 20315 23041
rect 19107 23001 19119 23004
rect 19061 22995 19119 23001
rect 20257 23001 20269 23035
rect 20303 23032 20315 23035
rect 20990 23032 20996 23044
rect 20303 23004 20996 23032
rect 20303 23001 20315 23004
rect 20257 22995 20315 23001
rect 20990 22992 20996 23004
rect 21048 22992 21054 23044
rect 21284 23032 21312 23131
rect 22112 23109 22140 23140
rect 22830 23128 22836 23140
rect 22888 23128 22894 23180
rect 24394 23128 24400 23180
rect 24452 23168 24458 23180
rect 26234 23168 26240 23180
rect 24452 23140 26240 23168
rect 24452 23128 24458 23140
rect 26234 23128 26240 23140
rect 26292 23128 26298 23180
rect 22097 23103 22155 23109
rect 22097 23069 22109 23103
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23069 22247 23103
rect 22189 23063 22247 23069
rect 22204 23032 22232 23063
rect 23934 23060 23940 23112
rect 23992 23060 23998 23112
rect 24213 23103 24271 23109
rect 24213 23069 24225 23103
rect 24259 23100 24271 23103
rect 24302 23100 24308 23112
rect 24259 23072 24308 23100
rect 24259 23069 24271 23072
rect 24213 23063 24271 23069
rect 24302 23060 24308 23072
rect 24360 23060 24366 23112
rect 26418 23060 26424 23112
rect 26476 23060 26482 23112
rect 26602 23060 26608 23112
rect 26660 23100 26666 23112
rect 26697 23103 26755 23109
rect 26697 23100 26709 23103
rect 26660 23072 26709 23100
rect 26660 23060 26666 23072
rect 26697 23069 26709 23072
rect 26743 23069 26755 23103
rect 26697 23063 26755 23069
rect 26786 23060 26792 23112
rect 26844 23100 26850 23112
rect 26988 23109 27016 23208
rect 27890 23196 27896 23208
rect 27948 23196 27954 23248
rect 30098 23196 30104 23248
rect 30156 23196 30162 23248
rect 37458 23196 37464 23248
rect 37516 23236 37522 23248
rect 37829 23239 37887 23245
rect 37829 23236 37841 23239
rect 37516 23208 37841 23236
rect 37516 23196 37522 23208
rect 37829 23205 37841 23208
rect 37875 23205 37887 23239
rect 37829 23199 37887 23205
rect 27341 23171 27399 23177
rect 27341 23137 27353 23171
rect 27387 23168 27399 23171
rect 28169 23171 28227 23177
rect 28169 23168 28181 23171
rect 27387 23140 28181 23168
rect 27387 23137 27399 23140
rect 27341 23131 27399 23137
rect 26881 23103 26939 23109
rect 26881 23100 26893 23103
rect 26844 23072 26893 23100
rect 26844 23060 26850 23072
rect 26881 23069 26893 23072
rect 26927 23069 26939 23103
rect 26881 23063 26939 23069
rect 26973 23103 27031 23109
rect 26973 23069 26985 23103
rect 27019 23069 27031 23103
rect 26973 23063 27031 23069
rect 27065 23103 27123 23109
rect 27065 23069 27077 23103
rect 27111 23100 27123 23103
rect 27111 23072 27200 23100
rect 27111 23069 27123 23072
rect 27065 23063 27123 23069
rect 21284 23004 22232 23032
rect 24673 23035 24731 23041
rect 24673 23001 24685 23035
rect 24719 23032 24731 23035
rect 24946 23032 24952 23044
rect 24719 23004 24952 23032
rect 24719 23001 24731 23004
rect 24673 22995 24731 23001
rect 24946 22992 24952 23004
rect 25004 22992 25010 23044
rect 25406 22992 25412 23044
rect 25464 22992 25470 23044
rect 2314 22924 2320 22976
rect 2372 22964 2378 22976
rect 3053 22967 3111 22973
rect 3053 22964 3065 22967
rect 2372 22936 3065 22964
rect 2372 22924 2378 22936
rect 3053 22933 3065 22936
rect 3099 22933 3111 22967
rect 3053 22927 3111 22933
rect 3142 22924 3148 22976
rect 3200 22964 3206 22976
rect 4062 22964 4068 22976
rect 3200 22936 4068 22964
rect 3200 22924 3206 22936
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 4985 22967 5043 22973
rect 4985 22933 4997 22967
rect 5031 22964 5043 22967
rect 5166 22964 5172 22976
rect 5031 22936 5172 22964
rect 5031 22933 5043 22936
rect 4985 22927 5043 22933
rect 5166 22924 5172 22936
rect 5224 22924 5230 22976
rect 5626 22924 5632 22976
rect 5684 22924 5690 22976
rect 5718 22924 5724 22976
rect 5776 22924 5782 22976
rect 7006 22924 7012 22976
rect 7064 22964 7070 22976
rect 7101 22967 7159 22973
rect 7101 22964 7113 22967
rect 7064 22936 7113 22964
rect 7064 22924 7070 22936
rect 7101 22933 7113 22936
rect 7147 22933 7159 22967
rect 7101 22927 7159 22933
rect 8389 22967 8447 22973
rect 8389 22933 8401 22967
rect 8435 22964 8447 22967
rect 8570 22964 8576 22976
rect 8435 22936 8576 22964
rect 8435 22933 8447 22936
rect 8389 22927 8447 22933
rect 8570 22924 8576 22936
rect 8628 22924 8634 22976
rect 8662 22924 8668 22976
rect 8720 22964 8726 22976
rect 8757 22967 8815 22973
rect 8757 22964 8769 22967
rect 8720 22936 8769 22964
rect 8720 22924 8726 22936
rect 8757 22933 8769 22936
rect 8803 22933 8815 22967
rect 8757 22927 8815 22933
rect 12066 22924 12072 22976
rect 12124 22924 12130 22976
rect 15746 22924 15752 22976
rect 15804 22924 15810 22976
rect 16114 22924 16120 22976
rect 16172 22924 16178 22976
rect 18138 22924 18144 22976
rect 18196 22964 18202 22976
rect 19242 22964 19248 22976
rect 18196 22936 19248 22964
rect 18196 22924 18202 22936
rect 19242 22924 19248 22936
rect 19300 22964 19306 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 19300 22936 19441 22964
rect 19300 22924 19306 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 19429 22927 19487 22933
rect 24121 22967 24179 22973
rect 24121 22933 24133 22967
rect 24167 22964 24179 22967
rect 24486 22964 24492 22976
rect 24167 22936 24492 22964
rect 24167 22933 24179 22936
rect 24121 22927 24179 22933
rect 24486 22924 24492 22936
rect 24544 22924 24550 22976
rect 27172 22964 27200 23072
rect 27246 23060 27252 23112
rect 27304 23102 27310 23112
rect 27540 23109 27568 23140
rect 28169 23137 28181 23140
rect 28215 23137 28227 23171
rect 28169 23131 28227 23137
rect 29825 23171 29883 23177
rect 29825 23137 29837 23171
rect 29871 23168 29883 23171
rect 30282 23168 30288 23180
rect 29871 23140 30288 23168
rect 29871 23137 29883 23140
rect 29825 23131 29883 23137
rect 30282 23128 30288 23140
rect 30340 23128 30346 23180
rect 31680 23140 32168 23168
rect 27433 23103 27491 23109
rect 27304 23100 27384 23102
rect 27433 23100 27445 23103
rect 27304 23074 27445 23100
rect 27304 23060 27310 23074
rect 27356 23072 27445 23074
rect 27433 23069 27445 23072
rect 27479 23069 27491 23103
rect 27433 23063 27491 23069
rect 27525 23103 27583 23109
rect 27525 23069 27537 23103
rect 27571 23069 27583 23103
rect 27525 23063 27583 23069
rect 27798 23060 27804 23112
rect 27856 23060 27862 23112
rect 27890 23060 27896 23112
rect 27948 23060 27954 23112
rect 28350 23060 28356 23112
rect 28408 23060 28414 23112
rect 28442 23060 28448 23112
rect 28500 23060 28506 23112
rect 28534 23060 28540 23112
rect 28592 23060 28598 23112
rect 29733 23103 29791 23109
rect 29733 23069 29745 23103
rect 29779 23100 29791 23103
rect 30834 23100 30840 23112
rect 29779 23072 30840 23100
rect 29779 23069 29791 23072
rect 29733 23063 29791 23069
rect 30834 23060 30840 23072
rect 30892 23060 30898 23112
rect 31680 23109 31708 23140
rect 32140 23112 32168 23140
rect 36630 23128 36636 23180
rect 36688 23168 36694 23180
rect 36817 23171 36875 23177
rect 36817 23168 36829 23171
rect 36688 23140 36829 23168
rect 36688 23128 36694 23140
rect 36817 23137 36829 23140
rect 36863 23137 36875 23171
rect 36817 23131 36875 23137
rect 31665 23103 31723 23109
rect 31665 23069 31677 23103
rect 31711 23069 31723 23103
rect 31665 23063 31723 23069
rect 31754 23060 31760 23112
rect 31812 23100 31818 23112
rect 31941 23103 31999 23109
rect 31941 23100 31953 23103
rect 31812 23072 31953 23100
rect 31812 23060 31818 23072
rect 31941 23069 31953 23072
rect 31987 23069 31999 23103
rect 31941 23063 31999 23069
rect 32122 23060 32128 23112
rect 32180 23060 32186 23112
rect 33134 23060 33140 23112
rect 33192 23060 33198 23112
rect 33226 23060 33232 23112
rect 33284 23060 33290 23112
rect 36541 23103 36599 23109
rect 36541 23069 36553 23103
rect 36587 23069 36599 23103
rect 36541 23063 36599 23069
rect 27709 23035 27767 23041
rect 27709 23001 27721 23035
rect 27755 23032 27767 23035
rect 28629 23035 28687 23041
rect 28629 23032 28641 23035
rect 27755 23004 28641 23032
rect 27755 23001 27767 23004
rect 27709 22995 27767 23001
rect 28629 23001 28641 23004
rect 28675 23001 28687 23035
rect 36556 23032 36584 23063
rect 36722 23060 36728 23112
rect 36780 23060 36786 23112
rect 36906 23060 36912 23112
rect 36964 23060 36970 23112
rect 37093 23103 37151 23109
rect 37093 23069 37105 23103
rect 37139 23069 37151 23103
rect 37093 23063 37151 23069
rect 36924 23032 36952 23060
rect 36556 23004 36952 23032
rect 37108 23032 37136 23063
rect 37182 23060 37188 23112
rect 37240 23100 37246 23112
rect 37366 23100 37372 23112
rect 37240 23072 37372 23100
rect 37240 23060 37246 23072
rect 37366 23060 37372 23072
rect 37424 23060 37430 23112
rect 37461 23103 37519 23109
rect 37461 23069 37473 23103
rect 37507 23100 37519 23103
rect 37642 23100 37648 23112
rect 37507 23072 37648 23100
rect 37507 23069 37519 23072
rect 37461 23063 37519 23069
rect 37642 23060 37648 23072
rect 37700 23060 37706 23112
rect 37918 23060 37924 23112
rect 37976 23060 37982 23112
rect 37108 23004 37320 23032
rect 28629 22995 28687 23001
rect 27724 22964 27752 22995
rect 37292 22973 37320 23004
rect 27172 22936 27752 22964
rect 37277 22967 37335 22973
rect 37277 22933 37289 22967
rect 37323 22964 37335 22967
rect 37366 22964 37372 22976
rect 37323 22936 37372 22964
rect 37323 22933 37335 22936
rect 37277 22927 37335 22933
rect 37366 22924 37372 22936
rect 37424 22964 37430 22976
rect 38102 22964 38108 22976
rect 37424 22936 38108 22964
rect 37424 22924 37430 22936
rect 38102 22924 38108 22936
rect 38160 22924 38166 22976
rect 1104 22874 38824 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 38824 22874
rect 1104 22800 38824 22822
rect 5626 22720 5632 22772
rect 5684 22760 5690 22772
rect 5684 22732 6776 22760
rect 5684 22720 5690 22732
rect 2314 22652 2320 22704
rect 2372 22652 2378 22704
rect 3050 22652 3056 22704
rect 3108 22652 3114 22704
rect 4062 22652 4068 22704
rect 4120 22692 4126 22704
rect 6457 22695 6515 22701
rect 4120 22664 4646 22692
rect 5736 22664 6408 22692
rect 4120 22652 4126 22664
rect 5736 22624 5764 22664
rect 5368 22596 5764 22624
rect 5813 22627 5871 22633
rect 1394 22516 1400 22568
rect 1452 22556 1458 22568
rect 2038 22556 2044 22568
rect 1452 22528 2044 22556
rect 1452 22516 1458 22528
rect 2038 22516 2044 22528
rect 2096 22556 2102 22568
rect 3878 22556 3884 22568
rect 2096 22528 3884 22556
rect 2096 22516 2102 22528
rect 3878 22516 3884 22528
rect 3936 22516 3942 22568
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22556 4215 22559
rect 4706 22556 4712 22568
rect 4203 22528 4712 22556
rect 4203 22525 4215 22528
rect 4157 22519 4215 22525
rect 4706 22516 4712 22528
rect 4764 22516 4770 22568
rect 4798 22516 4804 22568
rect 4856 22556 4862 22568
rect 5368 22556 5396 22596
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 5902 22624 5908 22636
rect 5859 22596 5908 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 5902 22584 5908 22596
rect 5960 22584 5966 22636
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6380 22633 6408 22664
rect 6457 22661 6469 22695
rect 6503 22692 6515 22695
rect 6638 22692 6644 22704
rect 6503 22664 6644 22692
rect 6503 22661 6515 22664
rect 6457 22655 6515 22661
rect 6638 22652 6644 22664
rect 6696 22652 6702 22704
rect 6748 22633 6776 22732
rect 6822 22720 6828 22772
rect 6880 22760 6886 22772
rect 8386 22760 8392 22772
rect 6880 22732 8392 22760
rect 6880 22720 6886 22732
rect 8386 22720 8392 22732
rect 8444 22760 8450 22772
rect 8481 22763 8539 22769
rect 8481 22760 8493 22763
rect 8444 22732 8493 22760
rect 8444 22720 8450 22732
rect 8481 22729 8493 22732
rect 8527 22729 8539 22763
rect 8481 22723 8539 22729
rect 8754 22720 8760 22772
rect 8812 22760 8818 22772
rect 8865 22763 8923 22769
rect 8865 22760 8877 22763
rect 8812 22732 8877 22760
rect 8812 22720 8818 22732
rect 8865 22729 8877 22732
rect 8911 22729 8923 22763
rect 8865 22723 8923 22729
rect 9033 22763 9091 22769
rect 9033 22729 9045 22763
rect 9079 22760 9091 22763
rect 9214 22760 9220 22772
rect 9079 22732 9220 22760
rect 9079 22729 9091 22732
rect 9033 22723 9091 22729
rect 9214 22720 9220 22732
rect 9272 22720 9278 22772
rect 11701 22763 11759 22769
rect 11701 22729 11713 22763
rect 11747 22760 11759 22763
rect 11790 22760 11796 22772
rect 11747 22732 11796 22760
rect 11747 22729 11759 22732
rect 11701 22723 11759 22729
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 12345 22763 12403 22769
rect 12345 22760 12357 22763
rect 11992 22732 12357 22760
rect 7006 22652 7012 22704
rect 7064 22652 7070 22704
rect 8018 22652 8024 22704
rect 8076 22652 8082 22704
rect 8662 22652 8668 22704
rect 8720 22652 8726 22704
rect 11992 22701 12020 22732
rect 12345 22729 12357 22732
rect 12391 22760 12403 22763
rect 12621 22763 12679 22769
rect 12621 22760 12633 22763
rect 12391 22732 12633 22760
rect 12391 22729 12403 22732
rect 12345 22723 12403 22729
rect 12621 22729 12633 22732
rect 12667 22760 12679 22763
rect 12805 22763 12863 22769
rect 12805 22760 12817 22763
rect 12667 22732 12817 22760
rect 12667 22729 12679 22732
rect 12621 22723 12679 22729
rect 12805 22729 12817 22732
rect 12851 22760 12863 22763
rect 14550 22760 14556 22772
rect 12851 22732 14556 22760
rect 12851 22729 12863 22732
rect 12805 22723 12863 22729
rect 14550 22720 14556 22732
rect 14608 22720 14614 22772
rect 19337 22763 19395 22769
rect 19337 22729 19349 22763
rect 19383 22760 19395 22763
rect 19610 22760 19616 22772
rect 19383 22732 19616 22760
rect 19383 22729 19395 22732
rect 19337 22723 19395 22729
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 19978 22720 19984 22772
rect 20036 22760 20042 22772
rect 20257 22763 20315 22769
rect 20257 22760 20269 22763
rect 20036 22732 20269 22760
rect 20036 22720 20042 22732
rect 20257 22729 20269 22732
rect 20303 22729 20315 22763
rect 20257 22723 20315 22729
rect 11977 22695 12035 22701
rect 11977 22661 11989 22695
rect 12023 22661 12035 22695
rect 11977 22655 12035 22661
rect 18782 22652 18788 22704
rect 18840 22692 18846 22704
rect 20272 22692 20300 22723
rect 20990 22720 20996 22772
rect 21048 22720 21054 22772
rect 21913 22763 21971 22769
rect 21913 22729 21925 22763
rect 21959 22760 21971 22763
rect 22278 22760 22284 22772
rect 21959 22732 22284 22760
rect 21959 22729 21971 22732
rect 21913 22723 21971 22729
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 25317 22763 25375 22769
rect 25317 22729 25329 22763
rect 25363 22760 25375 22763
rect 25498 22760 25504 22772
rect 25363 22732 25504 22760
rect 25363 22729 25375 22732
rect 25317 22723 25375 22729
rect 25498 22720 25504 22732
rect 25556 22720 25562 22772
rect 26786 22720 26792 22772
rect 26844 22720 26850 22772
rect 27617 22763 27675 22769
rect 27617 22729 27629 22763
rect 27663 22760 27675 22763
rect 27706 22760 27712 22772
rect 27663 22732 27712 22760
rect 27663 22729 27675 22732
rect 27617 22723 27675 22729
rect 27706 22720 27712 22732
rect 27764 22720 27770 22772
rect 28810 22720 28816 22772
rect 28868 22760 28874 22772
rect 28905 22763 28963 22769
rect 28905 22760 28917 22763
rect 28868 22732 28917 22760
rect 28868 22720 28874 22732
rect 28905 22729 28917 22732
rect 28951 22729 28963 22763
rect 28905 22723 28963 22729
rect 29362 22720 29368 22772
rect 29420 22720 29426 22772
rect 30190 22720 30196 22772
rect 30248 22720 30254 22772
rect 30282 22720 30288 22772
rect 30340 22720 30346 22772
rect 30834 22720 30840 22772
rect 30892 22720 30898 22772
rect 32122 22720 32128 22772
rect 32180 22720 32186 22772
rect 32585 22763 32643 22769
rect 32585 22729 32597 22763
rect 32631 22760 32643 22763
rect 33226 22760 33232 22772
rect 32631 22732 33232 22760
rect 32631 22729 32643 22732
rect 32585 22723 32643 22729
rect 33226 22720 33232 22732
rect 33284 22760 33290 22772
rect 33873 22763 33931 22769
rect 33284 22732 33732 22760
rect 33284 22720 33290 22732
rect 21358 22692 21364 22704
rect 18840 22664 19472 22692
rect 20272 22664 21364 22692
rect 18840 22652 18846 22664
rect 6365 22627 6423 22633
rect 6365 22593 6377 22627
rect 6411 22593 6423 22627
rect 6365 22587 6423 22593
rect 6733 22627 6791 22633
rect 6733 22593 6745 22627
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 12066 22624 12072 22636
rect 11388 22596 12072 22624
rect 11388 22584 11394 22596
rect 12066 22584 12072 22596
rect 12124 22624 12130 22636
rect 12161 22627 12219 22633
rect 12161 22624 12173 22627
rect 12124 22596 12173 22624
rect 12124 22584 12130 22596
rect 12161 22593 12173 22596
rect 12207 22593 12219 22627
rect 12161 22587 12219 22593
rect 19150 22584 19156 22636
rect 19208 22624 19214 22636
rect 19444 22633 19472 22664
rect 21358 22652 21364 22664
rect 21416 22692 21422 22704
rect 21416 22664 21864 22692
rect 21416 22652 21422 22664
rect 19251 22627 19309 22633
rect 19251 22624 19263 22627
rect 19208 22596 19263 22624
rect 19208 22584 19214 22596
rect 19251 22593 19263 22596
rect 19297 22593 19309 22627
rect 19251 22587 19309 22593
rect 19429 22627 19487 22633
rect 19429 22593 19441 22627
rect 19475 22624 19487 22627
rect 19705 22627 19763 22633
rect 19705 22624 19717 22627
rect 19475 22596 19717 22624
rect 19475 22593 19487 22596
rect 19429 22587 19487 22593
rect 19705 22593 19717 22596
rect 19751 22593 19763 22627
rect 19705 22587 19763 22593
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22624 20223 22627
rect 20254 22624 20260 22636
rect 20211 22596 20260 22624
rect 20211 22593 20223 22596
rect 20165 22587 20223 22593
rect 4856 22528 5396 22556
rect 4856 22516 4862 22528
rect 5718 22516 5724 22568
rect 5776 22556 5782 22568
rect 7466 22556 7472 22568
rect 5776 22528 7472 22556
rect 5776 22516 5782 22528
rect 7466 22516 7472 22528
rect 7524 22516 7530 22568
rect 13541 22559 13599 22565
rect 13541 22525 13553 22559
rect 13587 22556 13599 22559
rect 13722 22556 13728 22568
rect 13587 22528 13728 22556
rect 13587 22525 13599 22528
rect 13541 22519 13599 22525
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 19260 22556 19288 22587
rect 20254 22584 20260 22596
rect 20312 22584 20318 22636
rect 21836 22633 21864 22664
rect 23198 22652 23204 22704
rect 23256 22652 23262 22704
rect 23658 22652 23664 22704
rect 23716 22652 23722 22704
rect 24762 22652 24768 22704
rect 24820 22692 24826 22704
rect 24949 22695 25007 22701
rect 24949 22692 24961 22695
rect 24820 22664 24961 22692
rect 24820 22652 24826 22664
rect 24949 22661 24961 22664
rect 24995 22661 25007 22695
rect 24949 22655 25007 22661
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22624 20407 22627
rect 20625 22627 20683 22633
rect 20625 22624 20637 22627
rect 20395 22596 20637 22624
rect 20395 22593 20407 22596
rect 20349 22587 20407 22593
rect 20625 22593 20637 22596
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 19521 22559 19579 22565
rect 19521 22556 19533 22559
rect 19260 22528 19533 22556
rect 19521 22525 19533 22528
rect 19567 22525 19579 22559
rect 19521 22519 19579 22525
rect 18690 22448 18696 22500
rect 18748 22488 18754 22500
rect 20364 22488 20392 22587
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 25409 22627 25467 22633
rect 25409 22593 25421 22627
rect 25455 22593 25467 22627
rect 25516 22624 25544 22720
rect 28534 22692 28540 22704
rect 27632 22664 28540 22692
rect 26237 22627 26295 22633
rect 26237 22624 26249 22627
rect 25516 22596 26249 22624
rect 25409 22587 25467 22593
rect 26237 22593 26249 22596
rect 26283 22593 26295 22627
rect 26237 22587 26295 22593
rect 26513 22627 26571 22633
rect 26513 22593 26525 22627
rect 26559 22593 26571 22627
rect 26513 22587 26571 22593
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 18748 22460 20392 22488
rect 21836 22528 22293 22556
rect 18748 22448 18754 22460
rect 3789 22423 3847 22429
rect 3789 22389 3801 22423
rect 3835 22420 3847 22423
rect 3970 22420 3976 22432
rect 3835 22392 3976 22420
rect 3835 22389 3847 22392
rect 3789 22383 3847 22389
rect 3970 22380 3976 22392
rect 4028 22380 4034 22432
rect 5350 22380 5356 22432
rect 5408 22420 5414 22432
rect 5629 22423 5687 22429
rect 5629 22420 5641 22423
rect 5408 22392 5641 22420
rect 5408 22380 5414 22392
rect 5629 22389 5641 22392
rect 5675 22389 5687 22423
rect 5629 22383 5687 22389
rect 5902 22380 5908 22432
rect 5960 22420 5966 22432
rect 6181 22423 6239 22429
rect 6181 22420 6193 22423
rect 5960 22392 6193 22420
rect 5960 22380 5966 22392
rect 6181 22389 6193 22392
rect 6227 22389 6239 22423
rect 6181 22383 6239 22389
rect 8849 22423 8907 22429
rect 8849 22389 8861 22423
rect 8895 22420 8907 22423
rect 9582 22420 9588 22432
rect 8895 22392 9588 22420
rect 8895 22389 8907 22392
rect 8849 22383 8907 22389
rect 9582 22380 9588 22392
rect 9640 22380 9646 22432
rect 12897 22423 12955 22429
rect 12897 22389 12909 22423
rect 12943 22420 12955 22423
rect 12986 22420 12992 22432
rect 12943 22392 12992 22420
rect 12943 22389 12955 22392
rect 12897 22383 12955 22389
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19889 22423 19947 22429
rect 19889 22420 19901 22423
rect 19392 22392 19901 22420
rect 19392 22380 19398 22392
rect 19889 22389 19901 22392
rect 19935 22420 19947 22423
rect 20993 22423 21051 22429
rect 20993 22420 21005 22423
rect 19935 22392 21005 22420
rect 19935 22389 19947 22392
rect 19889 22383 19947 22389
rect 20993 22389 21005 22392
rect 21039 22389 21051 22423
rect 20993 22383 21051 22389
rect 21174 22380 21180 22432
rect 21232 22420 21238 22432
rect 21836 22420 21864 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 22281 22519 22339 22525
rect 22922 22516 22928 22568
rect 22980 22516 22986 22568
rect 25424 22556 25452 22587
rect 26418 22556 26424 22568
rect 25424 22528 26424 22556
rect 26418 22516 26424 22528
rect 26476 22516 26482 22568
rect 26528 22556 26556 22587
rect 26602 22584 26608 22636
rect 26660 22584 26666 22636
rect 27154 22584 27160 22636
rect 27212 22584 27218 22636
rect 27632 22624 27660 22664
rect 28534 22652 28540 22664
rect 28592 22652 28598 22704
rect 28721 22695 28779 22701
rect 28721 22661 28733 22695
rect 28767 22692 28779 22695
rect 28767 22664 29132 22692
rect 28767 22661 28779 22664
rect 28721 22655 28779 22661
rect 27264 22596 27660 22624
rect 27985 22627 28043 22633
rect 26694 22556 26700 22568
rect 26528 22528 26700 22556
rect 26694 22516 26700 22528
rect 26752 22556 26758 22568
rect 27264 22556 27292 22596
rect 27985 22593 27997 22627
rect 28031 22624 28043 22627
rect 28031 22596 28580 22624
rect 28031 22593 28043 22596
rect 27985 22587 28043 22593
rect 26752 22528 27292 22556
rect 26752 22516 26758 22528
rect 27338 22516 27344 22568
rect 27396 22516 27402 22568
rect 27525 22559 27583 22565
rect 27525 22525 27537 22559
rect 27571 22556 27583 22559
rect 27706 22556 27712 22568
rect 27571 22528 27712 22556
rect 27571 22525 27583 22528
rect 27525 22519 27583 22525
rect 27706 22516 27712 22528
rect 27764 22516 27770 22568
rect 28074 22516 28080 22568
rect 28132 22516 28138 22568
rect 28552 22556 28580 22596
rect 28626 22584 28632 22636
rect 28684 22584 28690 22636
rect 28813 22627 28871 22633
rect 28813 22593 28825 22627
rect 28859 22624 28871 22627
rect 28902 22624 28908 22636
rect 28859 22596 28908 22624
rect 28859 22593 28871 22596
rect 28813 22587 28871 22593
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 29104 22633 29132 22664
rect 29178 22652 29184 22704
rect 29236 22652 29242 22704
rect 29273 22695 29331 22701
rect 29273 22661 29285 22695
rect 29319 22692 29331 22695
rect 29380 22692 29408 22720
rect 33042 22692 33048 22704
rect 29319 22664 29408 22692
rect 30514 22664 30788 22692
rect 29319 22661 29331 22664
rect 29273 22655 29331 22661
rect 29089 22627 29147 22633
rect 29089 22593 29101 22627
rect 29135 22593 29147 22627
rect 29089 22587 29147 22593
rect 29411 22627 29469 22633
rect 29411 22593 29423 22627
rect 29457 22624 29469 22627
rect 30009 22627 30067 22633
rect 29457 22596 29868 22624
rect 29457 22593 29469 22596
rect 29411 22587 29469 22593
rect 28994 22556 29000 22568
rect 28552 22528 29000 22556
rect 28994 22516 29000 22528
rect 29052 22516 29058 22568
rect 29840 22565 29868 22596
rect 30009 22593 30021 22627
rect 30055 22624 30067 22627
rect 30374 22624 30380 22636
rect 30055 22596 30380 22624
rect 30055 22593 30067 22596
rect 30009 22587 30067 22593
rect 30374 22584 30380 22596
rect 30432 22624 30438 22636
rect 30514 22633 30542 22664
rect 30760 22633 30788 22664
rect 32508 22664 33048 22692
rect 30499 22630 30557 22633
rect 30484 22627 30557 22630
rect 30484 22624 30511 22627
rect 30432 22596 30511 22624
rect 30432 22584 30438 22596
rect 30499 22593 30511 22596
rect 30545 22593 30557 22627
rect 30499 22587 30557 22593
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22593 30711 22627
rect 30653 22587 30711 22593
rect 30745 22627 30803 22633
rect 30745 22593 30757 22627
rect 30791 22593 30803 22627
rect 30745 22587 30803 22593
rect 31021 22627 31079 22633
rect 31021 22593 31033 22627
rect 31067 22593 31079 22627
rect 31021 22587 31079 22593
rect 32125 22627 32183 22633
rect 32125 22593 32137 22627
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 29549 22559 29607 22565
rect 29549 22525 29561 22559
rect 29595 22556 29607 22559
rect 29733 22559 29791 22565
rect 29733 22556 29745 22559
rect 29595 22528 29745 22556
rect 29595 22525 29607 22528
rect 29549 22519 29607 22525
rect 29733 22525 29745 22528
rect 29779 22525 29791 22559
rect 29733 22519 29791 22525
rect 29825 22559 29883 22565
rect 29825 22525 29837 22559
rect 29871 22556 29883 22559
rect 30098 22556 30104 22568
rect 29871 22528 30104 22556
rect 29871 22525 29883 22528
rect 29825 22519 29883 22525
rect 22646 22488 22652 22500
rect 22296 22460 22652 22488
rect 21232 22392 21864 22420
rect 22189 22423 22247 22429
rect 21232 22380 21238 22392
rect 22189 22389 22201 22423
rect 22235 22420 22247 22423
rect 22296 22420 22324 22460
rect 22646 22448 22652 22460
rect 22704 22448 22710 22500
rect 26878 22448 26884 22500
rect 26936 22488 26942 22500
rect 27249 22491 27307 22497
rect 27249 22488 27261 22491
rect 26936 22460 27261 22488
rect 26936 22448 26942 22460
rect 27249 22457 27261 22460
rect 27295 22457 27307 22491
rect 27249 22451 27307 22457
rect 27430 22448 27436 22500
rect 27488 22488 27494 22500
rect 27488 22460 27752 22488
rect 27488 22448 27494 22460
rect 22235 22392 22324 22420
rect 22235 22389 22247 22392
rect 22189 22383 22247 22389
rect 22370 22380 22376 22432
rect 22428 22420 22434 22432
rect 22557 22423 22615 22429
rect 22557 22420 22569 22423
rect 22428 22392 22569 22420
rect 22428 22380 22434 22392
rect 22557 22389 22569 22392
rect 22603 22389 22615 22423
rect 22557 22383 22615 22389
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 24302 22420 24308 22432
rect 23716 22392 24308 22420
rect 23716 22380 23722 22392
rect 24302 22380 24308 22392
rect 24360 22380 24366 22432
rect 26329 22423 26387 22429
rect 26329 22389 26341 22423
rect 26375 22420 26387 22423
rect 26970 22420 26976 22432
rect 26375 22392 26976 22420
rect 26375 22389 26387 22392
rect 26329 22383 26387 22389
rect 26970 22380 26976 22392
rect 27028 22380 27034 22432
rect 27338 22380 27344 22432
rect 27396 22380 27402 22432
rect 27724 22420 27752 22460
rect 28810 22448 28816 22500
rect 28868 22488 28874 22500
rect 29564 22488 29592 22519
rect 30098 22516 30104 22528
rect 30156 22556 30162 22568
rect 30668 22556 30696 22587
rect 31036 22556 31064 22587
rect 30156 22528 31064 22556
rect 30156 22516 30162 22528
rect 32030 22516 32036 22568
rect 32088 22556 32094 22568
rect 32140 22556 32168 22587
rect 32306 22584 32312 22636
rect 32364 22584 32370 22636
rect 32508 22633 32536 22664
rect 33042 22652 33048 22664
rect 33100 22652 33106 22704
rect 32493 22627 32551 22633
rect 32493 22593 32505 22627
rect 32539 22593 32551 22627
rect 32493 22587 32551 22593
rect 32677 22627 32735 22633
rect 32677 22593 32689 22627
rect 32723 22624 32735 22627
rect 32858 22624 32864 22636
rect 32723 22596 32864 22624
rect 32723 22593 32735 22596
rect 32677 22587 32735 22593
rect 32858 22584 32864 22596
rect 32916 22584 32922 22636
rect 33704 22633 33732 22732
rect 33873 22729 33885 22763
rect 33919 22760 33931 22763
rect 34330 22760 34336 22772
rect 33919 22732 34336 22760
rect 33919 22729 33931 22732
rect 33873 22723 33931 22729
rect 34330 22720 34336 22732
rect 34388 22720 34394 22772
rect 34517 22763 34575 22769
rect 34517 22729 34529 22763
rect 34563 22760 34575 22763
rect 34606 22760 34612 22772
rect 34563 22732 34612 22760
rect 34563 22729 34575 22732
rect 34517 22723 34575 22729
rect 34606 22720 34612 22732
rect 34664 22720 34670 22772
rect 34790 22720 34796 22772
rect 34848 22720 34854 22772
rect 36081 22763 36139 22769
rect 36081 22729 36093 22763
rect 36127 22760 36139 22763
rect 36630 22760 36636 22772
rect 36127 22732 36636 22760
rect 36127 22729 36139 22732
rect 36081 22723 36139 22729
rect 36630 22720 36636 22732
rect 36688 22720 36694 22772
rect 36722 22720 36728 22772
rect 36780 22760 36786 22772
rect 36909 22763 36967 22769
rect 36909 22760 36921 22763
rect 36780 22732 36921 22760
rect 36780 22720 36786 22732
rect 36909 22729 36921 22732
rect 36955 22729 36967 22763
rect 36909 22723 36967 22729
rect 37826 22720 37832 22772
rect 37884 22720 37890 22772
rect 37918 22720 37924 22772
rect 37976 22720 37982 22772
rect 34945 22695 35003 22701
rect 34945 22692 34957 22695
rect 34440 22664 34957 22692
rect 34440 22636 34468 22664
rect 34945 22661 34957 22664
rect 34991 22692 35003 22695
rect 35161 22695 35219 22701
rect 34991 22664 35112 22692
rect 34991 22661 35003 22664
rect 34945 22655 35003 22661
rect 33137 22627 33195 22633
rect 33137 22593 33149 22627
rect 33183 22593 33195 22627
rect 33137 22587 33195 22593
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 33045 22559 33103 22565
rect 33045 22556 33057 22559
rect 32088 22528 33057 22556
rect 32088 22516 32094 22528
rect 33045 22525 33057 22528
rect 33091 22525 33103 22559
rect 33152 22556 33180 22587
rect 34422 22584 34428 22636
rect 34480 22584 34486 22636
rect 34606 22584 34612 22636
rect 34664 22584 34670 22636
rect 35084 22624 35112 22664
rect 35161 22661 35173 22695
rect 35207 22692 35219 22695
rect 37274 22692 37280 22704
rect 35207 22664 35572 22692
rect 35207 22661 35219 22664
rect 35161 22655 35219 22661
rect 35253 22627 35311 22633
rect 35253 22624 35265 22627
rect 35084 22596 35265 22624
rect 35253 22593 35265 22596
rect 35299 22593 35311 22627
rect 35253 22587 35311 22593
rect 35342 22584 35348 22636
rect 35400 22584 35406 22636
rect 35544 22633 35572 22664
rect 36280 22664 37280 22692
rect 35529 22627 35587 22633
rect 35529 22593 35541 22627
rect 35575 22624 35587 22627
rect 35894 22624 35900 22636
rect 35575 22596 35900 22624
rect 35575 22593 35587 22596
rect 35529 22587 35587 22593
rect 35894 22584 35900 22596
rect 35952 22584 35958 22636
rect 36280 22633 36308 22664
rect 37274 22652 37280 22664
rect 37332 22652 37338 22704
rect 35989 22627 36047 22633
rect 35989 22593 36001 22627
rect 36035 22593 36047 22627
rect 35989 22587 36047 22593
rect 36173 22627 36231 22633
rect 36173 22593 36185 22627
rect 36219 22593 36231 22627
rect 36173 22587 36231 22593
rect 36265 22627 36323 22633
rect 36265 22593 36277 22627
rect 36311 22593 36323 22627
rect 36265 22587 36323 22593
rect 33413 22559 33471 22565
rect 33413 22556 33425 22559
rect 33152 22528 33425 22556
rect 33045 22519 33103 22525
rect 33413 22525 33425 22528
rect 33459 22556 33471 22559
rect 33962 22556 33968 22568
rect 33459 22528 33968 22556
rect 33459 22525 33471 22528
rect 33413 22519 33471 22525
rect 28868 22460 29592 22488
rect 31021 22491 31079 22497
rect 28868 22448 28874 22460
rect 31021 22457 31033 22491
rect 31067 22488 31079 22491
rect 31754 22488 31760 22500
rect 31067 22460 31760 22488
rect 31067 22457 31079 22460
rect 31021 22451 31079 22457
rect 31754 22448 31760 22460
rect 31812 22448 31818 22500
rect 33060 22488 33088 22519
rect 33962 22516 33968 22528
rect 34020 22516 34026 22568
rect 33505 22491 33563 22497
rect 33505 22488 33517 22491
rect 33060 22460 33517 22488
rect 33505 22457 33517 22460
rect 33551 22457 33563 22491
rect 33505 22451 33563 22457
rect 35434 22448 35440 22500
rect 35492 22488 35498 22500
rect 35529 22491 35587 22497
rect 35529 22488 35541 22491
rect 35492 22460 35541 22488
rect 35492 22448 35498 22460
rect 35529 22457 35541 22460
rect 35575 22457 35587 22491
rect 36004 22488 36032 22587
rect 36188 22556 36216 22587
rect 36446 22584 36452 22636
rect 36504 22584 36510 22636
rect 36630 22584 36636 22636
rect 36688 22624 36694 22636
rect 36725 22627 36783 22633
rect 36725 22624 36737 22627
rect 36688 22596 36737 22624
rect 36688 22584 36694 22596
rect 36725 22593 36737 22596
rect 36771 22593 36783 22627
rect 36725 22587 36783 22593
rect 37550 22584 37556 22636
rect 37608 22624 37614 22636
rect 37645 22627 37703 22633
rect 37645 22624 37657 22627
rect 37608 22596 37657 22624
rect 37608 22584 37614 22596
rect 37645 22593 37657 22596
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 36357 22559 36415 22565
rect 36357 22556 36369 22559
rect 36188 22528 36369 22556
rect 36357 22525 36369 22528
rect 36403 22556 36415 22559
rect 36541 22559 36599 22565
rect 36541 22556 36553 22559
rect 36403 22528 36553 22556
rect 36403 22525 36415 22528
rect 36357 22519 36415 22525
rect 36541 22525 36553 22528
rect 36587 22525 36599 22559
rect 36541 22519 36599 22525
rect 37369 22559 37427 22565
rect 37369 22525 37381 22559
rect 37415 22556 37427 22559
rect 37458 22556 37464 22568
rect 37415 22528 37464 22556
rect 37415 22525 37427 22528
rect 37369 22519 37427 22525
rect 37458 22516 37464 22528
rect 37516 22516 37522 22568
rect 36630 22488 36636 22500
rect 36004 22460 36636 22488
rect 35529 22451 35587 22457
rect 36630 22448 36636 22460
rect 36688 22448 36694 22500
rect 37936 22488 37964 22720
rect 38010 22652 38016 22704
rect 38068 22701 38074 22704
rect 38068 22695 38131 22701
rect 38068 22661 38085 22695
rect 38119 22661 38131 22695
rect 38068 22655 38131 22661
rect 38289 22695 38347 22701
rect 38289 22661 38301 22695
rect 38335 22692 38347 22695
rect 38378 22692 38384 22704
rect 38335 22664 38384 22692
rect 38335 22661 38347 22664
rect 38289 22655 38347 22661
rect 38068 22652 38074 22655
rect 38378 22652 38384 22664
rect 38436 22652 38442 22704
rect 37476 22460 37964 22488
rect 29178 22420 29184 22432
rect 27724 22392 29184 22420
rect 29178 22380 29184 22392
rect 29236 22380 29242 22432
rect 32769 22423 32827 22429
rect 32769 22389 32781 22423
rect 32815 22420 32827 22423
rect 32858 22420 32864 22432
rect 32815 22392 32864 22420
rect 32815 22389 32827 22392
rect 32769 22383 32827 22389
rect 32858 22380 32864 22392
rect 32916 22380 32922 22432
rect 34977 22423 35035 22429
rect 34977 22389 34989 22423
rect 35023 22420 35035 22423
rect 35342 22420 35348 22432
rect 35023 22392 35348 22420
rect 35023 22389 35035 22392
rect 34977 22383 35035 22389
rect 35342 22380 35348 22392
rect 35400 22380 35406 22432
rect 37476 22429 37504 22460
rect 37461 22423 37519 22429
rect 37461 22389 37473 22423
rect 37507 22389 37519 22423
rect 37461 22383 37519 22389
rect 38102 22380 38108 22432
rect 38160 22380 38166 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 5166 22176 5172 22228
rect 5224 22216 5230 22228
rect 5353 22219 5411 22225
rect 5353 22216 5365 22219
rect 5224 22188 5365 22216
rect 5224 22176 5230 22188
rect 5353 22185 5365 22188
rect 5399 22216 5411 22219
rect 5442 22216 5448 22228
rect 5399 22188 5448 22216
rect 5399 22185 5411 22188
rect 5353 22179 5411 22185
rect 5442 22176 5448 22188
rect 5500 22216 5506 22228
rect 5902 22225 5908 22228
rect 5892 22219 5908 22225
rect 5500 22188 5764 22216
rect 5500 22176 5506 22188
rect 3878 22040 3884 22092
rect 3936 22080 3942 22092
rect 4341 22083 4399 22089
rect 4341 22080 4353 22083
rect 3936 22052 4353 22080
rect 3936 22040 3942 22052
rect 4341 22049 4353 22052
rect 4387 22080 4399 22083
rect 4614 22080 4620 22092
rect 4387 22052 4620 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 4614 22040 4620 22052
rect 4672 22080 4678 22092
rect 5736 22080 5764 22188
rect 5892 22185 5904 22219
rect 5892 22179 5908 22185
rect 5902 22176 5908 22179
rect 5960 22176 5966 22228
rect 7377 22219 7435 22225
rect 7377 22185 7389 22219
rect 7423 22216 7435 22219
rect 7466 22216 7472 22228
rect 7423 22188 7472 22216
rect 7423 22185 7435 22188
rect 7377 22179 7435 22185
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 14550 22216 14556 22228
rect 14332 22188 14556 22216
rect 14332 22176 14338 22188
rect 14550 22176 14556 22188
rect 14608 22216 14614 22228
rect 14921 22219 14979 22225
rect 14921 22216 14933 22219
rect 14608 22188 14933 22216
rect 14608 22176 14614 22188
rect 14921 22185 14933 22188
rect 14967 22216 14979 22219
rect 15102 22216 15108 22228
rect 14967 22188 15108 22216
rect 14967 22185 14979 22188
rect 14921 22179 14979 22185
rect 15102 22176 15108 22188
rect 15160 22176 15166 22228
rect 15368 22219 15426 22225
rect 15368 22185 15380 22219
rect 15414 22216 15426 22219
rect 15746 22216 15752 22228
rect 15414 22188 15752 22216
rect 15414 22185 15426 22188
rect 15368 22179 15426 22185
rect 15746 22176 15752 22188
rect 15804 22176 15810 22228
rect 20438 22176 20444 22228
rect 20496 22216 20502 22228
rect 22538 22219 22596 22225
rect 22538 22216 22550 22219
rect 20496 22188 22550 22216
rect 20496 22176 20502 22188
rect 22538 22185 22550 22188
rect 22584 22185 22596 22219
rect 22538 22179 22596 22185
rect 26970 22176 26976 22228
rect 27028 22216 27034 22228
rect 27430 22216 27436 22228
rect 27028 22188 27436 22216
rect 27028 22176 27034 22188
rect 27430 22176 27436 22188
rect 27488 22176 27494 22228
rect 28074 22176 28080 22228
rect 28132 22216 28138 22228
rect 28261 22219 28319 22225
rect 28261 22216 28273 22219
rect 28132 22188 28273 22216
rect 28132 22176 28138 22188
rect 28261 22185 28273 22188
rect 28307 22185 28319 22219
rect 28261 22179 28319 22185
rect 28626 22176 28632 22228
rect 28684 22176 28690 22228
rect 30098 22176 30104 22228
rect 30156 22176 30162 22228
rect 32030 22176 32036 22228
rect 32088 22176 32094 22228
rect 32306 22176 32312 22228
rect 32364 22216 32370 22228
rect 32585 22219 32643 22225
rect 32585 22216 32597 22219
rect 32364 22188 32597 22216
rect 32364 22176 32370 22188
rect 32585 22185 32597 22188
rect 32631 22185 32643 22219
rect 32585 22179 32643 22185
rect 33134 22176 33140 22228
rect 33192 22216 33198 22228
rect 33229 22219 33287 22225
rect 33229 22216 33241 22219
rect 33192 22188 33241 22216
rect 33192 22176 33198 22188
rect 33229 22185 33241 22188
rect 33275 22185 33287 22219
rect 33229 22179 33287 22185
rect 34422 22176 34428 22228
rect 34480 22176 34486 22228
rect 34606 22176 34612 22228
rect 34664 22216 34670 22228
rect 34701 22219 34759 22225
rect 34701 22216 34713 22219
rect 34664 22188 34713 22216
rect 34664 22176 34670 22188
rect 34701 22185 34713 22188
rect 34747 22185 34759 22219
rect 34701 22179 34759 22185
rect 36446 22176 36452 22228
rect 36504 22216 36510 22228
rect 36541 22219 36599 22225
rect 36541 22216 36553 22219
rect 36504 22188 36553 22216
rect 36504 22176 36510 22188
rect 36541 22185 36553 22188
rect 36587 22185 36599 22219
rect 36541 22179 36599 22185
rect 37550 22176 37556 22228
rect 37608 22216 37614 22228
rect 37829 22219 37887 22225
rect 37829 22216 37841 22219
rect 37608 22188 37841 22216
rect 37608 22176 37614 22188
rect 37829 22185 37841 22188
rect 37875 22185 37887 22219
rect 37829 22179 37887 22185
rect 8846 22148 8852 22160
rect 6932 22120 8852 22148
rect 6932 22080 6960 22120
rect 8846 22108 8852 22120
rect 8904 22108 8910 22160
rect 20898 22108 20904 22160
rect 20956 22148 20962 22160
rect 21634 22148 21640 22160
rect 20956 22120 21640 22148
rect 20956 22108 20962 22120
rect 21634 22108 21640 22120
rect 21692 22108 21698 22160
rect 4672 22052 5304 22080
rect 5736 22052 6960 22080
rect 8389 22083 8447 22089
rect 4672 22040 4678 22052
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 22012 3111 22015
rect 3786 22012 3792 22024
rect 3099 21984 3792 22012
rect 3099 21981 3111 21984
rect 3053 21975 3111 21981
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 5166 21972 5172 22024
rect 5224 21972 5230 22024
rect 5276 22012 5304 22052
rect 8389 22049 8401 22083
rect 8435 22080 8447 22083
rect 8478 22080 8484 22092
rect 8435 22052 8484 22080
rect 8435 22049 8447 22052
rect 8389 22043 8447 22049
rect 8478 22040 8484 22052
rect 8536 22040 8542 22092
rect 8665 22083 8723 22089
rect 8665 22049 8677 22083
rect 8711 22080 8723 22083
rect 9950 22080 9956 22092
rect 8711 22052 9956 22080
rect 8711 22049 8723 22052
rect 8665 22043 8723 22049
rect 9950 22040 9956 22052
rect 10008 22040 10014 22092
rect 11238 22040 11244 22092
rect 11296 22080 11302 22092
rect 11698 22080 11704 22092
rect 11296 22052 11704 22080
rect 11296 22040 11302 22052
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12161 22083 12219 22089
rect 12161 22080 12173 22083
rect 12115 22052 12173 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 12161 22049 12173 22052
rect 12207 22080 12219 22083
rect 12526 22080 12532 22092
rect 12207 22052 12532 22080
rect 12207 22049 12219 22052
rect 12161 22043 12219 22049
rect 12526 22040 12532 22052
rect 12584 22080 12590 22092
rect 12584 22052 13676 22080
rect 12584 22040 12590 22052
rect 5626 22012 5632 22024
rect 5276 21984 5632 22012
rect 5626 21972 5632 21984
rect 5684 21972 5690 22024
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 22012 8355 22015
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8343 21984 8953 22012
rect 8343 21981 8355 21984
rect 8297 21975 8355 21981
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 9030 21972 9036 22024
rect 9088 22012 9094 22024
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 9088 21984 9505 22012
rect 9088 21972 9094 21984
rect 9493 21981 9505 21984
rect 9539 21981 9551 22015
rect 13648 22012 13676 22052
rect 13722 22040 13728 22092
rect 13780 22080 13786 22092
rect 13909 22083 13967 22089
rect 13909 22080 13921 22083
rect 13780 22052 13921 22080
rect 13780 22040 13786 22052
rect 13909 22049 13921 22052
rect 13955 22049 13967 22083
rect 13909 22043 13967 22049
rect 16114 22040 16120 22092
rect 16172 22080 16178 22092
rect 17129 22083 17187 22089
rect 17129 22080 17141 22083
rect 16172 22052 17141 22080
rect 16172 22040 16178 22052
rect 17129 22049 17141 22052
rect 17175 22049 17187 22083
rect 17129 22043 17187 22049
rect 18969 22083 19027 22089
rect 18969 22049 18981 22083
rect 19015 22080 19027 22083
rect 19242 22080 19248 22092
rect 19015 22052 19248 22080
rect 19015 22049 19027 22052
rect 18969 22043 19027 22049
rect 19242 22040 19248 22052
rect 19300 22080 19306 22092
rect 20806 22080 20812 22092
rect 19300 22052 20812 22080
rect 19300 22040 19306 22052
rect 20806 22040 20812 22052
rect 20864 22080 20870 22092
rect 22281 22083 22339 22089
rect 22281 22080 22293 22083
rect 20864 22052 22293 22080
rect 20864 22040 20870 22052
rect 22281 22049 22293 22052
rect 22327 22080 22339 22083
rect 22922 22080 22928 22092
rect 22327 22052 22928 22080
rect 22327 22049 22339 22052
rect 22281 22043 22339 22049
rect 22922 22040 22928 22052
rect 22980 22040 22986 22092
rect 27065 22083 27123 22089
rect 27065 22049 27077 22083
rect 27111 22080 27123 22083
rect 27890 22080 27896 22092
rect 27111 22052 27896 22080
rect 27111 22049 27123 22052
rect 27065 22043 27123 22049
rect 27890 22040 27896 22052
rect 27948 22040 27954 22092
rect 28644 22080 28672 22176
rect 28276 22052 28672 22080
rect 14182 22012 14188 22024
rect 13648 21984 14188 22012
rect 9493 21975 9551 21981
rect 14182 21972 14188 21984
rect 14240 22012 14246 22024
rect 15105 22015 15163 22021
rect 15105 22012 15117 22015
rect 14240 21984 15117 22012
rect 14240 21972 14246 21984
rect 15105 21981 15117 21984
rect 15151 21981 15163 22015
rect 17402 22012 17408 22024
rect 16514 21984 17408 22012
rect 15105 21975 15163 21981
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 20070 22021 20076 22024
rect 20068 22012 20076 22021
rect 20031 21984 20076 22012
rect 20068 21975 20076 21984
rect 20070 21972 20076 21975
rect 20128 21972 20134 22024
rect 20440 22015 20498 22021
rect 20440 21981 20452 22015
rect 20486 21981 20498 22015
rect 20440 21975 20498 21981
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20622 22012 20628 22024
rect 20579 21984 20628 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 9674 21944 9680 21956
rect 7130 21916 9680 21944
rect 2866 21836 2872 21888
rect 2924 21836 2930 21888
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 3970 21876 3976 21888
rect 3752 21848 3976 21876
rect 3752 21836 3758 21848
rect 3970 21836 3976 21848
rect 4028 21876 4034 21888
rect 7208 21876 7236 21916
rect 9674 21904 9680 21916
rect 9732 21904 9738 21956
rect 11238 21904 11244 21956
rect 11296 21904 11302 21956
rect 11790 21904 11796 21956
rect 11848 21904 11854 21956
rect 12434 21904 12440 21956
rect 12492 21904 12498 21956
rect 13662 21916 14596 21944
rect 4028 21848 7236 21876
rect 10321 21879 10379 21885
rect 4028 21836 4034 21848
rect 10321 21845 10333 21879
rect 10367 21876 10379 21879
rect 11054 21876 11060 21888
rect 10367 21848 11060 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 11698 21836 11704 21888
rect 11756 21876 11762 21888
rect 13740 21876 13768 21916
rect 11756 21848 13768 21876
rect 14568 21876 14596 21916
rect 16666 21904 16672 21956
rect 16724 21944 16730 21956
rect 16724 21916 17526 21944
rect 16724 21904 16730 21916
rect 18690 21904 18696 21956
rect 18748 21904 18754 21956
rect 20165 21947 20223 21953
rect 20165 21913 20177 21947
rect 20211 21913 20223 21947
rect 20165 21907 20223 21913
rect 20257 21947 20315 21953
rect 20257 21913 20269 21947
rect 20303 21913 20315 21947
rect 20456 21944 20484 21975
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 20990 21972 20996 22024
rect 21048 22012 21054 22024
rect 21358 22021 21364 22024
rect 21177 22015 21235 22021
rect 21177 22012 21189 22015
rect 21048 21984 21189 22012
rect 21048 21972 21054 21984
rect 21177 21981 21189 21984
rect 21223 21981 21235 22015
rect 21177 21975 21235 21981
rect 21335 22015 21364 22021
rect 21335 21981 21347 22015
rect 21335 21975 21364 21981
rect 21358 21972 21364 21975
rect 21416 21972 21422 22024
rect 21634 21972 21640 22024
rect 21692 21972 21698 22024
rect 21818 21972 21824 22024
rect 21876 21972 21882 22024
rect 26602 21972 26608 22024
rect 26660 22012 26666 22024
rect 28276 22021 28304 22052
rect 28810 22040 28816 22092
rect 28868 22040 28874 22092
rect 30190 22040 30196 22092
rect 30248 22080 30254 22092
rect 30469 22083 30527 22089
rect 30469 22080 30481 22083
rect 30248 22052 30481 22080
rect 30248 22040 30254 22052
rect 30469 22049 30481 22052
rect 30515 22049 30527 22083
rect 30469 22043 30527 22049
rect 35250 22040 35256 22092
rect 35308 22080 35314 22092
rect 35529 22083 35587 22089
rect 35529 22080 35541 22083
rect 35308 22052 35541 22080
rect 35308 22040 35314 22052
rect 35529 22049 35541 22052
rect 35575 22049 35587 22083
rect 35529 22043 35587 22049
rect 37274 22040 37280 22092
rect 37332 22080 37338 22092
rect 37332 22052 37688 22080
rect 37332 22040 37338 22052
rect 26973 22015 27031 22021
rect 26973 22012 26985 22015
rect 26660 21984 26985 22012
rect 26660 21972 26666 21984
rect 26973 21981 26985 21984
rect 27019 21981 27031 22015
rect 26973 21975 27031 21981
rect 28077 22015 28135 22021
rect 28077 21981 28089 22015
rect 28123 21981 28135 22015
rect 28077 21975 28135 21981
rect 28261 22015 28319 22021
rect 28261 21981 28273 22015
rect 28307 21981 28319 22015
rect 28261 21975 28319 21981
rect 20714 21944 20720 21956
rect 20456 21916 20720 21944
rect 20257 21907 20315 21913
rect 16684 21876 16712 21904
rect 14568 21848 16712 21876
rect 17221 21879 17279 21885
rect 11756 21836 11762 21848
rect 17221 21845 17233 21879
rect 17267 21876 17279 21879
rect 18046 21876 18052 21888
rect 17267 21848 18052 21876
rect 17267 21845 17279 21848
rect 17221 21839 17279 21845
rect 18046 21836 18052 21848
rect 18104 21836 18110 21888
rect 19886 21836 19892 21888
rect 19944 21836 19950 21888
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 20180 21876 20208 21907
rect 20128 21848 20208 21876
rect 20272 21876 20300 21907
rect 20714 21904 20720 21916
rect 20772 21904 20778 21956
rect 21450 21904 21456 21956
rect 21508 21904 21514 21956
rect 21545 21947 21603 21953
rect 21545 21913 21557 21947
rect 21591 21944 21603 21947
rect 22094 21944 22100 21956
rect 21591 21916 22100 21944
rect 21591 21913 21603 21916
rect 21545 21907 21603 21913
rect 22094 21904 22100 21916
rect 22152 21904 22158 21956
rect 24302 21944 24308 21956
rect 23782 21916 24308 21944
rect 20898 21876 20904 21888
rect 20272 21848 20904 21876
rect 20128 21836 20134 21848
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 21818 21836 21824 21888
rect 21876 21876 21882 21888
rect 23860 21876 23888 21916
rect 24302 21904 24308 21916
rect 24360 21904 24366 21956
rect 25866 21904 25872 21956
rect 25924 21944 25930 21956
rect 28092 21944 28120 21975
rect 28442 21972 28448 22024
rect 28500 21972 28506 22024
rect 28626 21972 28632 22024
rect 28684 22012 28690 22024
rect 28828 22012 28856 22040
rect 28684 21984 28856 22012
rect 28684 21972 28690 21984
rect 29638 21972 29644 22024
rect 29696 22012 29702 22024
rect 30285 22015 30343 22021
rect 30285 22012 30297 22015
rect 29696 21984 30297 22012
rect 29696 21972 29702 21984
rect 30285 21981 30297 21984
rect 30331 21981 30343 22015
rect 32493 22015 32551 22021
rect 32493 22012 32505 22015
rect 30285 21975 30343 21981
rect 32232 21984 32505 22012
rect 28810 21944 28816 21956
rect 25924 21916 28816 21944
rect 25924 21904 25930 21916
rect 28810 21904 28816 21916
rect 28868 21904 28874 21956
rect 29454 21904 29460 21956
rect 29512 21944 29518 21956
rect 32232 21953 32260 21984
rect 32493 21981 32505 21984
rect 32539 21981 32551 22015
rect 32493 21975 32551 21981
rect 32674 21972 32680 22024
rect 32732 21972 32738 22024
rect 32858 21972 32864 22024
rect 32916 21972 32922 22024
rect 34333 22015 34391 22021
rect 34333 21981 34345 22015
rect 34379 22012 34391 22015
rect 34422 22012 34428 22024
rect 34379 21984 34428 22012
rect 34379 21981 34391 21984
rect 34333 21975 34391 21981
rect 34422 21972 34428 21984
rect 34480 21972 34486 22024
rect 34517 22015 34575 22021
rect 34517 21981 34529 22015
rect 34563 22012 34575 22015
rect 35069 22015 35127 22021
rect 35069 22012 35081 22015
rect 34563 21984 35081 22012
rect 34563 21981 34575 21984
rect 34517 21975 34575 21981
rect 35069 21981 35081 21984
rect 35115 22012 35127 22015
rect 35161 22015 35219 22021
rect 35161 22012 35173 22015
rect 35115 21984 35173 22012
rect 35115 21981 35127 21984
rect 35069 21975 35127 21981
rect 35161 21981 35173 21984
rect 35207 21981 35219 22015
rect 35161 21975 35219 21981
rect 35342 21972 35348 22024
rect 35400 21972 35406 22024
rect 36909 22015 36967 22021
rect 36909 21981 36921 22015
rect 36955 22012 36967 22015
rect 37090 22012 37096 22024
rect 36955 21984 37096 22012
rect 36955 21981 36967 21984
rect 36909 21975 36967 21981
rect 37090 21972 37096 21984
rect 37148 22012 37154 22024
rect 37185 22015 37243 22021
rect 37185 22012 37197 22015
rect 37148 21984 37197 22012
rect 37148 21972 37154 21984
rect 37185 21981 37197 21984
rect 37231 21981 37243 22015
rect 37185 21975 37243 21981
rect 37366 21972 37372 22024
rect 37424 21972 37430 22024
rect 37660 22021 37688 22052
rect 37645 22015 37703 22021
rect 37645 21981 37657 22015
rect 37691 21981 37703 22015
rect 37645 21975 37703 21981
rect 32217 21947 32275 21953
rect 32217 21944 32229 21947
rect 29512 21916 32229 21944
rect 29512 21904 29518 21916
rect 32217 21913 32229 21916
rect 32263 21913 32275 21947
rect 32217 21907 32275 21913
rect 32401 21947 32459 21953
rect 32401 21913 32413 21947
rect 32447 21944 32459 21947
rect 32692 21944 32720 21972
rect 32447 21916 32720 21944
rect 32447 21913 32459 21916
rect 32401 21907 32459 21913
rect 33042 21904 33048 21956
rect 33100 21904 33106 21956
rect 34440 21944 34468 21972
rect 34885 21947 34943 21953
rect 34885 21944 34897 21947
rect 34440 21916 34897 21944
rect 34885 21913 34897 21916
rect 34931 21913 34943 21947
rect 34885 21907 34943 21913
rect 36725 21947 36783 21953
rect 36725 21913 36737 21947
rect 36771 21944 36783 21947
rect 37384 21944 37412 21972
rect 36771 21916 37412 21944
rect 37461 21947 37519 21953
rect 36771 21913 36783 21916
rect 36725 21907 36783 21913
rect 37461 21913 37473 21947
rect 37507 21944 37519 21947
rect 37550 21944 37556 21956
rect 37507 21916 37556 21944
rect 37507 21913 37519 21916
rect 37461 21907 37519 21913
rect 21876 21848 23888 21876
rect 24029 21879 24087 21885
rect 21876 21836 21882 21848
rect 24029 21845 24041 21879
rect 24075 21876 24087 21879
rect 25774 21876 25780 21888
rect 24075 21848 25780 21876
rect 24075 21845 24087 21848
rect 24029 21839 24087 21845
rect 25774 21836 25780 21848
rect 25832 21836 25838 21888
rect 28350 21836 28356 21888
rect 28408 21876 28414 21888
rect 29472 21876 29500 21904
rect 28408 21848 29500 21876
rect 28408 21836 28414 21848
rect 34698 21836 34704 21888
rect 34756 21876 34762 21888
rect 36740 21876 36768 21907
rect 37550 21904 37556 21916
rect 37608 21904 37614 21956
rect 34756 21848 36768 21876
rect 34756 21836 34762 21848
rect 1104 21786 38824 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 38824 21786
rect 1104 21712 38824 21734
rect 4341 21675 4399 21681
rect 4341 21641 4353 21675
rect 4387 21672 4399 21675
rect 4706 21672 4712 21684
rect 4387 21644 4712 21672
rect 4387 21641 4399 21644
rect 4341 21635 4399 21641
rect 4706 21632 4712 21644
rect 4764 21632 4770 21684
rect 5997 21675 6055 21681
rect 5997 21641 6009 21675
rect 6043 21672 6055 21675
rect 6178 21672 6184 21684
rect 6043 21644 6184 21672
rect 6043 21641 6055 21644
rect 5997 21635 6055 21641
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 8757 21675 8815 21681
rect 8757 21641 8769 21675
rect 8803 21672 8815 21675
rect 8938 21672 8944 21684
rect 8803 21644 8944 21672
rect 8803 21641 8815 21644
rect 8757 21635 8815 21641
rect 8938 21632 8944 21644
rect 8996 21632 9002 21684
rect 11054 21632 11060 21684
rect 11112 21632 11118 21684
rect 11790 21632 11796 21684
rect 11848 21632 11854 21684
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 13173 21675 13231 21681
rect 13173 21672 13185 21675
rect 12492 21644 13185 21672
rect 12492 21632 12498 21644
rect 13173 21641 13185 21644
rect 13219 21641 13231 21675
rect 13173 21635 13231 21641
rect 13354 21632 13360 21684
rect 13412 21672 13418 21684
rect 14090 21672 14096 21684
rect 13412 21644 14096 21672
rect 13412 21632 13418 21644
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 15102 21632 15108 21684
rect 15160 21672 15166 21684
rect 17402 21672 17408 21684
rect 15160 21644 17408 21672
rect 15160 21632 15166 21644
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 17589 21675 17647 21681
rect 17589 21641 17601 21675
rect 17635 21672 17647 21675
rect 18690 21672 18696 21684
rect 17635 21644 18696 21672
rect 17635 21641 17647 21644
rect 17589 21635 17647 21641
rect 18690 21632 18696 21644
rect 18748 21632 18754 21684
rect 21726 21632 21732 21684
rect 21784 21672 21790 21684
rect 21821 21675 21879 21681
rect 21821 21672 21833 21675
rect 21784 21644 21833 21672
rect 21784 21632 21790 21644
rect 21821 21641 21833 21644
rect 21867 21641 21879 21675
rect 21821 21635 21879 21641
rect 26421 21675 26479 21681
rect 26421 21641 26433 21675
rect 26467 21672 26479 21675
rect 26786 21672 26792 21684
rect 26467 21644 26792 21672
rect 26467 21641 26479 21644
rect 26421 21635 26479 21641
rect 26786 21632 26792 21644
rect 26844 21672 26850 21684
rect 28350 21672 28356 21684
rect 26844 21644 28356 21672
rect 26844 21632 26850 21644
rect 28350 21632 28356 21644
rect 28408 21632 28414 21684
rect 28902 21632 28908 21684
rect 28960 21672 28966 21684
rect 29089 21675 29147 21681
rect 29089 21672 29101 21675
rect 28960 21644 29101 21672
rect 28960 21632 28966 21644
rect 29089 21641 29101 21644
rect 29135 21641 29147 21675
rect 29089 21635 29147 21641
rect 33962 21632 33968 21684
rect 34020 21632 34026 21684
rect 35069 21675 35127 21681
rect 35069 21641 35081 21675
rect 35115 21672 35127 21675
rect 35250 21672 35256 21684
rect 35115 21644 35256 21672
rect 35115 21641 35127 21644
rect 35069 21635 35127 21641
rect 35250 21632 35256 21644
rect 35308 21632 35314 21684
rect 35342 21632 35348 21684
rect 35400 21632 35406 21684
rect 3970 21564 3976 21616
rect 4028 21564 4034 21616
rect 4614 21564 4620 21616
rect 4672 21604 4678 21616
rect 5077 21607 5135 21613
rect 5077 21604 5089 21607
rect 4672 21576 5089 21604
rect 4672 21564 4678 21576
rect 5077 21573 5089 21576
rect 5123 21573 5135 21607
rect 5077 21567 5135 21573
rect 3789 21539 3847 21545
rect 3789 21505 3801 21539
rect 3835 21536 3847 21539
rect 4065 21539 4123 21545
rect 4065 21536 4077 21539
rect 3835 21508 4077 21536
rect 3835 21505 3847 21508
rect 3789 21499 3847 21505
rect 4065 21505 4077 21508
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4525 21539 4583 21545
rect 4525 21505 4537 21539
rect 4571 21505 4583 21539
rect 4525 21499 4583 21505
rect 4080 21400 4108 21499
rect 4540 21468 4568 21499
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21536 5043 21539
rect 5350 21536 5356 21548
rect 5031 21508 5356 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 5350 21496 5356 21508
rect 5408 21496 5414 21548
rect 5718 21496 5724 21548
rect 5776 21496 5782 21548
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 6196 21536 6224 21632
rect 9674 21564 9680 21616
rect 9732 21564 9738 21616
rect 9950 21564 9956 21616
rect 10008 21604 10014 21616
rect 10229 21607 10287 21613
rect 10229 21604 10241 21607
rect 10008 21576 10241 21604
rect 10008 21564 10014 21576
rect 10229 21573 10241 21576
rect 10275 21573 10287 21607
rect 11072 21604 11100 21632
rect 12158 21604 12164 21616
rect 11072 21576 12164 21604
rect 10229 21567 10287 21573
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 12253 21607 12311 21613
rect 12253 21573 12265 21607
rect 12299 21604 12311 21607
rect 12986 21604 12992 21616
rect 12299 21576 12992 21604
rect 12299 21573 12311 21576
rect 12253 21567 12311 21573
rect 12986 21564 12992 21576
rect 13044 21604 13050 21616
rect 13541 21607 13599 21613
rect 13541 21604 13553 21607
rect 13044 21576 13553 21604
rect 13044 21564 13050 21576
rect 13541 21573 13553 21576
rect 13587 21573 13599 21607
rect 16666 21604 16672 21616
rect 15686 21576 16672 21604
rect 13541 21567 13599 21573
rect 16666 21564 16672 21576
rect 16724 21564 16730 21616
rect 20714 21564 20720 21616
rect 20772 21604 20778 21616
rect 25958 21604 25964 21616
rect 20772 21576 22508 21604
rect 20772 21564 20778 21576
rect 21744 21548 21772 21576
rect 6365 21539 6423 21545
rect 6365 21536 6377 21539
rect 6196 21508 6377 21536
rect 6365 21505 6377 21508
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 6454 21496 6460 21548
rect 6512 21536 6518 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6512 21508 6561 21536
rect 6512 21496 6518 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21536 11023 21539
rect 11606 21536 11612 21548
rect 11011 21508 11612 21536
rect 11011 21505 11023 21508
rect 10965 21499 11023 21505
rect 11606 21496 11612 21508
rect 11664 21496 11670 21548
rect 12621 21539 12679 21545
rect 12621 21505 12633 21539
rect 12667 21505 12679 21539
rect 12621 21499 12679 21505
rect 5534 21468 5540 21480
rect 4540 21440 5540 21468
rect 5534 21428 5540 21440
rect 5592 21428 5598 21480
rect 8570 21428 8576 21480
rect 8628 21428 8634 21480
rect 10502 21428 10508 21480
rect 10560 21428 10566 21480
rect 10594 21428 10600 21480
rect 10652 21468 10658 21480
rect 11149 21471 11207 21477
rect 11149 21468 11161 21471
rect 10652 21440 11161 21468
rect 10652 21428 10658 21440
rect 11149 21437 11161 21440
rect 11195 21437 11207 21471
rect 11149 21431 11207 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21437 12495 21471
rect 12636 21468 12664 21499
rect 12710 21496 12716 21548
rect 12768 21536 12774 21548
rect 12805 21539 12863 21545
rect 12805 21536 12817 21539
rect 12768 21508 12817 21536
rect 12768 21496 12774 21508
rect 12805 21505 12817 21508
rect 12851 21505 12863 21539
rect 12805 21499 12863 21505
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21536 12955 21539
rect 13446 21536 13452 21548
rect 12943 21508 13452 21536
rect 12943 21505 12955 21508
rect 12897 21499 12955 21505
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 13630 21496 13636 21548
rect 13688 21536 13694 21548
rect 13688 21508 14136 21536
rect 13688 21496 13694 21508
rect 13538 21468 13544 21480
rect 12636 21440 13544 21468
rect 12437 21431 12495 21437
rect 5442 21400 5448 21412
rect 4080 21372 5448 21400
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 5994 21360 6000 21412
rect 6052 21400 6058 21412
rect 6365 21403 6423 21409
rect 6365 21400 6377 21403
rect 6052 21372 6377 21400
rect 6052 21360 6058 21372
rect 6365 21369 6377 21372
rect 6411 21369 6423 21403
rect 12452 21400 12480 21431
rect 13538 21428 13544 21440
rect 13596 21428 13602 21480
rect 13725 21471 13783 21477
rect 13725 21437 13737 21471
rect 13771 21437 13783 21471
rect 14108 21468 14136 21508
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 16684 21508 17233 21536
rect 14108 21440 14320 21468
rect 13725 21431 13783 21437
rect 13740 21400 13768 21431
rect 14182 21400 14188 21412
rect 12452 21372 14188 21400
rect 6365 21363 6423 21369
rect 14182 21360 14188 21372
rect 14240 21360 14246 21412
rect 4154 21292 4160 21344
rect 4212 21332 4218 21344
rect 4798 21332 4804 21344
rect 4212 21304 4804 21332
rect 4212 21292 4218 21304
rect 4798 21292 4804 21304
rect 4856 21292 4862 21344
rect 7926 21292 7932 21344
rect 7984 21332 7990 21344
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 7984 21304 8033 21332
rect 7984 21292 7990 21304
rect 8021 21301 8033 21304
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 10597 21335 10655 21341
rect 10597 21301 10609 21335
rect 10643 21332 10655 21335
rect 10686 21332 10692 21344
rect 10643 21304 10692 21332
rect 10643 21301 10655 21304
rect 10597 21295 10655 21301
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 12805 21335 12863 21341
rect 12805 21301 12817 21335
rect 12851 21332 12863 21335
rect 12986 21332 12992 21344
rect 12851 21304 12992 21332
rect 12851 21301 12863 21304
rect 12805 21295 12863 21301
rect 12986 21292 12992 21304
rect 13044 21292 13050 21344
rect 13081 21335 13139 21341
rect 13081 21301 13093 21335
rect 13127 21332 13139 21335
rect 13354 21332 13360 21344
rect 13127 21304 13360 21332
rect 13127 21301 13139 21304
rect 13081 21295 13139 21301
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 14292 21332 14320 21440
rect 14458 21428 14464 21480
rect 14516 21428 14522 21480
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 16684 21468 16712 21508
rect 17221 21505 17233 21508
rect 17267 21536 17279 21539
rect 17681 21539 17739 21545
rect 17681 21536 17693 21539
rect 17267 21508 17693 21536
rect 17267 21505 17279 21508
rect 17221 21499 17279 21505
rect 17681 21505 17693 21508
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21536 20683 21539
rect 20898 21536 20904 21548
rect 20671 21508 20904 21536
rect 20671 21505 20683 21508
rect 20625 21499 20683 21505
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21726 21496 21732 21548
rect 21784 21496 21790 21548
rect 21910 21496 21916 21548
rect 21968 21536 21974 21548
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 21968 21508 22201 21536
rect 21968 21496 21974 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22281 21539 22339 21545
rect 22281 21505 22293 21539
rect 22327 21536 22339 21539
rect 22370 21536 22376 21548
rect 22327 21508 22376 21536
rect 22327 21505 22339 21508
rect 22281 21499 22339 21505
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 22480 21545 22508 21576
rect 22756 21576 25964 21604
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 15252 21440 16712 21468
rect 15252 21428 15258 21440
rect 17034 21428 17040 21480
rect 17092 21428 17098 21480
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21468 17187 21471
rect 17954 21468 17960 21480
rect 17175 21440 17960 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 17954 21428 17960 21440
rect 18012 21428 18018 21480
rect 18138 21428 18144 21480
rect 18196 21468 18202 21480
rect 18233 21471 18291 21477
rect 18233 21468 18245 21471
rect 18196 21440 18245 21468
rect 18196 21428 18202 21440
rect 18233 21437 18245 21440
rect 18279 21437 18291 21471
rect 18233 21431 18291 21437
rect 21634 21428 21640 21480
rect 21692 21468 21698 21480
rect 22005 21471 22063 21477
rect 22005 21468 22017 21471
rect 21692 21440 22017 21468
rect 21692 21428 21698 21440
rect 22005 21437 22017 21440
rect 22051 21437 22063 21471
rect 22005 21431 22063 21437
rect 22094 21428 22100 21480
rect 22152 21468 22158 21480
rect 22554 21468 22560 21480
rect 22152 21440 22560 21468
rect 22152 21428 22158 21440
rect 22554 21428 22560 21440
rect 22612 21428 22618 21480
rect 21818 21400 21824 21412
rect 20364 21372 21824 21400
rect 20364 21344 20392 21372
rect 21818 21360 21824 21372
rect 21876 21360 21882 21412
rect 22756 21400 22784 21576
rect 25958 21564 25964 21576
rect 26016 21604 26022 21616
rect 29914 21604 29920 21616
rect 26016 21576 29920 21604
rect 26016 21564 26022 21576
rect 29914 21564 29920 21576
rect 29972 21564 29978 21616
rect 34330 21604 34336 21616
rect 34072 21576 34336 21604
rect 25041 21539 25099 21545
rect 25041 21505 25053 21539
rect 25087 21536 25099 21539
rect 25087 21508 25728 21536
rect 25087 21505 25099 21508
rect 25041 21499 25099 21505
rect 25130 21428 25136 21480
rect 25188 21428 25194 21480
rect 25317 21471 25375 21477
rect 25317 21437 25329 21471
rect 25363 21468 25375 21471
rect 25700 21468 25728 21508
rect 25774 21496 25780 21548
rect 25832 21496 25838 21548
rect 25866 21496 25872 21548
rect 25924 21496 25930 21548
rect 26329 21539 26387 21545
rect 26329 21505 26341 21539
rect 26375 21536 26387 21539
rect 26970 21536 26976 21548
rect 26375 21508 26976 21536
rect 26375 21505 26387 21508
rect 26329 21499 26387 21505
rect 25363 21440 25636 21468
rect 25700 21440 26096 21468
rect 25363 21437 25375 21440
rect 25317 21431 25375 21437
rect 22066 21372 22784 21400
rect 22066 21344 22094 21372
rect 15562 21332 15568 21344
rect 14292 21304 15568 21332
rect 15562 21292 15568 21304
rect 15620 21332 15626 21344
rect 15933 21335 15991 21341
rect 15933 21332 15945 21335
rect 15620 21304 15945 21332
rect 15620 21292 15626 21304
rect 15933 21301 15945 21304
rect 15979 21301 15991 21335
rect 15933 21295 15991 21301
rect 20346 21292 20352 21344
rect 20404 21292 20410 21344
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 21542 21332 21548 21344
rect 20956 21304 21548 21332
rect 20956 21292 20962 21304
rect 21542 21292 21548 21304
rect 21600 21332 21606 21344
rect 22002 21332 22008 21344
rect 21600 21304 22008 21332
rect 21600 21292 21606 21304
rect 22002 21292 22008 21304
rect 22060 21304 22094 21344
rect 22060 21292 22066 21304
rect 22554 21292 22560 21344
rect 22612 21292 22618 21344
rect 23842 21292 23848 21344
rect 23900 21332 23906 21344
rect 25608 21341 25636 21440
rect 26068 21409 26096 21440
rect 26053 21403 26111 21409
rect 26053 21369 26065 21403
rect 26099 21400 26111 21403
rect 26234 21400 26240 21412
rect 26099 21372 26240 21400
rect 26099 21369 26111 21372
rect 26053 21363 26111 21369
rect 26234 21360 26240 21372
rect 26292 21400 26298 21412
rect 26344 21400 26372 21499
rect 26970 21496 26976 21508
rect 27028 21496 27034 21548
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21536 27215 21539
rect 27798 21536 27804 21548
rect 27203 21508 27804 21536
rect 27203 21505 27215 21508
rect 27157 21499 27215 21505
rect 27798 21496 27804 21508
rect 27856 21536 27862 21548
rect 28626 21536 28632 21548
rect 27856 21508 28632 21536
rect 27856 21496 27862 21508
rect 28626 21496 28632 21508
rect 28684 21536 28690 21548
rect 28905 21539 28963 21545
rect 28905 21536 28917 21539
rect 28684 21508 28917 21536
rect 28684 21496 28690 21508
rect 28905 21505 28917 21508
rect 28951 21505 28963 21539
rect 28905 21499 28963 21505
rect 29270 21496 29276 21548
rect 29328 21496 29334 21548
rect 29454 21496 29460 21548
rect 29512 21496 29518 21548
rect 29638 21496 29644 21548
rect 29696 21536 29702 21548
rect 30009 21539 30067 21545
rect 30009 21536 30021 21539
rect 29696 21508 30021 21536
rect 29696 21496 29702 21508
rect 30009 21505 30021 21508
rect 30055 21505 30067 21539
rect 30009 21499 30067 21505
rect 30190 21496 30196 21548
rect 30248 21496 30254 21548
rect 32306 21496 32312 21548
rect 32364 21496 32370 21548
rect 33870 21496 33876 21548
rect 33928 21496 33934 21548
rect 34072 21545 34100 21576
rect 34330 21564 34336 21576
rect 34388 21604 34394 21616
rect 34701 21607 34759 21613
rect 34701 21604 34713 21607
rect 34388 21576 34713 21604
rect 34388 21564 34394 21576
rect 34701 21573 34713 21576
rect 34747 21604 34759 21607
rect 34747 21576 35204 21604
rect 34747 21573 34759 21576
rect 34701 21567 34759 21573
rect 35176 21545 35204 21576
rect 34057 21539 34115 21545
rect 34057 21505 34069 21539
rect 34103 21505 34115 21539
rect 34057 21499 34115 21505
rect 34885 21539 34943 21545
rect 34885 21505 34897 21539
rect 34931 21505 34943 21539
rect 34885 21499 34943 21505
rect 35161 21539 35219 21545
rect 35161 21505 35173 21539
rect 35207 21505 35219 21539
rect 35161 21499 35219 21505
rect 35345 21539 35403 21545
rect 35345 21505 35357 21539
rect 35391 21536 35403 21539
rect 36722 21536 36728 21548
rect 35391 21508 36728 21536
rect 35391 21505 35403 21508
rect 35345 21499 35403 21505
rect 28442 21428 28448 21480
rect 28500 21468 28506 21480
rect 28721 21471 28779 21477
rect 28721 21468 28733 21471
rect 28500 21440 28733 21468
rect 28500 21428 28506 21440
rect 28721 21437 28733 21440
rect 28767 21468 28779 21471
rect 29656 21468 29684 21496
rect 28767 21440 29684 21468
rect 28767 21437 28779 21440
rect 28721 21431 28779 21437
rect 26292 21372 26372 21400
rect 26292 21360 26298 21372
rect 28994 21360 29000 21412
rect 29052 21400 29058 21412
rect 30208 21400 30236 21496
rect 31754 21428 31760 21480
rect 31812 21468 31818 21480
rect 32217 21471 32275 21477
rect 32217 21468 32229 21471
rect 31812 21440 32229 21468
rect 31812 21428 31818 21440
rect 32217 21437 32229 21440
rect 32263 21437 32275 21471
rect 32217 21431 32275 21437
rect 32674 21428 32680 21480
rect 32732 21428 32738 21480
rect 34900 21468 34928 21499
rect 35360 21468 35388 21499
rect 36722 21496 36728 21508
rect 36780 21496 36786 21548
rect 34900 21440 35388 21468
rect 29052 21372 30236 21400
rect 29052 21360 29058 21372
rect 24673 21335 24731 21341
rect 24673 21332 24685 21335
rect 23900 21304 24685 21332
rect 23900 21292 23906 21304
rect 24673 21301 24685 21304
rect 24719 21301 24731 21335
rect 24673 21295 24731 21301
rect 25593 21335 25651 21341
rect 25593 21301 25605 21335
rect 25639 21332 25651 21335
rect 26694 21332 26700 21344
rect 25639 21304 26700 21332
rect 25639 21301 25651 21304
rect 25593 21295 25651 21301
rect 26694 21292 26700 21304
rect 26752 21292 26758 21344
rect 27065 21335 27123 21341
rect 27065 21301 27077 21335
rect 27111 21332 27123 21335
rect 27246 21332 27252 21344
rect 27111 21304 27252 21332
rect 27111 21301 27123 21304
rect 27065 21295 27123 21301
rect 27246 21292 27252 21304
rect 27304 21292 27310 21344
rect 29178 21292 29184 21344
rect 29236 21332 29242 21344
rect 29457 21335 29515 21341
rect 29457 21332 29469 21335
rect 29236 21304 29469 21332
rect 29236 21292 29242 21304
rect 29457 21301 29469 21304
rect 29503 21301 29515 21335
rect 29457 21295 29515 21301
rect 30374 21292 30380 21344
rect 30432 21292 30438 21344
rect 36354 21292 36360 21344
rect 36412 21332 36418 21344
rect 38194 21332 38200 21344
rect 36412 21304 38200 21332
rect 36412 21292 36418 21304
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 7561 21131 7619 21137
rect 7561 21097 7573 21131
rect 7607 21128 7619 21131
rect 9398 21128 9404 21140
rect 7607 21100 9404 21128
rect 7607 21097 7619 21100
rect 7561 21091 7619 21097
rect 9398 21088 9404 21100
rect 9456 21088 9462 21140
rect 13446 21088 13452 21140
rect 13504 21088 13510 21140
rect 13538 21088 13544 21140
rect 13596 21128 13602 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 13596 21100 13645 21128
rect 13596 21088 13602 21100
rect 13633 21097 13645 21100
rect 13679 21128 13691 21131
rect 13722 21128 13728 21140
rect 13679 21100 13728 21128
rect 13679 21097 13691 21100
rect 13633 21091 13691 21097
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 14182 21088 14188 21140
rect 14240 21128 14246 21140
rect 14240 21100 14412 21128
rect 14240 21088 14246 21100
rect 7929 21063 7987 21069
rect 7929 21029 7941 21063
rect 7975 21060 7987 21063
rect 7975 21032 8616 21060
rect 7975 21029 7987 21032
rect 7929 21023 7987 21029
rect 5626 20952 5632 21004
rect 5684 20952 5690 21004
rect 8478 20992 8484 21004
rect 7392 20964 8484 20992
rect 2866 20884 2872 20936
rect 2924 20884 2930 20936
rect 3053 20927 3111 20933
rect 3053 20893 3065 20927
rect 3099 20924 3111 20927
rect 3878 20924 3884 20936
rect 3099 20896 3884 20924
rect 3099 20893 3111 20896
rect 3053 20887 3111 20893
rect 3878 20884 3884 20896
rect 3936 20884 3942 20936
rect 7392 20933 7420 20964
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 8588 21001 8616 21032
rect 12820 21032 13768 21060
rect 8573 20995 8631 21001
rect 8573 20961 8585 20995
rect 8619 20961 8631 20995
rect 8573 20955 8631 20961
rect 10686 20952 10692 21004
rect 10744 20952 10750 21004
rect 7377 20927 7435 20933
rect 7377 20893 7389 20927
rect 7423 20893 7435 20927
rect 7377 20887 7435 20893
rect 7561 20927 7619 20933
rect 7561 20893 7573 20927
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 3513 20859 3571 20865
rect 3513 20825 3525 20859
rect 3559 20856 3571 20859
rect 3694 20856 3700 20868
rect 3559 20828 3700 20856
rect 3559 20825 3571 20828
rect 3513 20819 3571 20825
rect 3694 20816 3700 20828
rect 3752 20816 3758 20868
rect 4798 20816 4804 20868
rect 4856 20816 4862 20868
rect 5350 20816 5356 20868
rect 5408 20816 5414 20868
rect 7576 20856 7604 20887
rect 7650 20884 7656 20936
rect 7708 20884 7714 20936
rect 7926 20884 7932 20936
rect 7984 20884 7990 20936
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 10410 20924 10416 20936
rect 9732 20896 10416 20924
rect 9732 20884 9738 20896
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 12158 20884 12164 20936
rect 12216 20924 12222 20936
rect 12713 20927 12771 20933
rect 12713 20924 12725 20927
rect 12216 20896 12725 20924
rect 12216 20884 12222 20896
rect 12713 20893 12725 20896
rect 12759 20924 12771 20927
rect 12820 20924 12848 21032
rect 13078 20952 13084 21004
rect 13136 20992 13142 21004
rect 13740 21001 13768 21032
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 14277 21063 14335 21069
rect 14277 21060 14289 21063
rect 13872 21032 14289 21060
rect 13872 21020 13878 21032
rect 14277 21029 14289 21032
rect 14323 21029 14335 21063
rect 14384 21060 14412 21100
rect 14458 21088 14464 21140
rect 14516 21128 14522 21140
rect 14737 21131 14795 21137
rect 14737 21128 14749 21131
rect 14516 21100 14749 21128
rect 14516 21088 14522 21100
rect 14737 21097 14749 21100
rect 14783 21097 14795 21131
rect 15930 21128 15936 21140
rect 14737 21091 14795 21097
rect 15304 21100 15936 21128
rect 15304 21060 15332 21100
rect 15930 21088 15936 21100
rect 15988 21128 15994 21140
rect 17126 21128 17132 21140
rect 15988 21100 17132 21128
rect 15988 21088 15994 21100
rect 14384 21032 15332 21060
rect 14277 21023 14335 21029
rect 13725 20995 13783 21001
rect 13136 20964 13584 20992
rect 13136 20952 13142 20964
rect 12759 20896 12848 20924
rect 12897 20927 12955 20933
rect 12759 20893 12771 20896
rect 12713 20887 12771 20893
rect 12897 20893 12909 20927
rect 12943 20924 12955 20927
rect 12986 20924 12992 20936
rect 12943 20896 12992 20924
rect 12943 20893 12955 20896
rect 12897 20887 12955 20893
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20924 13231 20927
rect 13354 20924 13360 20936
rect 13219 20896 13360 20924
rect 13219 20893 13231 20896
rect 13173 20887 13231 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13556 20924 13584 20964
rect 13725 20961 13737 20995
rect 13771 20992 13783 20995
rect 14369 20995 14427 21001
rect 14369 20992 14381 20995
rect 13771 20964 14381 20992
rect 13771 20961 13783 20964
rect 13725 20955 13783 20961
rect 14369 20961 14381 20964
rect 14415 20961 14427 20995
rect 14369 20955 14427 20961
rect 15194 20952 15200 21004
rect 15252 20952 15258 21004
rect 15304 21001 15332 21032
rect 16209 21063 16267 21069
rect 16209 21029 16221 21063
rect 16255 21060 16267 21063
rect 16666 21060 16672 21072
rect 16255 21032 16672 21060
rect 16255 21029 16267 21032
rect 16209 21023 16267 21029
rect 16666 21020 16672 21032
rect 16724 21020 16730 21072
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20961 15347 20995
rect 16850 20992 16856 21004
rect 15289 20955 15347 20961
rect 15488 20964 15792 20992
rect 14185 20927 14243 20933
rect 14185 20924 14197 20927
rect 13556 20896 14197 20924
rect 14185 20893 14197 20896
rect 14231 20893 14243 20927
rect 14185 20887 14243 20893
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20893 14519 20927
rect 15488 20924 15516 20964
rect 14461 20887 14519 20893
rect 14568 20896 15516 20924
rect 8021 20859 8079 20865
rect 8021 20856 8033 20859
rect 7576 20828 8033 20856
rect 8021 20825 8033 20828
rect 8067 20825 8079 20859
rect 8021 20819 8079 20825
rect 11238 20816 11244 20868
rect 11296 20816 11302 20868
rect 13449 20859 13507 20865
rect 13449 20856 13461 20859
rect 12728 20828 13461 20856
rect 12728 20800 12756 20828
rect 13449 20825 13461 20828
rect 13495 20856 13507 20859
rect 13630 20856 13636 20868
rect 13495 20828 13636 20856
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 13630 20816 13636 20828
rect 13688 20816 13694 20868
rect 13722 20816 13728 20868
rect 13780 20856 13786 20868
rect 13817 20859 13875 20865
rect 13817 20856 13829 20859
rect 13780 20828 13829 20856
rect 13780 20816 13786 20828
rect 13817 20825 13829 20828
rect 13863 20856 13875 20859
rect 14476 20856 14504 20887
rect 13863 20828 14504 20856
rect 13863 20825 13875 20828
rect 13817 20819 13875 20825
rect 2774 20748 2780 20800
rect 2832 20788 2838 20800
rect 2961 20791 3019 20797
rect 2961 20788 2973 20791
rect 2832 20760 2973 20788
rect 2832 20748 2838 20760
rect 2961 20757 2973 20760
rect 3007 20757 3019 20791
rect 2961 20751 3019 20757
rect 3418 20748 3424 20800
rect 3476 20748 3482 20800
rect 3881 20791 3939 20797
rect 3881 20757 3893 20791
rect 3927 20788 3939 20791
rect 4706 20788 4712 20800
rect 3927 20760 4712 20788
rect 3927 20757 3939 20760
rect 3881 20751 3939 20757
rect 4706 20748 4712 20760
rect 4764 20748 4770 20800
rect 7742 20748 7748 20800
rect 7800 20748 7806 20800
rect 12158 20748 12164 20800
rect 12216 20748 12222 20800
rect 12710 20748 12716 20800
rect 12768 20748 12774 20800
rect 13357 20791 13415 20797
rect 13357 20757 13369 20791
rect 13403 20788 13415 20791
rect 14568 20788 14596 20896
rect 15562 20884 15568 20936
rect 15620 20884 15626 20936
rect 15764 20933 15792 20964
rect 16040 20964 16856 20992
rect 16040 20933 16068 20964
rect 16850 20952 16856 20964
rect 16908 20952 16914 21004
rect 16972 21001 17000 21100
rect 17126 21088 17132 21100
rect 17184 21088 17190 21140
rect 17954 21088 17960 21140
rect 18012 21088 18018 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 20990 21128 20996 21140
rect 19392 21100 20996 21128
rect 19392 21088 19398 21100
rect 20990 21088 20996 21100
rect 21048 21088 21054 21140
rect 21726 21088 21732 21140
rect 21784 21088 21790 21140
rect 22370 21088 22376 21140
rect 22428 21088 22434 21140
rect 25130 21088 25136 21140
rect 25188 21128 25194 21140
rect 26329 21131 26387 21137
rect 26329 21128 26341 21131
rect 25188 21100 26341 21128
rect 25188 21088 25194 21100
rect 26329 21097 26341 21100
rect 26375 21097 26387 21131
rect 26329 21091 26387 21097
rect 26878 21088 26884 21140
rect 26936 21128 26942 21140
rect 28166 21128 28172 21140
rect 26936 21100 28172 21128
rect 26936 21088 26942 21100
rect 28166 21088 28172 21100
rect 28224 21128 28230 21140
rect 28261 21131 28319 21137
rect 28261 21128 28273 21131
rect 28224 21100 28273 21128
rect 28224 21088 28230 21100
rect 28261 21097 28273 21100
rect 28307 21097 28319 21131
rect 28261 21091 28319 21097
rect 29362 21088 29368 21140
rect 29420 21128 29426 21140
rect 29641 21131 29699 21137
rect 29641 21128 29653 21131
rect 29420 21100 29653 21128
rect 29420 21088 29426 21100
rect 29641 21097 29653 21100
rect 29687 21097 29699 21131
rect 29641 21091 29699 21097
rect 31754 21088 31760 21140
rect 31812 21088 31818 21140
rect 32585 21131 32643 21137
rect 32585 21097 32597 21131
rect 32631 21128 32643 21131
rect 33042 21128 33048 21140
rect 32631 21100 33048 21128
rect 32631 21097 32643 21100
rect 32585 21091 32643 21097
rect 33042 21088 33048 21100
rect 33100 21088 33106 21140
rect 33781 21131 33839 21137
rect 33781 21097 33793 21131
rect 33827 21128 33839 21131
rect 33870 21128 33876 21140
rect 33827 21100 33876 21128
rect 33827 21097 33839 21100
rect 33781 21091 33839 21097
rect 33870 21088 33876 21100
rect 33928 21088 33934 21140
rect 34330 21088 34336 21140
rect 34388 21088 34394 21140
rect 35897 21131 35955 21137
rect 35897 21097 35909 21131
rect 35943 21128 35955 21131
rect 35986 21128 35992 21140
rect 35943 21100 35992 21128
rect 35943 21097 35955 21100
rect 35897 21091 35955 21097
rect 35986 21088 35992 21100
rect 36044 21088 36050 21140
rect 36722 21088 36728 21140
rect 36780 21088 36786 21140
rect 37550 21088 37556 21140
rect 37608 21088 37614 21140
rect 17034 21020 17040 21072
rect 17092 21060 17098 21072
rect 18509 21063 18567 21069
rect 18509 21060 18521 21063
rect 17092 21032 18521 21060
rect 17092 21020 17098 21032
rect 18509 21029 18521 21032
rect 18555 21029 18567 21063
rect 18509 21023 18567 21029
rect 21174 21020 21180 21072
rect 21232 21060 21238 21072
rect 21545 21063 21603 21069
rect 21545 21060 21557 21063
rect 21232 21032 21557 21060
rect 21232 21020 21238 21032
rect 21545 21029 21557 21032
rect 21591 21060 21603 21063
rect 22646 21060 22652 21072
rect 21591 21032 22652 21060
rect 21591 21029 21603 21032
rect 21545 21023 21603 21029
rect 22646 21020 22652 21032
rect 22704 21020 22710 21072
rect 28074 21060 28080 21072
rect 26804 21032 28080 21060
rect 16945 20995 17003 21001
rect 16945 20961 16957 20995
rect 16991 20961 17003 20995
rect 16945 20955 17003 20961
rect 17862 20952 17868 21004
rect 17920 20992 17926 21004
rect 18693 20995 18751 21001
rect 17920 20964 18460 20992
rect 17920 20952 17926 20964
rect 18432 20933 18460 20964
rect 18693 20961 18705 20995
rect 18739 20992 18751 20995
rect 18782 20992 18788 21004
rect 18739 20964 18788 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 19242 20952 19248 21004
rect 19300 20952 19306 21004
rect 21266 20952 21272 21004
rect 21324 20992 21330 21004
rect 21450 20992 21456 21004
rect 21324 20964 21456 20992
rect 21324 20952 21330 20964
rect 21450 20952 21456 20964
rect 21508 20992 21514 21004
rect 21508 20964 22140 20992
rect 21508 20952 21514 20964
rect 15749 20927 15807 20933
rect 15749 20893 15761 20927
rect 15795 20893 15807 20927
rect 15749 20887 15807 20893
rect 16025 20927 16083 20933
rect 16025 20893 16037 20927
rect 16071 20893 16083 20927
rect 17957 20927 18015 20933
rect 16025 20887 16083 20893
rect 16316 20896 17724 20924
rect 14645 20859 14703 20865
rect 14645 20825 14657 20859
rect 14691 20856 14703 20859
rect 16316 20856 16344 20896
rect 14691 20828 16344 20856
rect 16761 20859 16819 20865
rect 14691 20825 14703 20828
rect 14645 20819 14703 20825
rect 16761 20825 16773 20859
rect 16807 20856 16819 20859
rect 17221 20859 17279 20865
rect 17221 20856 17233 20859
rect 16807 20828 17233 20856
rect 16807 20825 16819 20828
rect 16761 20819 16819 20825
rect 17221 20825 17233 20828
rect 17267 20825 17279 20859
rect 17696 20856 17724 20896
rect 17957 20893 17969 20927
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 17972 20856 18000 20887
rect 17696 20828 18000 20856
rect 17221 20819 17279 20825
rect 13403 20760 14596 20788
rect 15105 20791 15163 20797
rect 13403 20757 13415 20760
rect 13357 20751 13415 20757
rect 15105 20757 15117 20791
rect 15151 20788 15163 20791
rect 15562 20788 15568 20800
rect 15151 20760 15568 20788
rect 15151 20757 15163 20760
rect 15105 20751 15163 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 16390 20748 16396 20800
rect 16448 20748 16454 20800
rect 16850 20748 16856 20800
rect 16908 20748 16914 20800
rect 16942 20748 16948 20800
rect 17000 20788 17006 20800
rect 18064 20788 18092 20887
rect 21818 20884 21824 20936
rect 21876 20884 21882 20936
rect 22112 20933 22140 20964
rect 24394 20952 24400 21004
rect 24452 20952 24458 21004
rect 24765 20995 24823 21001
rect 24765 20961 24777 20995
rect 24811 20992 24823 20995
rect 26804 20992 26832 21032
rect 28074 21020 28080 21032
rect 28132 21020 28138 21072
rect 28994 21020 29000 21072
rect 29052 21060 29058 21072
rect 29052 21032 29224 21060
rect 29052 21020 29058 21032
rect 24811 20964 26832 20992
rect 26881 20995 26939 21001
rect 24811 20961 24823 20964
rect 24765 20955 24823 20961
rect 26881 20961 26893 20995
rect 26927 20992 26939 20995
rect 27062 20992 27068 21004
rect 26927 20964 27068 20992
rect 26927 20961 26939 20964
rect 26881 20955 26939 20961
rect 27062 20952 27068 20964
rect 27120 20952 27126 21004
rect 29089 20995 29147 21001
rect 29089 20992 29101 20995
rect 28644 20964 29101 20992
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20924 22155 20927
rect 22373 20927 22431 20933
rect 22373 20924 22385 20927
rect 22143 20896 22385 20924
rect 22143 20893 22155 20896
rect 22097 20887 22155 20893
rect 22373 20893 22385 20896
rect 22419 20893 22431 20927
rect 22373 20887 22431 20893
rect 22462 20884 22468 20936
rect 22520 20924 22526 20936
rect 22741 20927 22799 20933
rect 22741 20924 22753 20927
rect 22520 20896 22753 20924
rect 22520 20884 22526 20896
rect 22741 20893 22753 20896
rect 22787 20924 22799 20927
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22787 20896 22845 20924
rect 22787 20893 22799 20896
rect 22741 20887 22799 20893
rect 22833 20893 22845 20896
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 23014 20884 23020 20936
rect 23072 20884 23078 20936
rect 23290 20884 23296 20936
rect 23348 20884 23354 20936
rect 26786 20884 26792 20936
rect 26844 20884 26850 20936
rect 26970 20884 26976 20936
rect 27028 20924 27034 20936
rect 27157 20927 27215 20933
rect 27157 20924 27169 20927
rect 27028 20896 27169 20924
rect 27028 20884 27034 20896
rect 27157 20893 27169 20896
rect 27203 20893 27215 20927
rect 27157 20887 27215 20893
rect 27341 20927 27399 20933
rect 27341 20893 27353 20927
rect 27387 20924 27399 20927
rect 27798 20924 27804 20936
rect 27387 20896 27804 20924
rect 27387 20893 27399 20896
rect 27341 20887 27399 20893
rect 18230 20816 18236 20868
rect 18288 20856 18294 20868
rect 18288 20828 19104 20856
rect 18288 20816 18294 20828
rect 18138 20788 18144 20800
rect 17000 20760 18144 20788
rect 17000 20748 17006 20760
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 18325 20791 18383 20797
rect 18325 20757 18337 20791
rect 18371 20788 18383 20791
rect 18506 20788 18512 20800
rect 18371 20760 18512 20788
rect 18371 20757 18383 20760
rect 18325 20751 18383 20757
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 18690 20748 18696 20800
rect 18748 20748 18754 20800
rect 19076 20797 19104 20828
rect 19518 20816 19524 20868
rect 19576 20816 19582 20868
rect 19628 20828 20010 20856
rect 19061 20791 19119 20797
rect 19061 20757 19073 20791
rect 19107 20788 19119 20791
rect 19628 20788 19656 20828
rect 20990 20816 20996 20868
rect 21048 20856 21054 20868
rect 23201 20859 23259 20865
rect 23201 20856 23213 20859
rect 21048 20828 23213 20856
rect 21048 20816 21054 20828
rect 23201 20825 23213 20828
rect 23247 20856 23259 20859
rect 23474 20856 23480 20868
rect 23247 20828 23480 20856
rect 23247 20825 23259 20828
rect 23201 20819 23259 20825
rect 23474 20816 23480 20828
rect 23532 20816 23538 20868
rect 25498 20816 25504 20868
rect 25556 20816 25562 20868
rect 26237 20859 26295 20865
rect 26237 20825 26249 20859
rect 26283 20856 26295 20859
rect 27356 20856 27384 20887
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 28077 20927 28135 20933
rect 28077 20893 28089 20927
rect 28123 20924 28135 20927
rect 28169 20927 28227 20933
rect 28169 20924 28181 20927
rect 28123 20896 28181 20924
rect 28123 20893 28135 20896
rect 28077 20887 28135 20893
rect 28169 20893 28181 20896
rect 28215 20893 28227 20927
rect 28169 20887 28227 20893
rect 28350 20884 28356 20936
rect 28408 20884 28414 20936
rect 28644 20933 28672 20964
rect 29089 20961 29101 20964
rect 29135 20961 29147 20995
rect 29196 20992 29224 21032
rect 29270 21020 29276 21072
rect 29328 21060 29334 21072
rect 36357 21063 36415 21069
rect 29328 21032 33732 21060
rect 29328 21020 29334 21032
rect 29196 20964 30512 20992
rect 29089 20955 29147 20961
rect 29472 20936 29500 20964
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28810 20884 28816 20936
rect 28868 20884 28874 20936
rect 28902 20884 28908 20936
rect 28960 20884 28966 20936
rect 28994 20884 29000 20936
rect 29052 20884 29058 20936
rect 29178 20884 29184 20936
rect 29236 20884 29242 20936
rect 29454 20884 29460 20936
rect 29512 20924 29518 20936
rect 29549 20927 29607 20933
rect 29549 20924 29561 20927
rect 29512 20896 29561 20924
rect 29512 20884 29518 20896
rect 29549 20893 29561 20896
rect 29595 20893 29607 20927
rect 29549 20887 29607 20893
rect 30009 20927 30067 20933
rect 30009 20893 30021 20927
rect 30055 20924 30067 20927
rect 30374 20924 30380 20936
rect 30055 20896 30380 20924
rect 30055 20893 30067 20896
rect 30009 20887 30067 20893
rect 30374 20884 30380 20896
rect 30432 20884 30438 20936
rect 30484 20924 30512 20964
rect 30834 20952 30840 21004
rect 30892 20992 30898 21004
rect 33704 20992 33732 21032
rect 36357 21029 36369 21063
rect 36403 21029 36415 21063
rect 36357 21023 36415 21029
rect 36372 20992 36400 21023
rect 37568 20992 37596 21088
rect 37918 21020 37924 21072
rect 37976 21060 37982 21072
rect 38105 21063 38163 21069
rect 38105 21060 38117 21063
rect 37976 21032 38117 21060
rect 37976 21020 37982 21032
rect 38105 21029 38117 21032
rect 38151 21029 38163 21063
rect 38105 21023 38163 21029
rect 38289 20995 38347 21001
rect 38289 20992 38301 20995
rect 30892 20964 31616 20992
rect 30892 20952 30898 20964
rect 31588 20936 31616 20964
rect 31864 20964 32444 20992
rect 31386 20924 31392 20936
rect 30484 20896 31392 20924
rect 31386 20884 31392 20896
rect 31444 20884 31450 20936
rect 31570 20884 31576 20936
rect 31628 20884 31634 20936
rect 31864 20933 31892 20964
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20893 31723 20927
rect 31665 20887 31723 20893
rect 31849 20927 31907 20933
rect 31849 20893 31861 20927
rect 31895 20893 31907 20927
rect 31849 20887 31907 20893
rect 26283 20828 27384 20856
rect 27525 20859 27583 20865
rect 26283 20825 26295 20828
rect 26237 20819 26295 20825
rect 27525 20825 27537 20859
rect 27571 20856 27583 20859
rect 27614 20856 27620 20868
rect 27571 20828 27620 20856
rect 27571 20825 27583 20828
rect 27525 20819 27583 20825
rect 27614 20816 27620 20828
rect 27672 20856 27678 20868
rect 27709 20859 27767 20865
rect 27709 20856 27721 20859
rect 27672 20828 27721 20856
rect 27672 20816 27678 20828
rect 27709 20825 27721 20828
rect 27755 20825 27767 20859
rect 27709 20819 27767 20825
rect 27893 20859 27951 20865
rect 27893 20825 27905 20859
rect 27939 20856 27951 20859
rect 29012 20856 29040 20884
rect 27939 20828 29040 20856
rect 29196 20856 29224 20884
rect 29825 20859 29883 20865
rect 29825 20856 29837 20859
rect 29196 20828 29837 20856
rect 27939 20825 27951 20828
rect 27893 20819 27951 20825
rect 29825 20825 29837 20828
rect 29871 20825 29883 20859
rect 29825 20819 29883 20825
rect 31481 20859 31539 20865
rect 31481 20825 31493 20859
rect 31527 20856 31539 20859
rect 31680 20856 31708 20887
rect 32306 20884 32312 20936
rect 32364 20884 32370 20936
rect 32416 20933 32444 20964
rect 33704 20964 34192 20992
rect 36372 20964 36676 20992
rect 37568 20964 38301 20992
rect 33704 20933 33732 20964
rect 32401 20927 32459 20933
rect 32401 20893 32413 20927
rect 32447 20924 32459 20927
rect 32677 20927 32735 20933
rect 32677 20924 32689 20927
rect 32447 20896 32689 20924
rect 32447 20893 32459 20896
rect 32401 20887 32459 20893
rect 32677 20893 32689 20896
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 33689 20927 33747 20933
rect 33689 20893 33701 20927
rect 33735 20893 33747 20927
rect 33689 20887 33747 20893
rect 33870 20884 33876 20936
rect 33928 20924 33934 20936
rect 34164 20933 34192 20964
rect 33965 20927 34023 20933
rect 33965 20924 33977 20927
rect 33928 20896 33977 20924
rect 33928 20884 33934 20896
rect 33965 20893 33977 20896
rect 34011 20893 34023 20927
rect 33965 20887 34023 20893
rect 34149 20927 34207 20933
rect 34149 20893 34161 20927
rect 34195 20893 34207 20927
rect 34149 20887 34207 20893
rect 35434 20884 35440 20936
rect 35492 20924 35498 20936
rect 35805 20927 35863 20933
rect 35805 20924 35817 20927
rect 35492 20896 35817 20924
rect 35492 20884 35498 20896
rect 35805 20893 35817 20896
rect 35851 20893 35863 20927
rect 35805 20887 35863 20893
rect 35986 20884 35992 20936
rect 36044 20884 36050 20936
rect 36538 20933 36544 20936
rect 36081 20927 36139 20933
rect 36081 20893 36093 20927
rect 36127 20893 36139 20927
rect 36081 20887 36139 20893
rect 36357 20927 36415 20933
rect 36357 20893 36369 20927
rect 36403 20893 36415 20927
rect 36357 20887 36415 20893
rect 36495 20927 36544 20933
rect 36495 20893 36507 20927
rect 36541 20893 36544 20927
rect 36495 20887 36544 20893
rect 31938 20856 31944 20868
rect 31527 20828 31944 20856
rect 31527 20825 31539 20828
rect 31481 20819 31539 20825
rect 31938 20816 31944 20828
rect 31996 20816 32002 20868
rect 32324 20856 32352 20884
rect 32582 20856 32588 20868
rect 32324 20828 32588 20856
rect 32582 20816 32588 20828
rect 32640 20816 32646 20868
rect 32861 20859 32919 20865
rect 32861 20825 32873 20859
rect 32907 20825 32919 20859
rect 32861 20819 32919 20825
rect 19107 20760 19656 20788
rect 19107 20757 19119 20760
rect 19061 20751 19119 20757
rect 22186 20748 22192 20800
rect 22244 20748 22250 20800
rect 26326 20748 26332 20800
rect 26384 20788 26390 20800
rect 26697 20791 26755 20797
rect 26697 20788 26709 20791
rect 26384 20760 26709 20788
rect 26384 20748 26390 20760
rect 26697 20757 26709 20760
rect 26743 20757 26755 20791
rect 26697 20751 26755 20757
rect 28442 20748 28448 20800
rect 28500 20748 28506 20800
rect 30190 20748 30196 20800
rect 30248 20748 30254 20800
rect 31570 20748 31576 20800
rect 31628 20788 31634 20800
rect 32306 20788 32312 20800
rect 31628 20760 32312 20788
rect 31628 20748 31634 20760
rect 32306 20748 32312 20760
rect 32364 20788 32370 20800
rect 32876 20788 32904 20819
rect 33042 20816 33048 20868
rect 33100 20816 33106 20868
rect 32364 20760 32904 20788
rect 32364 20748 32370 20760
rect 35986 20748 35992 20800
rect 36044 20788 36050 20800
rect 36096 20788 36124 20887
rect 36044 20760 36124 20788
rect 36372 20788 36400 20887
rect 36538 20884 36544 20887
rect 36596 20884 36602 20936
rect 36648 20933 36676 20964
rect 36633 20927 36691 20933
rect 36633 20893 36645 20927
rect 36679 20893 36691 20927
rect 36633 20887 36691 20893
rect 36722 20884 36728 20936
rect 36780 20924 36786 20936
rect 36817 20927 36875 20933
rect 36817 20924 36829 20927
rect 36780 20896 36829 20924
rect 36780 20884 36786 20896
rect 36817 20893 36829 20896
rect 36863 20893 36875 20927
rect 37826 20924 37832 20936
rect 36817 20887 36875 20893
rect 37660 20896 37832 20924
rect 37537 20859 37595 20865
rect 37537 20825 37549 20859
rect 37583 20856 37595 20859
rect 37660 20856 37688 20896
rect 37826 20884 37832 20896
rect 37884 20884 37890 20936
rect 37936 20933 37964 20964
rect 38289 20961 38301 20964
rect 38335 20961 38347 20995
rect 38289 20955 38347 20961
rect 37921 20927 37979 20933
rect 37921 20893 37933 20927
rect 37967 20893 37979 20927
rect 37921 20887 37979 20893
rect 38102 20884 38108 20936
rect 38160 20884 38166 20936
rect 38194 20884 38200 20936
rect 38252 20884 38258 20936
rect 38378 20884 38384 20936
rect 38436 20884 38442 20936
rect 37583 20828 37688 20856
rect 37583 20825 37595 20828
rect 37537 20819 37595 20825
rect 37734 20816 37740 20868
rect 37792 20856 37798 20868
rect 38120 20856 38148 20884
rect 37792 20828 38148 20856
rect 37792 20816 37798 20828
rect 36446 20788 36452 20800
rect 36372 20760 36452 20788
rect 36044 20748 36050 20760
rect 36446 20748 36452 20760
rect 36504 20788 36510 20800
rect 37369 20791 37427 20797
rect 37369 20788 37381 20791
rect 36504 20760 37381 20788
rect 36504 20748 36510 20760
rect 37369 20757 37381 20760
rect 37415 20757 37427 20791
rect 37369 20751 37427 20757
rect 1104 20698 38824 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 38824 20698
rect 1104 20624 38824 20646
rect 3418 20544 3424 20596
rect 3476 20584 3482 20596
rect 3476 20556 4936 20584
rect 3476 20544 3482 20556
rect 2501 20519 2559 20525
rect 2501 20485 2513 20519
rect 2547 20516 2559 20519
rect 2774 20516 2780 20528
rect 2547 20488 2780 20516
rect 2547 20485 2559 20488
rect 2501 20479 2559 20485
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 4798 20516 4804 20528
rect 3726 20488 4804 20516
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 4908 20525 4936 20556
rect 5350 20544 5356 20596
rect 5408 20544 5414 20596
rect 7929 20587 7987 20593
rect 7929 20553 7941 20587
rect 7975 20584 7987 20587
rect 8570 20584 8576 20596
rect 7975 20556 8576 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 9582 20584 9588 20596
rect 9048 20556 9588 20584
rect 4893 20519 4951 20525
rect 4893 20485 4905 20519
rect 4939 20516 4951 20519
rect 8018 20516 8024 20528
rect 4939 20488 8024 20516
rect 4939 20485 4951 20488
rect 4893 20479 4951 20485
rect 8018 20476 8024 20488
rect 8076 20476 8082 20528
rect 9048 20516 9076 20556
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 11606 20544 11612 20596
rect 11664 20544 11670 20596
rect 12158 20544 12164 20596
rect 12216 20584 12222 20596
rect 12894 20584 12900 20596
rect 12216 20556 12900 20584
rect 12216 20544 12222 20556
rect 8970 20488 9076 20516
rect 9398 20476 9404 20528
rect 9456 20476 9462 20528
rect 2038 20408 2044 20460
rect 2096 20448 2102 20460
rect 2225 20451 2283 20457
rect 2225 20448 2237 20451
rect 2096 20420 2237 20448
rect 2096 20408 2102 20420
rect 2225 20417 2237 20420
rect 2271 20417 2283 20451
rect 2225 20411 2283 20417
rect 5534 20408 5540 20460
rect 5592 20408 5598 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5644 20420 5825 20448
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 3804 20352 4629 20380
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 3804 20244 3832 20352
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 4617 20343 4675 20349
rect 4706 20340 4712 20392
rect 4764 20380 4770 20392
rect 5644 20380 5672 20420
rect 5813 20417 5825 20420
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20417 6055 20451
rect 5997 20411 6055 20417
rect 6917 20451 6975 20457
rect 6917 20417 6929 20451
rect 6963 20448 6975 20451
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 6963 20420 7205 20448
rect 6963 20417 6975 20420
rect 6917 20411 6975 20417
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 4764 20352 5672 20380
rect 4764 20340 4770 20352
rect 5718 20340 5724 20392
rect 5776 20380 5782 20392
rect 5905 20383 5963 20389
rect 5905 20380 5917 20383
rect 5776 20352 5917 20380
rect 5776 20340 5782 20352
rect 5905 20349 5917 20352
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 3878 20272 3884 20324
rect 3936 20312 3942 20324
rect 6012 20312 6040 20411
rect 7742 20408 7748 20460
rect 7800 20408 7806 20460
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 12268 20457 12296 20556
rect 12894 20544 12900 20556
rect 12952 20584 12958 20596
rect 13722 20584 13728 20596
rect 12952 20556 13728 20584
rect 12952 20544 12958 20556
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 15933 20587 15991 20593
rect 14292 20556 15240 20584
rect 12805 20519 12863 20525
rect 12805 20485 12817 20519
rect 12851 20516 12863 20519
rect 14292 20516 14320 20556
rect 15212 20516 15240 20556
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 16850 20584 16856 20596
rect 15979 20556 16856 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 16850 20544 16856 20556
rect 16908 20584 16914 20596
rect 17313 20587 17371 20593
rect 17313 20584 17325 20587
rect 16908 20556 17325 20584
rect 16908 20544 16914 20556
rect 17313 20553 17325 20556
rect 17359 20553 17371 20587
rect 17313 20547 17371 20553
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 18230 20584 18236 20596
rect 17552 20556 18236 20584
rect 17552 20544 17558 20556
rect 18230 20544 18236 20556
rect 18288 20544 18294 20596
rect 18325 20587 18383 20593
rect 18325 20553 18337 20587
rect 18371 20584 18383 20587
rect 19518 20584 19524 20596
rect 18371 20556 19524 20584
rect 18371 20553 18383 20556
rect 18325 20547 18383 20553
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 25317 20587 25375 20593
rect 25317 20553 25329 20587
rect 25363 20584 25375 20587
rect 25866 20584 25872 20596
rect 25363 20556 25872 20584
rect 25363 20553 25375 20556
rect 25317 20547 25375 20553
rect 25866 20544 25872 20556
rect 25924 20544 25930 20596
rect 25958 20544 25964 20596
rect 26016 20544 26022 20596
rect 26602 20544 26608 20596
rect 26660 20584 26666 20596
rect 27249 20587 27307 20593
rect 27249 20584 27261 20587
rect 26660 20556 27261 20584
rect 26660 20544 26666 20556
rect 27249 20553 27261 20556
rect 27295 20584 27307 20587
rect 27522 20584 27528 20596
rect 27295 20556 27528 20584
rect 27295 20553 27307 20556
rect 27249 20547 27307 20553
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 34422 20544 34428 20596
rect 34480 20544 34486 20596
rect 35434 20544 35440 20596
rect 35492 20584 35498 20596
rect 35529 20587 35587 20593
rect 35529 20584 35541 20587
rect 35492 20556 35541 20584
rect 35492 20544 35498 20556
rect 35529 20553 35541 20556
rect 35575 20553 35587 20587
rect 35529 20547 35587 20553
rect 36170 20544 36176 20596
rect 36228 20584 36234 20596
rect 37093 20587 37151 20593
rect 37093 20584 37105 20587
rect 36228 20556 37105 20584
rect 36228 20544 36234 20556
rect 37093 20553 37105 20556
rect 37139 20553 37151 20587
rect 37093 20547 37151 20553
rect 37826 20544 37832 20596
rect 37884 20544 37890 20596
rect 16393 20519 16451 20525
rect 12851 20488 14320 20516
rect 15134 20488 16344 20516
rect 12851 20485 12863 20488
rect 12805 20479 12863 20485
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20417 12311 20451
rect 12253 20411 12311 20417
rect 12526 20408 12532 20460
rect 12584 20448 12590 20460
rect 13633 20451 13691 20457
rect 13633 20448 13645 20451
rect 12584 20420 13645 20448
rect 12584 20408 12590 20420
rect 13633 20417 13645 20420
rect 13679 20417 13691 20451
rect 13633 20411 13691 20417
rect 15838 20408 15844 20460
rect 15896 20408 15902 20460
rect 16316 20448 16344 20488
rect 16393 20485 16405 20519
rect 16439 20516 16451 20519
rect 17681 20519 17739 20525
rect 17681 20516 17693 20519
rect 16439 20488 17693 20516
rect 16439 20485 16451 20488
rect 16393 20479 16451 20485
rect 16485 20451 16543 20457
rect 16316 20420 16436 20448
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7466 20380 7472 20392
rect 7055 20352 7472 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7466 20340 7472 20352
rect 7524 20380 7530 20392
rect 7650 20380 7656 20392
rect 7524 20352 7656 20380
rect 7524 20340 7530 20352
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13035 20352 13768 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 3936 20284 6040 20312
rect 3936 20272 3942 20284
rect 3973 20247 4031 20253
rect 3973 20244 3985 20247
rect 3752 20216 3985 20244
rect 3752 20204 3758 20216
rect 3973 20213 3985 20216
rect 4019 20213 4031 20247
rect 3973 20207 4031 20213
rect 4062 20204 4068 20256
rect 4120 20204 4126 20256
rect 4982 20204 4988 20256
rect 5040 20204 5046 20256
rect 6549 20247 6607 20253
rect 6549 20213 6561 20247
rect 6595 20244 6607 20247
rect 6638 20244 6644 20256
rect 6595 20216 6644 20244
rect 6595 20213 6607 20216
rect 6549 20207 6607 20213
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 13541 20247 13599 20253
rect 13541 20244 13553 20247
rect 13504 20216 13553 20244
rect 13504 20204 13510 20216
rect 13541 20213 13553 20216
rect 13587 20213 13599 20247
rect 13740 20244 13768 20352
rect 13906 20340 13912 20392
rect 13964 20340 13970 20392
rect 15654 20340 15660 20392
rect 15712 20380 15718 20392
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 15712 20352 16037 20380
rect 15712 20340 15718 20352
rect 16025 20349 16037 20352
rect 16071 20349 16083 20383
rect 16408 20380 16436 20420
rect 16485 20417 16497 20451
rect 16531 20448 16543 20451
rect 16574 20448 16580 20460
rect 16531 20420 16580 20448
rect 16531 20417 16543 20420
rect 16485 20411 16543 20417
rect 16574 20408 16580 20420
rect 16632 20448 16638 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16632 20420 16681 20448
rect 16632 20408 16638 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 17310 20380 17316 20392
rect 16408 20352 17316 20380
rect 16025 20343 16083 20349
rect 17310 20340 17316 20352
rect 17368 20340 17374 20392
rect 17512 20380 17540 20488
rect 17681 20485 17693 20488
rect 17727 20485 17739 20519
rect 17681 20479 17739 20485
rect 17954 20476 17960 20528
rect 18012 20516 18018 20528
rect 18141 20519 18199 20525
rect 18141 20516 18153 20519
rect 18012 20488 18153 20516
rect 18012 20476 18018 20488
rect 18141 20485 18153 20488
rect 18187 20485 18199 20519
rect 19242 20516 19248 20528
rect 18141 20479 18199 20485
rect 18248 20488 18644 20516
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20448 17647 20451
rect 18248 20448 18276 20488
rect 18616 20460 18644 20488
rect 19076 20488 19248 20516
rect 17635 20420 18276 20448
rect 17635 20417 17647 20420
rect 17589 20411 17647 20417
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 18598 20408 18604 20460
rect 18656 20408 18662 20460
rect 18874 20457 18880 20460
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 18831 20451 18880 20457
rect 18831 20417 18843 20451
rect 18877 20417 18880 20451
rect 18831 20411 18880 20417
rect 18708 20380 18736 20411
rect 18874 20408 18880 20411
rect 18932 20408 18938 20460
rect 19076 20457 19104 20488
rect 19242 20476 19248 20488
rect 19300 20476 19306 20528
rect 20346 20476 20352 20528
rect 20404 20476 20410 20528
rect 21174 20476 21180 20528
rect 21232 20476 21238 20528
rect 21542 20476 21548 20528
rect 21600 20516 21606 20528
rect 21600 20488 22581 20516
rect 21600 20476 21606 20488
rect 19061 20451 19119 20457
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 20990 20408 20996 20460
rect 21048 20448 21054 20460
rect 22112 20457 22140 20488
rect 21453 20451 21511 20457
rect 21453 20448 21465 20451
rect 21048 20420 21465 20448
rect 21048 20408 21054 20420
rect 21453 20417 21465 20420
rect 21499 20448 21511 20451
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21499 20420 21833 20448
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20417 22155 20451
rect 22097 20411 22155 20417
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 17512 20352 18736 20380
rect 18138 20272 18144 20324
rect 18196 20272 18202 20324
rect 18708 20312 18736 20352
rect 18969 20383 19027 20389
rect 18969 20349 18981 20383
rect 19015 20349 19027 20383
rect 18969 20343 19027 20349
rect 19337 20383 19395 20389
rect 19337 20349 19349 20383
rect 19383 20380 19395 20383
rect 19794 20380 19800 20392
rect 19383 20352 19800 20380
rect 19383 20349 19395 20352
rect 19337 20343 19395 20349
rect 18782 20312 18788 20324
rect 18708 20284 18788 20312
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 14366 20244 14372 20256
rect 13740 20216 14372 20244
rect 13541 20207 13599 20213
rect 14366 20204 14372 20216
rect 14424 20244 14430 20256
rect 15381 20247 15439 20253
rect 15381 20244 15393 20247
rect 14424 20216 15393 20244
rect 14424 20204 14430 20216
rect 15381 20213 15393 20216
rect 15427 20213 15439 20247
rect 15381 20207 15439 20213
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 17402 20204 17408 20256
rect 17460 20204 17466 20256
rect 18984 20244 19012 20343
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 20070 20340 20076 20392
rect 20128 20380 20134 20392
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 20128 20352 21281 20380
rect 20128 20340 20134 20352
rect 21269 20349 21281 20352
rect 21315 20380 21327 20383
rect 21542 20380 21548 20392
rect 21315 20352 21548 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 21542 20340 21548 20352
rect 21600 20340 21606 20392
rect 21910 20340 21916 20392
rect 21968 20340 21974 20392
rect 22278 20340 22284 20392
rect 22336 20380 22342 20392
rect 22394 20380 22422 20411
rect 22336 20352 22422 20380
rect 22465 20383 22523 20389
rect 22336 20340 22342 20352
rect 22465 20349 22477 20383
rect 22511 20349 22523 20383
rect 22553 20380 22581 20488
rect 23842 20476 23848 20528
rect 23900 20476 23906 20528
rect 24302 20476 24308 20528
rect 24360 20476 24366 20528
rect 25498 20476 25504 20528
rect 25556 20476 25562 20528
rect 25685 20519 25743 20525
rect 25685 20485 25697 20519
rect 25731 20516 25743 20519
rect 25976 20516 26004 20544
rect 25731 20488 26004 20516
rect 27065 20519 27123 20525
rect 25731 20485 25743 20488
rect 25685 20479 25743 20485
rect 27065 20485 27077 20519
rect 27111 20516 27123 20519
rect 29270 20516 29276 20528
rect 27111 20488 29276 20516
rect 27111 20485 27123 20488
rect 27065 20479 27123 20485
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 23109 20451 23167 20457
rect 23109 20448 23121 20451
rect 22704 20420 23121 20448
rect 22704 20408 22710 20420
rect 23109 20417 23121 20420
rect 23155 20417 23167 20451
rect 23109 20411 23167 20417
rect 23201 20451 23259 20457
rect 23201 20417 23213 20451
rect 23247 20417 23259 20451
rect 23201 20411 23259 20417
rect 22925 20383 22983 20389
rect 22925 20380 22937 20383
rect 22553 20352 22937 20380
rect 22465 20343 22523 20349
rect 22925 20349 22937 20352
rect 22971 20380 22983 20383
rect 23014 20380 23020 20392
rect 22971 20352 23020 20380
rect 22971 20349 22983 20352
rect 22925 20343 22983 20349
rect 21634 20272 21640 20324
rect 21692 20272 21698 20324
rect 21928 20312 21956 20340
rect 22480 20312 22508 20343
rect 23014 20340 23020 20352
rect 23072 20340 23078 20392
rect 23216 20380 23244 20411
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23474 20408 23480 20460
rect 23532 20408 23538 20460
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20448 26203 20451
rect 26234 20448 26240 20460
rect 26191 20420 26240 20448
rect 26191 20417 26203 20420
rect 26145 20411 26203 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 26326 20408 26332 20460
rect 26384 20408 26390 20460
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20417 26479 20451
rect 26421 20411 26479 20417
rect 26513 20451 26571 20457
rect 26513 20417 26525 20451
rect 26559 20448 26571 20451
rect 27080 20448 27108 20479
rect 29270 20476 29276 20488
rect 29328 20476 29334 20528
rect 29641 20519 29699 20525
rect 29641 20485 29653 20519
rect 29687 20516 29699 20519
rect 31846 20516 31852 20528
rect 29687 20488 31852 20516
rect 29687 20485 29699 20488
rect 29641 20479 29699 20485
rect 31846 20476 31852 20488
rect 31904 20516 31910 20528
rect 33042 20516 33048 20528
rect 31904 20488 33048 20516
rect 31904 20476 31910 20488
rect 33042 20476 33048 20488
rect 33100 20476 33106 20528
rect 36078 20476 36084 20528
rect 36136 20516 36142 20528
rect 36136 20488 36952 20516
rect 36136 20476 36142 20488
rect 26559 20420 27108 20448
rect 27157 20451 27215 20457
rect 26559 20417 26571 20420
rect 26513 20411 26571 20417
rect 27157 20417 27169 20451
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 23382 20380 23388 20392
rect 23216 20352 23388 20380
rect 23382 20340 23388 20352
rect 23440 20340 23446 20392
rect 23569 20383 23627 20389
rect 23569 20349 23581 20383
rect 23615 20349 23627 20383
rect 23569 20343 23627 20349
rect 21744 20284 21956 20312
rect 22204 20284 22508 20312
rect 19334 20244 19340 20256
rect 18984 20216 19340 20244
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 20809 20247 20867 20253
rect 20809 20244 20821 20247
rect 19576 20216 20821 20244
rect 19576 20204 19582 20216
rect 20809 20213 20821 20216
rect 20855 20244 20867 20247
rect 21177 20247 21235 20253
rect 21177 20244 21189 20247
rect 20855 20216 21189 20244
rect 20855 20213 20867 20216
rect 20809 20207 20867 20213
rect 21177 20213 21189 20216
rect 21223 20244 21235 20247
rect 21744 20244 21772 20284
rect 21223 20216 21772 20244
rect 21223 20213 21235 20216
rect 21177 20207 21235 20213
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 22204 20244 22232 20284
rect 21968 20216 22232 20244
rect 22281 20247 22339 20253
rect 21968 20204 21974 20216
rect 22281 20213 22293 20247
rect 22327 20244 22339 20247
rect 22370 20244 22376 20256
rect 22327 20216 22376 20244
rect 22327 20213 22339 20216
rect 22281 20207 22339 20213
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 22554 20204 22560 20256
rect 22612 20204 22618 20256
rect 22738 20204 22744 20256
rect 22796 20204 22802 20256
rect 23014 20204 23020 20256
rect 23072 20204 23078 20256
rect 23584 20244 23612 20343
rect 26050 20340 26056 20392
rect 26108 20380 26114 20392
rect 26436 20380 26464 20411
rect 26108 20352 26464 20380
rect 27172 20380 27200 20411
rect 27246 20408 27252 20460
rect 27304 20408 27310 20460
rect 27433 20451 27491 20457
rect 27433 20417 27445 20451
rect 27479 20448 27491 20451
rect 27614 20448 27620 20460
rect 27479 20420 27620 20448
rect 27479 20417 27491 20420
rect 27433 20411 27491 20417
rect 27614 20408 27620 20420
rect 27672 20448 27678 20460
rect 27893 20451 27951 20457
rect 27893 20448 27905 20451
rect 27672 20420 27905 20448
rect 27672 20408 27678 20420
rect 27893 20417 27905 20420
rect 27939 20417 27951 20451
rect 27893 20411 27951 20417
rect 28077 20451 28135 20457
rect 28077 20417 28089 20451
rect 28123 20448 28135 20451
rect 28994 20448 29000 20460
rect 28123 20420 29000 20448
rect 28123 20417 28135 20420
rect 28077 20411 28135 20417
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 29362 20408 29368 20460
rect 29420 20448 29426 20460
rect 29546 20448 29552 20460
rect 29420 20420 29552 20448
rect 29420 20408 29426 20420
rect 29546 20408 29552 20420
rect 29604 20448 29610 20460
rect 30009 20451 30067 20457
rect 30009 20448 30021 20451
rect 29604 20420 30021 20448
rect 29604 20408 29610 20420
rect 30009 20417 30021 20420
rect 30055 20417 30067 20451
rect 30009 20411 30067 20417
rect 30193 20451 30251 20457
rect 30193 20417 30205 20451
rect 30239 20448 30251 20451
rect 31573 20451 31631 20457
rect 31573 20448 31585 20451
rect 30239 20420 31585 20448
rect 30239 20417 30251 20420
rect 30193 20411 30251 20417
rect 31573 20417 31585 20420
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20448 31815 20451
rect 31938 20448 31944 20460
rect 31803 20420 31944 20448
rect 31803 20417 31815 20420
rect 31757 20411 31815 20417
rect 27798 20380 27804 20392
rect 27172 20352 27804 20380
rect 26108 20340 26114 20352
rect 27798 20340 27804 20352
rect 27856 20340 27862 20392
rect 27985 20383 28043 20389
rect 27985 20349 27997 20383
rect 28031 20380 28043 20383
rect 28350 20380 28356 20392
rect 28031 20352 28356 20380
rect 28031 20349 28043 20352
rect 27985 20343 28043 20349
rect 28350 20340 28356 20352
rect 28408 20380 28414 20392
rect 29730 20380 29736 20392
rect 28408 20352 29736 20380
rect 28408 20340 28414 20352
rect 29730 20340 29736 20352
rect 29788 20380 29794 20392
rect 30208 20380 30236 20411
rect 31938 20408 31944 20420
rect 31996 20408 32002 20460
rect 33505 20451 33563 20457
rect 33505 20417 33517 20451
rect 33551 20448 33563 20451
rect 33551 20420 33732 20448
rect 33551 20417 33563 20420
rect 33505 20411 33563 20417
rect 29788 20352 30236 20380
rect 29788 20340 29794 20352
rect 33594 20340 33600 20392
rect 33652 20340 33658 20392
rect 33704 20324 33732 20420
rect 33962 20408 33968 20460
rect 34020 20408 34026 20460
rect 34057 20451 34115 20457
rect 34057 20417 34069 20451
rect 34103 20417 34115 20451
rect 34057 20411 34115 20417
rect 33870 20340 33876 20392
rect 33928 20340 33934 20392
rect 34072 20380 34100 20411
rect 34146 20408 34152 20460
rect 34204 20448 34210 20460
rect 34241 20451 34299 20457
rect 34241 20448 34253 20451
rect 34204 20420 34253 20448
rect 34204 20408 34210 20420
rect 34241 20417 34253 20420
rect 34287 20417 34299 20451
rect 34241 20411 34299 20417
rect 35897 20451 35955 20457
rect 35897 20417 35909 20451
rect 35943 20417 35955 20451
rect 35897 20411 35955 20417
rect 34072 20352 34192 20380
rect 33686 20272 33692 20324
rect 33744 20312 33750 20324
rect 34164 20312 34192 20352
rect 35802 20340 35808 20392
rect 35860 20340 35866 20392
rect 35912 20380 35940 20411
rect 36170 20408 36176 20460
rect 36228 20448 36234 20460
rect 36924 20457 36952 20488
rect 37458 20476 37464 20528
rect 37516 20476 37522 20528
rect 37642 20476 37648 20528
rect 37700 20476 37706 20528
rect 36357 20451 36415 20457
rect 36357 20448 36369 20451
rect 36228 20420 36369 20448
rect 36228 20408 36234 20420
rect 36357 20417 36369 20420
rect 36403 20448 36415 20451
rect 36633 20451 36691 20457
rect 36633 20448 36645 20451
rect 36403 20420 36645 20448
rect 36403 20417 36415 20420
rect 36357 20411 36415 20417
rect 36633 20417 36645 20420
rect 36679 20417 36691 20451
rect 36633 20411 36691 20417
rect 36909 20451 36967 20457
rect 36909 20417 36921 20451
rect 36955 20417 36967 20451
rect 36909 20411 36967 20417
rect 35986 20380 35992 20392
rect 35912 20352 35992 20380
rect 35986 20340 35992 20352
rect 36044 20340 36050 20392
rect 36449 20383 36507 20389
rect 36449 20349 36461 20383
rect 36495 20349 36507 20383
rect 36449 20343 36507 20349
rect 36354 20312 36360 20324
rect 33744 20284 36360 20312
rect 33744 20272 33750 20284
rect 36354 20272 36360 20284
rect 36412 20272 36418 20324
rect 36464 20312 36492 20343
rect 36464 20284 36768 20312
rect 36740 20256 36768 20284
rect 24946 20244 24952 20256
rect 23584 20216 24952 20244
rect 24946 20204 24952 20216
rect 25004 20204 25010 20256
rect 26786 20204 26792 20256
rect 26844 20204 26850 20256
rect 29549 20247 29607 20253
rect 29549 20213 29561 20247
rect 29595 20244 29607 20247
rect 29638 20244 29644 20256
rect 29595 20216 29644 20244
rect 29595 20213 29607 20216
rect 29549 20207 29607 20213
rect 29638 20204 29644 20216
rect 29696 20204 29702 20256
rect 30098 20204 30104 20256
rect 30156 20244 30162 20256
rect 30193 20247 30251 20253
rect 30193 20244 30205 20247
rect 30156 20216 30205 20244
rect 30156 20204 30162 20216
rect 30193 20213 30205 20216
rect 30239 20213 30251 20247
rect 30193 20207 30251 20213
rect 31570 20204 31576 20256
rect 31628 20204 31634 20256
rect 35894 20204 35900 20256
rect 35952 20204 35958 20256
rect 35986 20204 35992 20256
rect 36044 20204 36050 20256
rect 36722 20204 36728 20256
rect 36780 20204 36786 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 3694 20040 3700 20052
rect 3467 20012 3700 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 3786 20000 3792 20052
rect 3844 20000 3850 20052
rect 4433 20043 4491 20049
rect 4433 20009 4445 20043
rect 4479 20040 4491 20043
rect 5534 20040 5540 20052
rect 4479 20012 5540 20040
rect 4479 20009 4491 20012
rect 4433 20003 4491 20009
rect 5534 20000 5540 20012
rect 5592 20000 5598 20052
rect 7742 20000 7748 20052
rect 7800 20040 7806 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7800 20012 8125 20040
rect 7800 20000 7806 20012
rect 8113 20009 8125 20012
rect 8159 20040 8171 20043
rect 8389 20043 8447 20049
rect 8389 20040 8401 20043
rect 8159 20012 8401 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8389 20009 8401 20012
rect 8435 20009 8447 20043
rect 8389 20003 8447 20009
rect 8478 20000 8484 20052
rect 8536 20040 8542 20052
rect 8573 20043 8631 20049
rect 8573 20040 8585 20043
rect 8536 20012 8585 20040
rect 8536 20000 8542 20012
rect 8573 20009 8585 20012
rect 8619 20009 8631 20043
rect 8573 20003 8631 20009
rect 13906 20000 13912 20052
rect 13964 20000 13970 20052
rect 14274 20000 14280 20052
rect 14332 20000 14338 20052
rect 16666 20040 16672 20052
rect 15856 20012 16672 20040
rect 3237 19975 3295 19981
rect 3237 19941 3249 19975
rect 3283 19972 3295 19975
rect 3878 19972 3884 19984
rect 3283 19944 3884 19972
rect 3283 19941 3295 19944
rect 3237 19935 3295 19941
rect 3878 19932 3884 19944
rect 3936 19932 3942 19984
rect 13372 19944 13584 19972
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2038 19904 2044 19916
rect 1443 19876 2044 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 5684 19876 6285 19904
rect 5684 19864 5690 19876
rect 6273 19873 6285 19876
rect 6319 19904 6331 19907
rect 6365 19907 6423 19913
rect 6365 19904 6377 19907
rect 6319 19876 6377 19904
rect 6319 19873 6331 19876
rect 6273 19867 6331 19873
rect 6365 19873 6377 19876
rect 6411 19873 6423 19907
rect 6365 19867 6423 19873
rect 6638 19864 6644 19916
rect 6696 19864 6702 19916
rect 10594 19864 10600 19916
rect 10652 19864 10658 19916
rect 12526 19864 12532 19916
rect 12584 19864 12590 19916
rect 13372 19913 13400 19944
rect 13357 19907 13415 19913
rect 13357 19873 13369 19907
rect 13403 19873 13415 19907
rect 13357 19867 13415 19873
rect 13446 19864 13452 19916
rect 13504 19864 13510 19916
rect 13556 19904 13584 19944
rect 14090 19932 14096 19984
rect 14148 19972 14154 19984
rect 15856 19972 15884 20012
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 17497 20043 17555 20049
rect 17497 20009 17509 20043
rect 17543 20040 17555 20043
rect 17954 20040 17960 20052
rect 17543 20012 17960 20040
rect 17543 20009 17555 20012
rect 17497 20003 17555 20009
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 19794 20000 19800 20052
rect 19852 20000 19858 20052
rect 21450 20000 21456 20052
rect 21508 20040 21514 20052
rect 21726 20040 21732 20052
rect 21508 20012 21732 20040
rect 21508 20000 21514 20012
rect 21726 20000 21732 20012
rect 21784 20000 21790 20052
rect 22833 20043 22891 20049
rect 22833 20009 22845 20043
rect 22879 20040 22891 20043
rect 22879 20012 23244 20040
rect 22879 20009 22891 20012
rect 22833 20003 22891 20009
rect 14148 19944 15884 19972
rect 22925 19975 22983 19981
rect 14148 19932 14154 19944
rect 22925 19941 22937 19975
rect 22971 19941 22983 19975
rect 22925 19935 22983 19941
rect 15654 19904 15660 19916
rect 13556 19876 15660 19904
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16390 19904 16396 19916
rect 16071 19876 16396 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19904 17739 19907
rect 18598 19904 18604 19916
rect 17727 19876 18604 19904
rect 17727 19873 17739 19876
rect 17681 19867 17739 19873
rect 18598 19864 18604 19876
rect 18656 19904 18662 19916
rect 18656 19876 19472 19904
rect 18656 19864 18662 19876
rect 2774 19796 2780 19848
rect 2832 19796 2838 19848
rect 3970 19796 3976 19848
rect 4028 19796 4034 19848
rect 4249 19839 4307 19845
rect 4249 19805 4261 19839
rect 4295 19836 4307 19839
rect 4706 19836 4712 19848
rect 4295 19808 4712 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 8570 19796 8576 19848
rect 8628 19796 8634 19848
rect 12544 19836 12572 19864
rect 14369 19839 14427 19845
rect 14369 19836 14381 19839
rect 12544 19808 14381 19836
rect 14369 19805 14381 19808
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 1670 19728 1676 19780
rect 1728 19728 1734 19780
rect 3510 19768 3516 19780
rect 3160 19740 3516 19768
rect 3160 19709 3188 19740
rect 3510 19728 3516 19740
rect 3568 19768 3574 19780
rect 3605 19771 3663 19777
rect 3605 19768 3617 19771
rect 3568 19740 3617 19768
rect 3568 19728 3574 19740
rect 3605 19737 3617 19740
rect 3651 19737 3663 19771
rect 3605 19731 3663 19737
rect 3878 19728 3884 19780
rect 3936 19768 3942 19780
rect 4065 19771 4123 19777
rect 4065 19768 4077 19771
rect 3936 19740 4077 19768
rect 3936 19728 3942 19740
rect 4065 19737 4077 19740
rect 4111 19737 4123 19771
rect 4065 19731 4123 19737
rect 4982 19728 4988 19780
rect 5040 19728 5046 19780
rect 5994 19728 6000 19780
rect 6052 19728 6058 19780
rect 7926 19768 7932 19780
rect 7866 19740 7932 19768
rect 7926 19728 7932 19740
rect 7984 19728 7990 19780
rect 8205 19771 8263 19777
rect 8205 19737 8217 19771
rect 8251 19768 8263 19771
rect 8588 19768 8616 19796
rect 8251 19740 8616 19768
rect 8251 19737 8263 19740
rect 8205 19731 8263 19737
rect 11790 19728 11796 19780
rect 11848 19728 11854 19780
rect 12250 19728 12256 19780
rect 12308 19728 12314 19780
rect 14384 19768 14412 19799
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 14700 19808 14749 19836
rect 14700 19796 14706 19808
rect 14737 19805 14749 19808
rect 14783 19805 14795 19839
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 14737 19799 14795 19805
rect 15488 19808 15761 19836
rect 15488 19777 15516 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 17586 19796 17592 19848
rect 17644 19796 17650 19848
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 15473 19771 15531 19777
rect 15473 19768 15485 19771
rect 14384 19740 15485 19768
rect 14752 19712 14780 19740
rect 15473 19737 15485 19740
rect 15519 19737 15531 19771
rect 17494 19768 17500 19780
rect 17250 19740 17500 19768
rect 15473 19731 15531 19737
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 17678 19728 17684 19780
rect 17736 19768 17742 19780
rect 17788 19768 17816 19799
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19444 19845 19472 19876
rect 21634 19864 21640 19916
rect 21692 19904 21698 19916
rect 22189 19907 22247 19913
rect 22189 19904 22201 19907
rect 21692 19876 22201 19904
rect 21692 19864 21698 19876
rect 22189 19873 22201 19876
rect 22235 19873 22247 19907
rect 22189 19867 22247 19873
rect 22649 19907 22707 19913
rect 22649 19873 22661 19907
rect 22695 19904 22707 19907
rect 22940 19904 22968 19935
rect 22695 19876 22968 19904
rect 23216 19904 23244 20012
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 23477 20043 23535 20049
rect 23477 20040 23489 20043
rect 23440 20012 23489 20040
rect 23440 20000 23446 20012
rect 23477 20009 23489 20012
rect 23523 20009 23535 20043
rect 23477 20003 23535 20009
rect 28074 20000 28080 20052
rect 28132 20000 28138 20052
rect 29178 20000 29184 20052
rect 29236 20000 29242 20052
rect 29638 20000 29644 20052
rect 29696 20040 29702 20052
rect 29696 20012 36400 20040
rect 29696 20000 29702 20012
rect 23658 19932 23664 19984
rect 23716 19972 23722 19984
rect 29822 19972 29828 19984
rect 23716 19944 29828 19972
rect 23716 19932 23722 19944
rect 29822 19932 29828 19944
rect 29880 19932 29886 19984
rect 31846 19981 31852 19984
rect 31803 19975 31852 19981
rect 31803 19941 31815 19975
rect 31849 19941 31852 19975
rect 31803 19935 31852 19941
rect 31846 19932 31852 19935
rect 31904 19932 31910 19984
rect 33594 19932 33600 19984
rect 33652 19932 33658 19984
rect 33962 19932 33968 19984
rect 34020 19932 34026 19984
rect 35802 19932 35808 19984
rect 35860 19972 35866 19984
rect 35860 19944 36308 19972
rect 35860 19932 35866 19944
rect 23474 19904 23480 19916
rect 23216 19876 23480 19904
rect 22695 19873 22707 19876
rect 22649 19867 22707 19873
rect 23474 19864 23480 19876
rect 23532 19864 23538 19916
rect 25976 19876 27844 19904
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18748 19808 19257 19836
rect 18748 19796 18754 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 19518 19796 19524 19848
rect 19576 19796 19582 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 21729 19839 21787 19845
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 17736 19740 17816 19768
rect 17736 19728 17742 19740
rect 18874 19728 18880 19780
rect 18932 19768 18938 19780
rect 19628 19768 19656 19799
rect 18932 19740 19656 19768
rect 21744 19768 21772 19799
rect 21818 19796 21824 19848
rect 21876 19796 21882 19848
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19836 22615 19839
rect 22738 19836 22744 19848
rect 22603 19808 22744 19836
rect 22603 19805 22615 19808
rect 22557 19799 22615 19805
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 22922 19796 22928 19848
rect 22980 19836 22986 19848
rect 23050 19839 23108 19845
rect 23050 19836 23062 19839
rect 22980 19808 23062 19836
rect 22980 19796 22986 19808
rect 23050 19805 23062 19808
rect 23096 19805 23108 19839
rect 23050 19799 23108 19805
rect 23198 19796 23204 19848
rect 23256 19836 23262 19848
rect 23569 19839 23627 19845
rect 23569 19836 23581 19839
rect 23256 19808 23581 19836
rect 23256 19796 23262 19808
rect 23569 19805 23581 19808
rect 23615 19836 23627 19839
rect 24026 19836 24032 19848
rect 23615 19808 24032 19836
rect 23615 19805 23627 19808
rect 23569 19799 23627 19805
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 25976 19845 26004 19876
rect 27816 19848 27844 19876
rect 29362 19864 29368 19916
rect 29420 19864 29426 19916
rect 29546 19864 29552 19916
rect 29604 19864 29610 19916
rect 30006 19864 30012 19916
rect 30064 19864 30070 19916
rect 30190 19864 30196 19916
rect 30248 19904 30254 19916
rect 33980 19904 34008 19932
rect 34425 19907 34483 19913
rect 34425 19904 34437 19907
rect 30248 19876 31524 19904
rect 30248 19864 30254 19876
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19805 26019 19839
rect 25961 19799 26019 19805
rect 26050 19796 26056 19848
rect 26108 19796 26114 19848
rect 26234 19796 26240 19848
rect 26292 19796 26298 19848
rect 26326 19796 26332 19848
rect 26384 19796 26390 19848
rect 27525 19839 27583 19845
rect 27525 19805 27537 19839
rect 27571 19836 27583 19839
rect 27614 19836 27620 19848
rect 27571 19808 27620 19836
rect 27571 19805 27583 19808
rect 27525 19799 27583 19805
rect 27614 19796 27620 19808
rect 27672 19796 27678 19848
rect 27798 19796 27804 19848
rect 27856 19796 27862 19848
rect 27893 19839 27951 19845
rect 27893 19805 27905 19839
rect 27939 19836 27951 19839
rect 27939 19808 28764 19836
rect 27939 19805 27951 19808
rect 27893 19799 27951 19805
rect 22186 19768 22192 19780
rect 21744 19740 22192 19768
rect 18932 19728 18938 19740
rect 22186 19728 22192 19740
rect 22244 19728 22250 19780
rect 23934 19768 23940 19780
rect 22756 19740 23940 19768
rect 3418 19709 3424 19712
rect 3145 19703 3203 19709
rect 3145 19669 3157 19703
rect 3191 19669 3203 19703
rect 3145 19663 3203 19669
rect 3405 19703 3424 19709
rect 3405 19669 3417 19703
rect 3405 19663 3424 19669
rect 3418 19660 3424 19663
rect 3476 19660 3482 19712
rect 4525 19703 4583 19709
rect 4525 19669 4537 19703
rect 4571 19700 4583 19703
rect 4706 19700 4712 19712
rect 4571 19672 4712 19700
rect 4571 19669 4583 19672
rect 4525 19663 4583 19669
rect 4706 19660 4712 19672
rect 4764 19700 4770 19712
rect 5258 19700 5264 19712
rect 4764 19672 5264 19700
rect 4764 19660 4770 19672
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 7466 19660 7472 19712
rect 7524 19700 7530 19712
rect 8389 19703 8447 19709
rect 8389 19700 8401 19703
rect 7524 19672 8401 19700
rect 7524 19660 7530 19672
rect 8389 19669 8401 19672
rect 8435 19669 8447 19703
rect 8389 19663 8447 19669
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 9953 19703 10011 19709
rect 9953 19700 9965 19703
rect 9824 19672 9965 19700
rect 9824 19660 9830 19672
rect 9953 19669 9965 19672
rect 9999 19669 10011 19703
rect 9953 19663 10011 19669
rect 10318 19660 10324 19712
rect 10376 19660 10382 19712
rect 10413 19703 10471 19709
rect 10413 19669 10425 19703
rect 10459 19700 10471 19703
rect 10781 19703 10839 19709
rect 10781 19700 10793 19703
rect 10459 19672 10793 19700
rect 10459 19669 10471 19672
rect 10413 19663 10471 19669
rect 10781 19669 10793 19672
rect 10827 19700 10839 19703
rect 11882 19700 11888 19712
rect 10827 19672 11888 19700
rect 10827 19669 10839 19672
rect 10781 19663 10839 19669
rect 11882 19660 11888 19672
rect 11940 19700 11946 19712
rect 12434 19700 12440 19712
rect 11940 19672 12440 19700
rect 11940 19660 11946 19672
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19700 13599 19703
rect 13998 19700 14004 19712
rect 13587 19672 14004 19700
rect 13587 19669 13599 19672
rect 13541 19663 13599 19669
rect 13998 19660 14004 19672
rect 14056 19660 14062 19712
rect 14734 19660 14740 19712
rect 14792 19660 14798 19712
rect 18782 19660 18788 19712
rect 18840 19700 18846 19712
rect 21450 19700 21456 19712
rect 18840 19672 21456 19700
rect 18840 19660 18846 19672
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 22097 19703 22155 19709
rect 22097 19669 22109 19703
rect 22143 19700 22155 19703
rect 22756 19700 22784 19740
rect 23934 19728 23940 19740
rect 23992 19728 23998 19780
rect 27706 19728 27712 19780
rect 27764 19728 27770 19780
rect 28736 19777 28764 19808
rect 28810 19796 28816 19848
rect 28868 19796 28874 19848
rect 28994 19796 29000 19848
rect 29052 19836 29058 19848
rect 29089 19839 29147 19845
rect 29089 19836 29101 19839
rect 29052 19808 29101 19836
rect 29052 19796 29058 19808
rect 29089 19805 29101 19808
rect 29135 19836 29147 19839
rect 29638 19836 29644 19848
rect 29135 19808 29644 19836
rect 29135 19805 29147 19808
rect 29089 19799 29147 19805
rect 29638 19796 29644 19808
rect 29696 19796 29702 19848
rect 29730 19796 29736 19848
rect 29788 19796 29794 19848
rect 29822 19796 29828 19848
rect 29880 19836 29886 19848
rect 30377 19839 30435 19845
rect 30377 19836 30389 19839
rect 29880 19808 30389 19836
rect 29880 19796 29886 19808
rect 30377 19805 30389 19808
rect 30423 19805 30435 19839
rect 30377 19799 30435 19805
rect 28721 19771 28779 19777
rect 28721 19737 28733 19771
rect 28767 19768 28779 19771
rect 29454 19768 29460 19780
rect 28767 19740 29460 19768
rect 28767 19737 28779 19740
rect 28721 19731 28779 19737
rect 29454 19728 29460 19740
rect 29512 19728 29518 19780
rect 31202 19728 31208 19780
rect 31260 19728 31266 19780
rect 31496 19768 31524 19876
rect 33796 19876 34437 19904
rect 31570 19796 31576 19848
rect 31628 19836 31634 19848
rect 32582 19845 32588 19848
rect 32401 19839 32459 19845
rect 32401 19836 32413 19839
rect 31628 19808 32413 19836
rect 31628 19796 31634 19808
rect 32401 19805 32413 19808
rect 32447 19805 32459 19839
rect 32579 19836 32588 19845
rect 32543 19808 32588 19836
rect 32401 19799 32459 19805
rect 32579 19799 32588 19808
rect 32582 19796 32588 19799
rect 32640 19796 32646 19848
rect 32674 19796 32680 19848
rect 32732 19836 32738 19848
rect 33796 19845 33824 19876
rect 34425 19873 34437 19876
rect 34471 19873 34483 19907
rect 34425 19867 34483 19873
rect 35986 19864 35992 19916
rect 36044 19864 36050 19916
rect 36280 19848 36308 19944
rect 33796 19839 33869 19845
rect 33796 19836 33823 19839
rect 32732 19808 33823 19836
rect 32732 19796 32738 19808
rect 33796 19805 33823 19808
rect 33857 19805 33869 19839
rect 33796 19802 33869 19805
rect 33811 19799 33869 19802
rect 33965 19839 34023 19845
rect 33965 19805 33977 19839
rect 34011 19836 34023 19839
rect 34146 19836 34152 19848
rect 34011 19808 34152 19836
rect 34011 19805 34023 19808
rect 33965 19799 34023 19805
rect 34146 19796 34152 19808
rect 34204 19796 34210 19848
rect 35894 19796 35900 19848
rect 35952 19836 35958 19848
rect 36173 19839 36231 19845
rect 36173 19836 36185 19839
rect 35952 19808 36185 19836
rect 35952 19796 35958 19808
rect 36173 19805 36185 19808
rect 36219 19805 36231 19839
rect 36173 19799 36231 19805
rect 32122 19768 32128 19780
rect 31496 19740 32128 19768
rect 32122 19728 32128 19740
rect 32180 19728 32186 19780
rect 32306 19728 32312 19780
rect 32364 19768 32370 19780
rect 34057 19771 34115 19777
rect 34057 19768 34069 19771
rect 32364 19740 34069 19768
rect 32364 19728 32370 19740
rect 33796 19712 33824 19740
rect 34057 19737 34069 19740
rect 34103 19737 34115 19771
rect 34057 19731 34115 19737
rect 34241 19771 34299 19777
rect 34241 19737 34253 19771
rect 34287 19768 34299 19771
rect 34330 19768 34336 19780
rect 34287 19740 34336 19768
rect 34287 19737 34299 19740
rect 34241 19731 34299 19737
rect 34330 19728 34336 19740
rect 34388 19728 34394 19780
rect 35989 19771 36047 19777
rect 35989 19737 36001 19771
rect 36035 19768 36047 19771
rect 36078 19768 36084 19780
rect 36035 19740 36084 19768
rect 36035 19737 36047 19740
rect 35989 19731 36047 19737
rect 36078 19728 36084 19740
rect 36136 19728 36142 19780
rect 36188 19768 36216 19799
rect 36262 19796 36268 19848
rect 36320 19796 36326 19848
rect 36372 19845 36400 20012
rect 36446 20000 36452 20052
rect 36504 20000 36510 20052
rect 36722 20000 36728 20052
rect 36780 20040 36786 20052
rect 36909 20043 36967 20049
rect 36909 20040 36921 20043
rect 36780 20012 36921 20040
rect 36780 20000 36786 20012
rect 36909 20009 36921 20012
rect 36955 20009 36967 20043
rect 36909 20003 36967 20009
rect 36538 19864 36544 19916
rect 36596 19904 36602 19916
rect 36633 19907 36691 19913
rect 36633 19904 36645 19907
rect 36596 19876 36645 19904
rect 36596 19864 36602 19876
rect 36633 19873 36645 19876
rect 36679 19904 36691 19907
rect 37918 19904 37924 19916
rect 36679 19876 37924 19904
rect 36679 19873 36691 19876
rect 36633 19867 36691 19873
rect 37918 19864 37924 19876
rect 37976 19864 37982 19916
rect 36357 19839 36415 19845
rect 36357 19805 36369 19839
rect 36403 19805 36415 19839
rect 36357 19799 36415 19805
rect 36446 19768 36452 19780
rect 36188 19740 36452 19768
rect 36446 19728 36452 19740
rect 36504 19728 36510 19780
rect 22143 19672 22784 19700
rect 23109 19703 23167 19709
rect 22143 19669 22155 19672
rect 22097 19663 22155 19669
rect 23109 19669 23121 19703
rect 23155 19700 23167 19703
rect 23198 19700 23204 19712
rect 23155 19672 23204 19700
rect 23155 19669 23167 19672
rect 23109 19663 23167 19669
rect 23198 19660 23204 19672
rect 23256 19660 23262 19712
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 26513 19703 26571 19709
rect 26513 19669 26525 19703
rect 26559 19700 26571 19703
rect 26878 19700 26884 19712
rect 26559 19672 26884 19700
rect 26559 19669 26571 19672
rect 26513 19663 26571 19669
rect 26878 19660 26884 19672
rect 26936 19660 26942 19712
rect 27154 19660 27160 19712
rect 27212 19700 27218 19712
rect 27982 19700 27988 19712
rect 27212 19672 27988 19700
rect 27212 19660 27218 19672
rect 27982 19660 27988 19672
rect 28040 19660 28046 19712
rect 29365 19703 29423 19709
rect 29365 19669 29377 19703
rect 29411 19700 29423 19703
rect 29546 19700 29552 19712
rect 29411 19672 29552 19700
rect 29411 19669 29423 19672
rect 29365 19663 29423 19669
rect 29546 19660 29552 19672
rect 29604 19660 29610 19712
rect 29914 19660 29920 19712
rect 29972 19660 29978 19712
rect 32493 19703 32551 19709
rect 32493 19669 32505 19703
rect 32539 19700 32551 19703
rect 33226 19700 33232 19712
rect 32539 19672 33232 19700
rect 32539 19669 32551 19672
rect 32493 19663 32551 19669
rect 33226 19660 33232 19672
rect 33284 19660 33290 19712
rect 33778 19660 33784 19712
rect 33836 19660 33842 19712
rect 35434 19660 35440 19712
rect 35492 19700 35498 19712
rect 36170 19700 36176 19712
rect 35492 19672 36176 19700
rect 35492 19660 35498 19672
rect 36170 19660 36176 19672
rect 36228 19660 36234 19712
rect 1104 19610 38824 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 38824 19610
rect 1104 19536 38824 19558
rect 21545 19499 21603 19505
rect 21545 19496 21557 19499
rect 2746 19468 21557 19496
rect 106 19388 112 19440
rect 164 19428 170 19440
rect 2746 19428 2774 19468
rect 21545 19465 21557 19468
rect 21591 19496 21603 19499
rect 25869 19499 25927 19505
rect 21591 19468 21864 19496
rect 21591 19465 21603 19468
rect 21545 19459 21603 19465
rect 164 19400 2774 19428
rect 164 19388 170 19400
rect 2866 19388 2872 19440
rect 2924 19428 2930 19440
rect 3697 19431 3755 19437
rect 2924 19400 3648 19428
rect 2924 19388 2930 19400
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 2685 19363 2743 19369
rect 2685 19360 2697 19363
rect 2179 19332 2697 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 2685 19329 2697 19332
rect 2731 19329 2743 19363
rect 3418 19360 3424 19372
rect 2685 19323 2743 19329
rect 3160 19332 3424 19360
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1728 19264 1777 19292
rect 1728 19252 1734 19264
rect 1765 19261 1777 19264
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2225 19295 2283 19301
rect 2225 19261 2237 19295
rect 2271 19292 2283 19295
rect 3160 19292 3188 19332
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 3510 19320 3516 19372
rect 3568 19320 3574 19372
rect 3620 19360 3648 19400
rect 3697 19397 3709 19431
rect 3743 19428 3755 19431
rect 4062 19428 4068 19440
rect 3743 19400 4068 19428
rect 3743 19397 3755 19400
rect 3697 19391 3755 19397
rect 4062 19388 4068 19400
rect 4120 19388 4126 19440
rect 7926 19388 7932 19440
rect 7984 19428 7990 19440
rect 11793 19431 11851 19437
rect 7984 19400 10258 19428
rect 7984 19388 7990 19400
rect 11793 19397 11805 19431
rect 11839 19428 11851 19431
rect 12713 19431 12771 19437
rect 11839 19400 12572 19428
rect 11839 19397 11851 19400
rect 11793 19391 11851 19397
rect 4249 19363 4307 19369
rect 3620 19332 3740 19360
rect 2271 19264 3188 19292
rect 3329 19295 3387 19301
rect 2271 19261 2283 19264
rect 2225 19255 2283 19261
rect 3329 19261 3341 19295
rect 3375 19292 3387 19295
rect 3528 19292 3556 19320
rect 3375 19264 3556 19292
rect 3375 19261 3387 19264
rect 3329 19255 3387 19261
rect 3712 19233 3740 19332
rect 4249 19329 4261 19363
rect 4295 19360 4307 19363
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4295 19332 4721 19360
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 4709 19329 4721 19332
rect 4755 19329 4767 19363
rect 5718 19360 5724 19372
rect 4709 19323 4767 19329
rect 5184 19332 5724 19360
rect 4341 19295 4399 19301
rect 4341 19261 4353 19295
rect 4387 19292 4399 19295
rect 5184 19292 5212 19332
rect 5718 19320 5724 19332
rect 5776 19320 5782 19372
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 7653 19363 7711 19369
rect 7653 19329 7665 19363
rect 7699 19360 7711 19363
rect 8478 19360 8484 19372
rect 7699 19332 8484 19360
rect 7699 19329 7711 19332
rect 7653 19323 7711 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 11882 19320 11888 19372
rect 11940 19320 11946 19372
rect 12250 19320 12256 19372
rect 12308 19320 12314 19372
rect 12544 19334 12572 19400
rect 12713 19397 12725 19431
rect 12759 19428 12771 19431
rect 12986 19428 12992 19440
rect 12759 19400 12992 19428
rect 12759 19397 12771 19400
rect 12713 19391 12771 19397
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 13449 19431 13507 19437
rect 13449 19428 13461 19431
rect 13096 19400 13461 19428
rect 4387 19264 5212 19292
rect 4387 19261 4399 19264
rect 4341 19255 4399 19261
rect 5258 19252 5264 19304
rect 5316 19252 5322 19304
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 9493 19295 9551 19301
rect 9493 19292 9505 19295
rect 9272 19264 9505 19292
rect 9272 19252 9278 19264
rect 9493 19261 9505 19264
rect 9539 19261 9551 19295
rect 9493 19255 9551 19261
rect 9766 19252 9772 19304
rect 9824 19252 9830 19304
rect 10318 19252 10324 19304
rect 10376 19292 10382 19304
rect 10962 19292 10968 19304
rect 10376 19264 10968 19292
rect 10376 19252 10382 19264
rect 10962 19252 10968 19264
rect 11020 19292 11026 19304
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 11020 19264 11253 19292
rect 11020 19252 11026 19264
rect 11241 19261 11253 19264
rect 11287 19261 11299 19295
rect 11241 19255 11299 19261
rect 11609 19295 11667 19301
rect 11609 19261 11621 19295
rect 11655 19261 11667 19295
rect 11609 19255 11667 19261
rect 3697 19227 3755 19233
rect 3697 19193 3709 19227
rect 3743 19193 3755 19227
rect 3697 19187 3755 19193
rect 4617 19227 4675 19233
rect 4617 19193 4629 19227
rect 4663 19224 4675 19227
rect 5994 19224 6000 19236
rect 4663 19196 6000 19224
rect 4663 19193 4675 19196
rect 4617 19187 4675 19193
rect 5994 19184 6000 19196
rect 6052 19184 6058 19236
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 11624 19224 11652 19255
rect 12268 19233 12296 19320
rect 12544 19306 12664 19334
rect 12894 19320 12900 19372
rect 12952 19320 12958 19372
rect 13096 19360 13124 19400
rect 13449 19397 13461 19400
rect 13495 19397 13507 19431
rect 14185 19431 14243 19437
rect 14185 19428 14197 19431
rect 13449 19391 13507 19397
rect 14108 19400 14197 19428
rect 14108 19372 14136 19400
rect 14185 19397 14197 19400
rect 14231 19428 14243 19431
rect 14366 19428 14372 19440
rect 14231 19400 14372 19428
rect 14231 19397 14243 19400
rect 14185 19391 14243 19397
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 18782 19388 18788 19440
rect 18840 19388 18846 19440
rect 20806 19388 20812 19440
rect 20864 19388 20870 19440
rect 21836 19437 21864 19468
rect 25869 19465 25881 19499
rect 25915 19496 25927 19499
rect 26050 19496 26056 19508
rect 25915 19468 26056 19496
rect 25915 19465 25927 19468
rect 25869 19459 25927 19465
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 27062 19456 27068 19508
rect 27120 19496 27126 19508
rect 28445 19499 28503 19505
rect 27120 19468 28120 19496
rect 27120 19456 27126 19468
rect 21821 19431 21879 19437
rect 21821 19397 21833 19431
rect 21867 19397 21879 19431
rect 21821 19391 21879 19397
rect 22922 19388 22928 19440
rect 22980 19428 22986 19440
rect 22980 19400 23888 19428
rect 22980 19388 22986 19400
rect 13004 19332 13124 19360
rect 12636 19292 12664 19306
rect 13004 19292 13032 19332
rect 13170 19320 13176 19372
rect 13228 19320 13234 19372
rect 13357 19363 13415 19369
rect 13357 19329 13369 19363
rect 13403 19360 13415 19363
rect 13998 19360 14004 19372
rect 13403 19332 14004 19360
rect 13403 19329 13415 19332
rect 13357 19323 13415 19329
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 14090 19320 14096 19372
rect 14148 19320 14154 19372
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 12636 19264 13032 19292
rect 13446 19252 13452 19304
rect 13504 19292 13510 19304
rect 14277 19295 14335 19301
rect 14277 19292 14289 19295
rect 13504 19264 14289 19292
rect 13504 19252 13510 19264
rect 14277 19261 14289 19264
rect 14323 19261 14335 19295
rect 14277 19255 14335 19261
rect 10836 19196 11652 19224
rect 12253 19227 12311 19233
rect 10836 19184 10842 19196
rect 12253 19193 12265 19227
rect 12299 19193 12311 19227
rect 12253 19187 12311 19193
rect 12434 19184 12440 19236
rect 12492 19224 12498 19236
rect 13464 19224 13492 19252
rect 12492 19196 13492 19224
rect 12492 19184 12498 19196
rect 13998 19184 14004 19236
rect 14056 19224 14062 19236
rect 14476 19224 14504 19323
rect 14734 19320 14740 19372
rect 14792 19320 14798 19372
rect 16114 19320 16120 19372
rect 16172 19320 16178 19372
rect 16574 19360 16580 19372
rect 16500 19332 16580 19360
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15470 19292 15476 19304
rect 15059 19264 15476 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 16500 19301 16528 19332
rect 16574 19320 16580 19332
rect 16632 19320 16638 19372
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 18506 19320 18512 19372
rect 18564 19320 18570 19372
rect 18690 19320 18696 19372
rect 18748 19320 18754 19372
rect 18874 19320 18880 19372
rect 18932 19320 18938 19372
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 18984 19332 19533 19360
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18984 19292 19012 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 23014 19320 23020 19372
rect 23072 19360 23078 19372
rect 23860 19369 23888 19400
rect 24210 19388 24216 19440
rect 24268 19428 24274 19440
rect 24305 19431 24363 19437
rect 24305 19428 24317 19431
rect 24268 19400 24317 19428
rect 24268 19388 24274 19400
rect 24305 19397 24317 19400
rect 24351 19397 24363 19431
rect 25225 19431 25283 19437
rect 25225 19428 25237 19431
rect 24305 19391 24363 19397
rect 24688 19400 25237 19428
rect 23661 19363 23719 19369
rect 23661 19360 23673 19363
rect 23072 19332 23673 19360
rect 23072 19320 23078 19332
rect 23661 19329 23673 19332
rect 23707 19329 23719 19363
rect 23661 19323 23719 19329
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 23934 19320 23940 19372
rect 23992 19320 23998 19372
rect 24026 19320 24032 19372
rect 24084 19320 24090 19372
rect 24688 19369 24716 19400
rect 25225 19397 25237 19400
rect 25271 19397 25283 19431
rect 25225 19391 25283 19397
rect 26786 19388 26792 19440
rect 26844 19428 26850 19440
rect 28092 19437 28120 19468
rect 28445 19465 28457 19499
rect 28491 19496 28503 19499
rect 28994 19496 29000 19508
rect 28491 19468 29000 19496
rect 28491 19465 28503 19468
rect 28445 19459 28503 19465
rect 28994 19456 29000 19468
rect 29052 19456 29058 19508
rect 31754 19496 31760 19508
rect 29288 19468 31760 19496
rect 28077 19431 28135 19437
rect 26844 19400 27844 19428
rect 26844 19388 26850 19400
rect 24673 19363 24731 19369
rect 24673 19329 24685 19363
rect 24719 19329 24731 19363
rect 24673 19323 24731 19329
rect 25133 19363 25191 19369
rect 25133 19329 25145 19363
rect 25179 19329 25191 19363
rect 25133 19323 25191 19329
rect 18012 19264 19012 19292
rect 18012 19252 18018 19264
rect 19794 19252 19800 19304
rect 19852 19252 19858 19304
rect 24765 19295 24823 19301
rect 24765 19261 24777 19295
rect 24811 19292 24823 19295
rect 24854 19292 24860 19304
rect 24811 19264 24860 19292
rect 24811 19261 24823 19264
rect 24765 19255 24823 19261
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 25148 19292 25176 19323
rect 25314 19320 25320 19372
rect 25372 19320 25378 19372
rect 25774 19320 25780 19372
rect 25832 19320 25838 19372
rect 25958 19320 25964 19372
rect 26016 19320 26022 19372
rect 26694 19320 26700 19372
rect 26752 19360 26758 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26752 19332 26985 19360
rect 26752 19320 26758 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 25406 19292 25412 19304
rect 25148 19264 25412 19292
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 14056 19196 14504 19224
rect 25041 19227 25099 19233
rect 14056 19184 14062 19196
rect 25041 19193 25053 19227
rect 25087 19224 25099 19227
rect 26326 19224 26332 19236
rect 25087 19196 26332 19224
rect 25087 19193 25099 19196
rect 25041 19187 25099 19193
rect 26326 19184 26332 19196
rect 26384 19184 26390 19236
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 7653 19159 7711 19165
rect 7653 19156 7665 19159
rect 6972 19128 7665 19156
rect 6972 19116 6978 19128
rect 7653 19125 7665 19128
rect 7699 19125 7711 19159
rect 7653 19119 7711 19125
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 14185 19159 14243 19165
rect 14185 19156 14197 19159
rect 13412 19128 14197 19156
rect 13412 19116 13418 19128
rect 14185 19125 14197 19128
rect 14231 19125 14243 19159
rect 14185 19119 14243 19125
rect 14645 19159 14703 19165
rect 14645 19125 14657 19159
rect 14691 19156 14703 19159
rect 15010 19156 15016 19168
rect 14691 19128 15016 19156
rect 14691 19125 14703 19128
rect 14645 19119 14703 19125
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 16853 19159 16911 19165
rect 16853 19125 16865 19159
rect 16899 19156 16911 19159
rect 17034 19156 17040 19168
rect 16899 19128 17040 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 19061 19159 19119 19165
rect 19061 19125 19073 19159
rect 19107 19156 19119 19159
rect 19334 19156 19340 19168
rect 19107 19128 19340 19156
rect 19107 19125 19119 19128
rect 19061 19119 19119 19125
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 21266 19116 21272 19168
rect 21324 19116 21330 19168
rect 23106 19116 23112 19168
rect 23164 19156 23170 19168
rect 23658 19156 23664 19168
rect 23164 19128 23664 19156
rect 23164 19116 23170 19128
rect 23658 19116 23664 19128
rect 23716 19116 23722 19168
rect 26988 19156 27016 19323
rect 27154 19320 27160 19372
rect 27212 19320 27218 19372
rect 27522 19320 27528 19372
rect 27580 19320 27586 19372
rect 27816 19369 27844 19400
rect 28077 19397 28089 19431
rect 28123 19397 28135 19431
rect 28077 19391 28135 19397
rect 28166 19388 28172 19440
rect 28224 19388 28230 19440
rect 29288 19437 29316 19468
rect 31754 19456 31760 19468
rect 31812 19456 31818 19508
rect 32122 19456 32128 19508
rect 32180 19496 32186 19508
rect 32180 19468 32536 19496
rect 32180 19456 32186 19468
rect 29273 19431 29331 19437
rect 29273 19397 29285 19431
rect 29319 19397 29331 19431
rect 29273 19391 29331 19397
rect 29365 19431 29423 19437
rect 29365 19397 29377 19431
rect 29411 19428 29423 19431
rect 29638 19428 29644 19440
rect 29411 19400 29644 19428
rect 29411 19397 29423 19400
rect 29365 19391 29423 19397
rect 29638 19388 29644 19400
rect 29696 19388 29702 19440
rect 29914 19388 29920 19440
rect 29972 19388 29978 19440
rect 30098 19388 30104 19440
rect 30156 19388 30162 19440
rect 31570 19388 31576 19440
rect 31628 19428 31634 19440
rect 32508 19437 32536 19468
rect 32582 19456 32588 19508
rect 32640 19496 32646 19508
rect 33318 19496 33324 19508
rect 32640 19468 33324 19496
rect 32640 19456 32646 19468
rect 33318 19456 33324 19468
rect 33376 19456 33382 19508
rect 33413 19499 33471 19505
rect 33413 19465 33425 19499
rect 33459 19496 33471 19499
rect 33594 19496 33600 19508
rect 33459 19468 33600 19496
rect 33459 19465 33471 19468
rect 33413 19459 33471 19465
rect 33594 19456 33600 19468
rect 33652 19496 33658 19508
rect 33965 19499 34023 19505
rect 33965 19496 33977 19499
rect 33652 19468 33977 19496
rect 33652 19456 33658 19468
rect 33965 19465 33977 19468
rect 34011 19496 34023 19499
rect 34146 19496 34152 19508
rect 34011 19468 34152 19496
rect 34011 19465 34023 19468
rect 33965 19459 34023 19465
rect 34146 19456 34152 19468
rect 34204 19456 34210 19508
rect 35434 19456 35440 19508
rect 35492 19496 35498 19508
rect 35621 19499 35679 19505
rect 35621 19496 35633 19499
rect 35492 19468 35633 19496
rect 35492 19456 35498 19468
rect 35621 19465 35633 19468
rect 35667 19465 35679 19499
rect 35621 19459 35679 19465
rect 35710 19456 35716 19508
rect 35768 19496 35774 19508
rect 36262 19496 36268 19508
rect 35768 19468 36268 19496
rect 35768 19456 35774 19468
rect 36262 19456 36268 19468
rect 36320 19496 36326 19508
rect 36357 19499 36415 19505
rect 36357 19496 36369 19499
rect 36320 19468 36369 19496
rect 36320 19456 36326 19468
rect 36357 19465 36369 19468
rect 36403 19465 36415 19499
rect 36357 19459 36415 19465
rect 36630 19456 36636 19508
rect 36688 19496 36694 19508
rect 36817 19499 36875 19505
rect 36817 19496 36829 19499
rect 36688 19468 36829 19496
rect 36688 19456 36694 19468
rect 36817 19465 36829 19468
rect 36863 19465 36875 19499
rect 36817 19459 36875 19465
rect 31665 19431 31723 19437
rect 31665 19428 31677 19431
rect 31628 19400 31677 19428
rect 31628 19388 31634 19400
rect 31665 19397 31677 19400
rect 31711 19397 31723 19431
rect 31665 19391 31723 19397
rect 31849 19431 31907 19437
rect 31849 19397 31861 19431
rect 31895 19428 31907 19431
rect 32217 19431 32275 19437
rect 32217 19428 32229 19431
rect 31895 19400 32229 19428
rect 31895 19397 31907 19400
rect 31849 19391 31907 19397
rect 32217 19397 32229 19400
rect 32263 19397 32275 19431
rect 32217 19391 32275 19397
rect 32493 19431 32551 19437
rect 32493 19397 32505 19431
rect 32539 19397 32551 19431
rect 32493 19391 32551 19397
rect 32674 19388 32680 19440
rect 32732 19388 32738 19440
rect 33336 19428 33364 19456
rect 35805 19431 35863 19437
rect 35805 19428 35817 19431
rect 33336 19400 33640 19428
rect 27801 19363 27859 19369
rect 27801 19329 27813 19363
rect 27847 19329 27859 19363
rect 27801 19323 27859 19329
rect 27890 19320 27896 19372
rect 27948 19360 27954 19372
rect 28307 19363 28365 19369
rect 27948 19332 27993 19360
rect 27948 19320 27954 19332
rect 28307 19329 28319 19363
rect 28353 19360 28365 19363
rect 28353 19332 29040 19360
rect 28353 19329 28365 19332
rect 28307 19323 28365 19329
rect 27062 19252 27068 19304
rect 27120 19292 27126 19304
rect 27249 19295 27307 19301
rect 27249 19292 27261 19295
rect 27120 19264 27261 19292
rect 27120 19252 27126 19264
rect 27249 19261 27261 19264
rect 27295 19261 27307 19295
rect 27249 19255 27307 19261
rect 27341 19295 27399 19301
rect 27341 19261 27353 19295
rect 27387 19261 27399 19295
rect 27341 19255 27399 19261
rect 27356 19224 27384 19255
rect 27614 19252 27620 19304
rect 27672 19292 27678 19304
rect 27709 19295 27767 19301
rect 27709 19292 27721 19295
rect 27672 19264 27721 19292
rect 27672 19252 27678 19264
rect 27709 19261 27721 19264
rect 27755 19261 27767 19295
rect 29012 19292 29040 19332
rect 29086 19320 29092 19372
rect 29144 19320 29150 19372
rect 29454 19320 29460 19372
rect 29512 19320 29518 19372
rect 29822 19360 29828 19372
rect 29656 19332 29828 19360
rect 29270 19292 29276 19304
rect 29012 19264 29276 19292
rect 27709 19255 27767 19261
rect 29270 19252 29276 19264
rect 29328 19252 29334 19304
rect 28074 19224 28080 19236
rect 27356 19196 28080 19224
rect 28074 19184 28080 19196
rect 28132 19184 28138 19236
rect 29656 19233 29684 19332
rect 29822 19320 29828 19332
rect 29880 19320 29886 19372
rect 30116 19360 30144 19388
rect 32125 19363 32183 19369
rect 32125 19360 32137 19363
rect 30116 19332 32137 19360
rect 32125 19329 32137 19332
rect 32171 19360 32183 19363
rect 32171 19332 32260 19360
rect 32171 19329 32183 19332
rect 32125 19323 32183 19329
rect 32232 19292 32260 19332
rect 32306 19320 32312 19372
rect 32364 19320 32370 19372
rect 32416 19332 33180 19360
rect 32416 19292 32444 19332
rect 32232 19264 32444 19292
rect 33152 19292 33180 19332
rect 33226 19320 33232 19372
rect 33284 19320 33290 19372
rect 33502 19320 33508 19372
rect 33560 19320 33566 19372
rect 33520 19292 33548 19320
rect 33612 19301 33640 19400
rect 35544 19400 35817 19428
rect 33778 19320 33784 19372
rect 33836 19320 33842 19372
rect 34609 19363 34667 19369
rect 34609 19329 34621 19363
rect 34655 19360 34667 19363
rect 34790 19360 34796 19372
rect 34655 19332 34796 19360
rect 34655 19329 34667 19332
rect 34609 19323 34667 19329
rect 34790 19320 34796 19332
rect 34848 19320 34854 19372
rect 35544 19369 35572 19400
rect 35805 19397 35817 19400
rect 35851 19397 35863 19431
rect 35805 19391 35863 19397
rect 36078 19388 36084 19440
rect 36136 19428 36142 19440
rect 36173 19431 36231 19437
rect 36173 19428 36185 19431
rect 36136 19400 36185 19428
rect 36136 19388 36142 19400
rect 36173 19397 36185 19400
rect 36219 19428 36231 19431
rect 36906 19428 36912 19440
rect 36219 19400 36912 19428
rect 36219 19397 36231 19400
rect 36173 19391 36231 19397
rect 36906 19388 36912 19400
rect 36964 19388 36970 19440
rect 35529 19363 35587 19369
rect 35529 19329 35541 19363
rect 35575 19329 35587 19363
rect 35529 19323 35587 19329
rect 35713 19363 35771 19369
rect 35713 19329 35725 19363
rect 35759 19329 35771 19363
rect 35713 19323 35771 19329
rect 33152 19264 33548 19292
rect 33597 19295 33655 19301
rect 33597 19261 33609 19295
rect 33643 19292 33655 19295
rect 34330 19292 34336 19304
rect 33643 19264 34336 19292
rect 33643 19261 33655 19264
rect 33597 19255 33655 19261
rect 34330 19252 34336 19264
rect 34388 19252 34394 19304
rect 29641 19227 29699 19233
rect 29641 19193 29653 19227
rect 29687 19193 29699 19227
rect 29641 19187 29699 19193
rect 33134 19184 33140 19236
rect 33192 19224 33198 19236
rect 35728 19224 35756 19323
rect 35986 19320 35992 19372
rect 36044 19320 36050 19372
rect 36262 19320 36268 19372
rect 36320 19320 36326 19372
rect 36354 19320 36360 19372
rect 36412 19360 36418 19372
rect 36541 19363 36599 19369
rect 36541 19360 36553 19363
rect 36412 19332 36553 19360
rect 36412 19320 36418 19332
rect 36541 19329 36553 19332
rect 36587 19329 36599 19363
rect 36541 19323 36599 19329
rect 36814 19320 36820 19372
rect 36872 19320 36878 19372
rect 36998 19320 37004 19372
rect 37056 19360 37062 19372
rect 37093 19363 37151 19369
rect 37093 19360 37105 19363
rect 37056 19332 37105 19360
rect 37056 19320 37062 19332
rect 37093 19329 37105 19332
rect 37139 19329 37151 19363
rect 37093 19323 37151 19329
rect 36725 19295 36783 19301
rect 36725 19261 36737 19295
rect 36771 19292 36783 19295
rect 37366 19292 37372 19304
rect 36771 19264 37372 19292
rect 36771 19261 36783 19264
rect 36725 19255 36783 19261
rect 37366 19252 37372 19264
rect 37424 19292 37430 19304
rect 38378 19292 38384 19304
rect 37424 19264 38384 19292
rect 37424 19252 37430 19264
rect 38378 19252 38384 19264
rect 38436 19252 38442 19304
rect 36630 19224 36636 19236
rect 33192 19196 35664 19224
rect 35728 19196 36636 19224
rect 33192 19184 33198 19196
rect 27798 19156 27804 19168
rect 26988 19128 27804 19156
rect 27798 19116 27804 19128
rect 27856 19156 27862 19168
rect 28810 19156 28816 19168
rect 27856 19128 28816 19156
rect 27856 19116 27862 19128
rect 28810 19116 28816 19128
rect 28868 19116 28874 19168
rect 29178 19116 29184 19168
rect 29236 19156 29242 19168
rect 30285 19159 30343 19165
rect 30285 19156 30297 19159
rect 29236 19128 30297 19156
rect 29236 19116 29242 19128
rect 30285 19125 30297 19128
rect 30331 19125 30343 19159
rect 30285 19119 30343 19125
rect 31386 19116 31392 19168
rect 31444 19156 31450 19168
rect 31481 19159 31539 19165
rect 31481 19156 31493 19159
rect 31444 19128 31493 19156
rect 31444 19116 31450 19128
rect 31481 19125 31493 19128
rect 31527 19125 31539 19159
rect 31481 19119 31539 19125
rect 32766 19116 32772 19168
rect 32824 19116 32830 19168
rect 33042 19116 33048 19168
rect 33100 19156 33106 19168
rect 34146 19156 34152 19168
rect 33100 19128 34152 19156
rect 33100 19116 33106 19128
rect 34146 19116 34152 19128
rect 34204 19116 34210 19168
rect 34698 19116 34704 19168
rect 34756 19156 34762 19168
rect 34793 19159 34851 19165
rect 34793 19156 34805 19159
rect 34756 19128 34805 19156
rect 34756 19116 34762 19128
rect 34793 19125 34805 19128
rect 34839 19125 34851 19159
rect 35636 19156 35664 19196
rect 36630 19184 36636 19196
rect 36688 19184 36694 19236
rect 36170 19156 36176 19168
rect 35636 19128 36176 19156
rect 34793 19119 34851 19125
rect 36170 19116 36176 19128
rect 36228 19156 36234 19168
rect 36998 19156 37004 19168
rect 36228 19128 37004 19156
rect 36228 19116 36234 19128
rect 36998 19116 37004 19128
rect 37056 19116 37062 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 3510 18952 3516 18964
rect 3467 18924 3516 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 3970 18952 3976 18964
rect 3927 18924 3976 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 4157 18955 4215 18961
rect 4157 18921 4169 18955
rect 4203 18952 4215 18955
rect 4617 18955 4675 18961
rect 4203 18924 4568 18952
rect 4203 18921 4215 18924
rect 4157 18915 4215 18921
rect 3528 18816 3556 18912
rect 4540 18896 4568 18924
rect 4617 18921 4629 18955
rect 4663 18921 4675 18955
rect 4617 18915 4675 18921
rect 3605 18887 3663 18893
rect 3605 18853 3617 18887
rect 3651 18884 3663 18887
rect 4249 18887 4307 18893
rect 4249 18884 4261 18887
rect 3651 18856 4261 18884
rect 3651 18853 3663 18856
rect 3605 18847 3663 18853
rect 4249 18853 4261 18856
rect 4295 18853 4307 18887
rect 4249 18847 4307 18853
rect 4522 18844 4528 18896
rect 4580 18844 4586 18896
rect 4632 18816 4660 18915
rect 8478 18912 8484 18964
rect 8536 18912 8542 18964
rect 13081 18955 13139 18961
rect 13081 18921 13093 18955
rect 13127 18952 13139 18955
rect 13170 18952 13176 18964
rect 13127 18924 13176 18952
rect 13127 18921 13139 18924
rect 13081 18915 13139 18921
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 14642 18912 14648 18964
rect 14700 18912 14706 18964
rect 15838 18912 15844 18964
rect 15896 18952 15902 18964
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 15896 18924 16129 18952
rect 15896 18912 15902 18924
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16117 18915 16175 18921
rect 17037 18955 17095 18961
rect 17037 18921 17049 18955
rect 17083 18952 17095 18955
rect 17126 18952 17132 18964
rect 17083 18924 17132 18952
rect 17083 18921 17095 18924
rect 17037 18915 17095 18921
rect 17126 18912 17132 18924
rect 17184 18952 17190 18964
rect 17402 18952 17408 18964
rect 17184 18924 17408 18952
rect 17184 18912 17190 18924
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 23569 18955 23627 18961
rect 23569 18921 23581 18955
rect 23615 18952 23627 18955
rect 23934 18952 23940 18964
rect 23615 18924 23940 18952
rect 23615 18921 23627 18924
rect 23569 18915 23627 18921
rect 23934 18912 23940 18924
rect 23992 18912 23998 18964
rect 25133 18955 25191 18961
rect 25133 18921 25145 18955
rect 25179 18952 25191 18955
rect 25774 18952 25780 18964
rect 25179 18924 25780 18952
rect 25179 18921 25191 18924
rect 25133 18915 25191 18921
rect 25774 18912 25780 18924
rect 25832 18912 25838 18964
rect 27433 18955 27491 18961
rect 27433 18921 27445 18955
rect 27479 18952 27491 18955
rect 27706 18952 27712 18964
rect 27479 18924 27712 18952
rect 27479 18921 27491 18924
rect 27433 18915 27491 18921
rect 27706 18912 27712 18924
rect 27764 18912 27770 18964
rect 28721 18955 28779 18961
rect 28721 18921 28733 18955
rect 28767 18952 28779 18955
rect 29086 18952 29092 18964
rect 28767 18924 29092 18952
rect 28767 18921 28779 18924
rect 28721 18915 28779 18921
rect 29086 18912 29092 18924
rect 29144 18912 29150 18964
rect 33502 18952 33508 18964
rect 33336 18924 33508 18952
rect 10962 18844 10968 18896
rect 11020 18884 11026 18896
rect 13354 18884 13360 18896
rect 11020 18856 13360 18884
rect 11020 18844 11026 18856
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 15856 18884 15884 18912
rect 15764 18856 15884 18884
rect 17221 18887 17279 18893
rect 3528 18788 4660 18816
rect 6914 18776 6920 18828
rect 6972 18776 6978 18828
rect 13173 18819 13231 18825
rect 13173 18816 13185 18819
rect 12636 18788 13185 18816
rect 3234 18708 3240 18760
rect 3292 18708 3298 18760
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 3436 18680 3464 18711
rect 3694 18708 3700 18760
rect 3752 18748 3758 18760
rect 3970 18748 3976 18760
rect 3752 18720 3976 18748
rect 3752 18708 3758 18720
rect 3970 18708 3976 18720
rect 4028 18748 4034 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 4028 18720 4077 18748
rect 4028 18708 4034 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 4338 18708 4344 18760
rect 4396 18708 4402 18760
rect 4522 18708 4528 18760
rect 4580 18748 4586 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 4580 18720 4629 18748
rect 4580 18708 4586 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 4724 18680 4752 18708
rect 3436 18652 4752 18680
rect 6656 18680 6684 18711
rect 8018 18708 8024 18760
rect 8076 18708 8082 18760
rect 8478 18708 8484 18760
rect 8536 18708 8542 18760
rect 8662 18708 8668 18760
rect 8720 18708 8726 18760
rect 9122 18708 9128 18760
rect 9180 18708 9186 18760
rect 12434 18708 12440 18760
rect 12492 18708 12498 18760
rect 12636 18757 12664 18788
rect 13173 18785 13185 18788
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 13998 18776 14004 18828
rect 14056 18816 14062 18828
rect 14056 18788 14320 18816
rect 14056 18776 14062 18788
rect 14292 18760 14320 18788
rect 12621 18751 12679 18757
rect 12621 18717 12633 18751
rect 12667 18717 12679 18751
rect 12621 18711 12679 18717
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 6822 18680 6828 18692
rect 6656 18652 6828 18680
rect 6822 18640 6828 18652
rect 6880 18640 6886 18692
rect 9398 18640 9404 18692
rect 9456 18640 9462 18692
rect 10410 18640 10416 18692
rect 10468 18640 10474 18692
rect 12912 18680 12940 18711
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 13630 18708 13636 18760
rect 13688 18708 13694 18760
rect 13817 18751 13875 18757
rect 13817 18717 13829 18751
rect 13863 18748 13875 18751
rect 13906 18748 13912 18760
rect 13863 18720 13912 18748
rect 13863 18717 13875 18720
rect 13817 18711 13875 18717
rect 13906 18708 13912 18720
rect 13964 18708 13970 18760
rect 14090 18708 14096 18760
rect 14148 18708 14154 18760
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 15194 18708 15200 18760
rect 15252 18708 15258 18760
rect 15657 18751 15715 18757
rect 15657 18717 15669 18751
rect 15703 18748 15715 18751
rect 15764 18748 15792 18856
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 18690 18884 18696 18896
rect 17267 18856 18696 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 25593 18887 25651 18893
rect 25593 18853 25605 18887
rect 25639 18884 25651 18887
rect 27062 18884 27068 18896
rect 25639 18856 27068 18884
rect 25639 18853 25651 18856
rect 25593 18847 25651 18853
rect 27062 18844 27068 18856
rect 27120 18844 27126 18896
rect 31754 18844 31760 18896
rect 31812 18884 31818 18896
rect 32490 18884 32496 18896
rect 31812 18856 32496 18884
rect 31812 18844 31818 18856
rect 32490 18844 32496 18856
rect 32548 18844 32554 18896
rect 15930 18776 15936 18828
rect 15988 18776 15994 18828
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17586 18816 17592 18828
rect 16816 18788 17592 18816
rect 16816 18776 16822 18788
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 18874 18816 18880 18828
rect 17696 18788 18880 18816
rect 15703 18720 15792 18748
rect 15703 18717 15715 18720
rect 15657 18711 15715 18717
rect 16022 18708 16028 18760
rect 16080 18748 16086 18760
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 16080 18720 17325 18748
rect 16080 18708 16086 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17696 18757 17724 18788
rect 18874 18776 18880 18788
rect 18932 18776 18938 18828
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 19392 18788 19717 18816
rect 19392 18776 19398 18788
rect 19705 18785 19717 18788
rect 19751 18785 19763 18819
rect 22002 18816 22008 18828
rect 19705 18779 19763 18785
rect 20824 18788 22008 18816
rect 20824 18760 20852 18788
rect 22002 18776 22008 18788
rect 22060 18776 22066 18828
rect 22373 18819 22431 18825
rect 22373 18785 22385 18819
rect 22419 18816 22431 18819
rect 22462 18816 22468 18828
rect 22419 18788 22468 18816
rect 22419 18785 22431 18788
rect 22373 18779 22431 18785
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 23293 18819 23351 18825
rect 23293 18785 23305 18819
rect 23339 18816 23351 18819
rect 23382 18816 23388 18828
rect 23339 18788 23388 18816
rect 23339 18785 23351 18788
rect 23293 18779 23351 18785
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 25501 18819 25559 18825
rect 25501 18816 25513 18819
rect 24872 18788 25513 18816
rect 24872 18760 24900 18788
rect 25501 18785 25513 18788
rect 25547 18785 25559 18819
rect 25501 18779 25559 18785
rect 25685 18819 25743 18825
rect 25685 18785 25697 18819
rect 25731 18816 25743 18819
rect 25958 18816 25964 18828
rect 25731 18788 25964 18816
rect 25731 18785 25743 18788
rect 25685 18779 25743 18785
rect 25958 18776 25964 18788
rect 26016 18816 26022 18828
rect 26016 18788 27016 18816
rect 26016 18776 26022 18788
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 17460 18720 17509 18748
rect 17460 18708 17466 18720
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 17681 18751 17739 18757
rect 17681 18717 17693 18751
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18472 18720 18521 18748
rect 18472 18708 18478 18720
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 14108 18680 14136 18708
rect 12912 18652 14136 18680
rect 15105 18683 15163 18689
rect 15105 18649 15117 18683
rect 15151 18680 15163 18683
rect 16298 18680 16304 18692
rect 15151 18652 16304 18680
rect 15151 18649 15163 18652
rect 15105 18643 15163 18649
rect 16298 18640 16304 18652
rect 16356 18680 16362 18692
rect 16853 18683 16911 18689
rect 16853 18680 16865 18683
rect 16356 18652 16865 18680
rect 16356 18640 16362 18652
rect 16853 18649 16865 18652
rect 16899 18649 16911 18683
rect 16853 18643 16911 18649
rect 17034 18640 17040 18692
rect 17092 18689 17098 18692
rect 17092 18683 17111 18689
rect 17099 18649 17111 18683
rect 17092 18643 17111 18649
rect 17092 18640 17098 18643
rect 17586 18640 17592 18692
rect 17644 18640 17650 18692
rect 17770 18640 17776 18692
rect 17828 18680 17834 18692
rect 17957 18683 18015 18689
rect 17957 18680 17969 18683
rect 17828 18652 17969 18680
rect 17828 18640 17834 18652
rect 17957 18649 17969 18652
rect 18003 18649 18015 18683
rect 17957 18643 18015 18649
rect 4433 18615 4491 18621
rect 4433 18581 4445 18615
rect 4479 18612 4491 18615
rect 4614 18612 4620 18624
rect 4479 18584 4620 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 4614 18572 4620 18584
rect 4672 18572 4678 18624
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 4985 18615 5043 18621
rect 4985 18612 4997 18615
rect 4856 18584 4997 18612
rect 4856 18572 4862 18584
rect 4985 18581 4997 18584
rect 5031 18581 5043 18615
rect 4985 18575 5043 18581
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8389 18615 8447 18621
rect 8389 18612 8401 18615
rect 8352 18584 8401 18612
rect 8352 18572 8358 18584
rect 8389 18581 8401 18584
rect 8435 18581 8447 18615
rect 8389 18575 8447 18581
rect 10870 18572 10876 18624
rect 10928 18572 10934 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 13320 18584 14197 18612
rect 13320 18572 13326 18584
rect 14185 18581 14197 18584
rect 14231 18581 14243 18615
rect 14185 18575 14243 18581
rect 15286 18572 15292 18624
rect 15344 18572 15350 18624
rect 15746 18572 15752 18624
rect 15804 18572 15810 18624
rect 17862 18572 17868 18624
rect 17920 18572 17926 18624
rect 18524 18612 18552 18711
rect 19426 18708 19432 18760
rect 19484 18708 19490 18760
rect 20806 18708 20812 18760
rect 20864 18708 20870 18760
rect 21266 18708 21272 18760
rect 21324 18748 21330 18760
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 21324 18720 21557 18748
rect 21324 18708 21330 18720
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 21726 18708 21732 18760
rect 21784 18708 21790 18760
rect 21910 18748 21916 18760
rect 21836 18720 21916 18748
rect 21450 18640 21456 18692
rect 21508 18680 21514 18692
rect 21836 18680 21864 18720
rect 21910 18708 21916 18720
rect 21968 18748 21974 18760
rect 22097 18751 22155 18757
rect 22097 18748 22109 18751
rect 21968 18720 22109 18748
rect 21968 18708 21974 18720
rect 22097 18717 22109 18720
rect 22143 18717 22155 18751
rect 22097 18711 22155 18717
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 21508 18652 21864 18680
rect 22005 18683 22063 18689
rect 21508 18640 21514 18652
rect 22005 18649 22017 18683
rect 22051 18680 22063 18683
rect 22572 18680 22600 18711
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22796 18720 23029 18748
rect 22796 18708 22802 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 23198 18708 23204 18760
rect 23256 18748 23262 18760
rect 23845 18751 23903 18757
rect 23845 18748 23857 18751
rect 23256 18720 23857 18748
rect 23256 18708 23262 18720
rect 23216 18680 23244 18708
rect 23584 18689 23612 18720
rect 23845 18717 23857 18720
rect 23891 18717 23903 18751
rect 23845 18711 23903 18717
rect 23934 18708 23940 18760
rect 23992 18748 23998 18760
rect 24029 18751 24087 18757
rect 24029 18748 24041 18751
rect 23992 18720 24041 18748
rect 23992 18708 23998 18720
rect 24029 18717 24041 18720
rect 24075 18717 24087 18751
rect 24029 18711 24087 18717
rect 24118 18708 24124 18760
rect 24176 18708 24182 18760
rect 24854 18708 24860 18760
rect 24912 18708 24918 18760
rect 25314 18708 25320 18760
rect 25372 18708 25378 18760
rect 25406 18708 25412 18760
rect 25464 18708 25470 18760
rect 26878 18708 26884 18760
rect 26936 18708 26942 18760
rect 22051 18652 23244 18680
rect 23385 18683 23443 18689
rect 22051 18649 22063 18652
rect 22005 18643 22063 18649
rect 23385 18649 23397 18683
rect 23431 18649 23443 18683
rect 23584 18683 23643 18689
rect 23584 18652 23597 18683
rect 23385 18643 23443 18649
rect 23585 18649 23597 18652
rect 23631 18649 23643 18683
rect 24136 18680 24164 18708
rect 23585 18643 23643 18649
rect 23676 18652 24164 18680
rect 24949 18683 25007 18689
rect 21726 18612 21732 18624
rect 18524 18584 21732 18612
rect 21726 18572 21732 18584
rect 21784 18572 21790 18624
rect 23400 18612 23428 18643
rect 23676 18612 23704 18652
rect 24949 18649 24961 18683
rect 24995 18680 25007 18683
rect 25424 18680 25452 18708
rect 26988 18692 27016 18788
rect 27246 18776 27252 18828
rect 27304 18776 27310 18828
rect 27798 18776 27804 18828
rect 27856 18816 27862 18828
rect 28353 18819 28411 18825
rect 27856 18788 28028 18816
rect 27856 18776 27862 18788
rect 27065 18751 27123 18757
rect 27065 18717 27077 18751
rect 27111 18748 27123 18751
rect 27264 18748 27292 18776
rect 27111 18720 27292 18748
rect 27111 18717 27123 18720
rect 27065 18711 27123 18717
rect 27338 18708 27344 18760
rect 27396 18708 27402 18760
rect 27617 18751 27675 18757
rect 27617 18717 27629 18751
rect 27663 18748 27675 18751
rect 27890 18748 27896 18760
rect 27663 18720 27896 18748
rect 27663 18717 27675 18720
rect 27617 18711 27675 18717
rect 27890 18708 27896 18720
rect 27948 18708 27954 18760
rect 28000 18757 28028 18788
rect 28353 18785 28365 18819
rect 28399 18816 28411 18819
rect 31018 18816 31024 18828
rect 28399 18788 31024 18816
rect 28399 18785 28411 18788
rect 28353 18779 28411 18785
rect 27985 18751 28043 18757
rect 27985 18717 27997 18751
rect 28031 18717 28043 18751
rect 27985 18711 28043 18717
rect 28074 18708 28080 18760
rect 28132 18748 28138 18760
rect 28169 18751 28227 18757
rect 28169 18748 28181 18751
rect 28132 18720 28181 18748
rect 28132 18708 28138 18720
rect 28169 18717 28181 18720
rect 28215 18717 28227 18751
rect 28169 18711 28227 18717
rect 28258 18708 28264 18760
rect 28316 18708 28322 18760
rect 24995 18652 25452 18680
rect 24995 18649 25007 18652
rect 24949 18643 25007 18649
rect 26970 18640 26976 18692
rect 27028 18640 27034 18692
rect 27203 18683 27261 18689
rect 27203 18649 27215 18683
rect 27249 18680 27261 18683
rect 27706 18680 27712 18692
rect 27249 18652 27712 18680
rect 27249 18649 27261 18652
rect 27203 18643 27261 18649
rect 27706 18640 27712 18652
rect 27764 18640 27770 18692
rect 27801 18683 27859 18689
rect 27801 18649 27813 18683
rect 27847 18680 27859 18683
rect 28368 18680 28396 18779
rect 31018 18776 31024 18788
rect 31076 18776 31082 18828
rect 31478 18776 31484 18828
rect 31536 18816 31542 18828
rect 31849 18819 31907 18825
rect 31849 18816 31861 18819
rect 31536 18788 31861 18816
rect 31536 18776 31542 18788
rect 31849 18785 31861 18788
rect 31895 18785 31907 18819
rect 31849 18779 31907 18785
rect 33134 18776 33140 18828
rect 33192 18776 33198 18828
rect 28442 18708 28448 18760
rect 28500 18748 28506 18760
rect 28537 18751 28595 18757
rect 28537 18748 28549 18751
rect 28500 18720 28549 18748
rect 28500 18708 28506 18720
rect 28537 18717 28549 18720
rect 28583 18717 28595 18751
rect 28537 18711 28595 18717
rect 28810 18708 28816 18760
rect 28868 18708 28874 18760
rect 28994 18708 29000 18760
rect 29052 18708 29058 18760
rect 29178 18708 29184 18760
rect 29236 18708 29242 18760
rect 29546 18708 29552 18760
rect 29604 18708 29610 18760
rect 29733 18751 29791 18757
rect 29733 18717 29745 18751
rect 29779 18748 29791 18751
rect 30190 18748 30196 18760
rect 29779 18720 30196 18748
rect 29779 18717 29791 18720
rect 29733 18711 29791 18717
rect 30190 18708 30196 18720
rect 30248 18708 30254 18760
rect 32122 18708 32128 18760
rect 32180 18708 32186 18760
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32401 18751 32459 18757
rect 32401 18748 32413 18751
rect 32272 18720 32413 18748
rect 32272 18708 32278 18720
rect 32401 18717 32413 18720
rect 32447 18717 32459 18751
rect 32401 18711 32459 18717
rect 32766 18708 32772 18760
rect 32824 18708 32830 18760
rect 33336 18748 33364 18924
rect 33502 18912 33508 18924
rect 33560 18952 33566 18964
rect 34422 18952 34428 18964
rect 33560 18924 34428 18952
rect 33560 18912 33566 18924
rect 34422 18912 34428 18924
rect 34480 18912 34486 18964
rect 34885 18955 34943 18961
rect 34885 18921 34897 18955
rect 34931 18952 34943 18955
rect 35710 18952 35716 18964
rect 34931 18924 35716 18952
rect 34931 18921 34943 18924
rect 34885 18915 34943 18921
rect 35710 18912 35716 18924
rect 35768 18912 35774 18964
rect 35989 18955 36047 18961
rect 35989 18921 36001 18955
rect 36035 18952 36047 18955
rect 36078 18952 36084 18964
rect 36035 18924 36084 18952
rect 36035 18921 36047 18924
rect 35989 18915 36047 18921
rect 33410 18844 33416 18896
rect 33468 18884 33474 18896
rect 33689 18887 33747 18893
rect 33689 18884 33701 18887
rect 33468 18856 33701 18884
rect 33468 18844 33474 18856
rect 33689 18853 33701 18856
rect 33735 18853 33747 18887
rect 33689 18847 33747 18853
rect 34701 18887 34759 18893
rect 34701 18853 34713 18887
rect 34747 18853 34759 18887
rect 36004 18884 36032 18915
rect 36078 18912 36084 18924
rect 36136 18912 36142 18964
rect 34701 18847 34759 18853
rect 35544 18856 36032 18884
rect 33704 18816 33732 18847
rect 33704 18788 34100 18816
rect 33413 18751 33471 18757
rect 33413 18748 33425 18751
rect 33336 18720 33425 18748
rect 33413 18717 33425 18720
rect 33459 18717 33471 18751
rect 33413 18711 33471 18717
rect 33502 18708 33508 18760
rect 33560 18748 33566 18760
rect 33965 18751 34023 18757
rect 33965 18748 33977 18751
rect 33560 18720 33977 18748
rect 33560 18708 33566 18720
rect 33965 18717 33977 18720
rect 34011 18717 34023 18751
rect 33965 18711 34023 18717
rect 27847 18652 28396 18680
rect 27847 18649 27859 18652
rect 27801 18643 27859 18649
rect 29086 18640 29092 18692
rect 29144 18640 29150 18692
rect 29270 18640 29276 18692
rect 29328 18680 29334 18692
rect 29328 18652 29960 18680
rect 29328 18640 29334 18652
rect 29932 18624 29960 18652
rect 30834 18640 30840 18692
rect 30892 18680 30898 18692
rect 31389 18683 31447 18689
rect 31389 18680 31401 18683
rect 30892 18652 31401 18680
rect 30892 18640 30898 18652
rect 31389 18649 31401 18652
rect 31435 18680 31447 18683
rect 31478 18680 31484 18692
rect 31435 18652 31484 18680
rect 31435 18649 31447 18652
rect 31389 18643 31447 18649
rect 31478 18640 31484 18652
rect 31536 18640 31542 18692
rect 31573 18683 31631 18689
rect 31573 18649 31585 18683
rect 31619 18680 31631 18683
rect 32582 18680 32588 18692
rect 31619 18652 32588 18680
rect 31619 18649 31631 18652
rect 31573 18643 31631 18649
rect 23400 18584 23704 18612
rect 23750 18572 23756 18624
rect 23808 18572 23814 18624
rect 24118 18572 24124 18624
rect 24176 18572 24182 18624
rect 26697 18615 26755 18621
rect 26697 18581 26709 18615
rect 26743 18612 26755 18615
rect 28902 18612 28908 18624
rect 26743 18584 28908 18612
rect 26743 18581 26755 18584
rect 26697 18575 26755 18581
rect 28902 18572 28908 18584
rect 28960 18572 28966 18624
rect 29362 18572 29368 18624
rect 29420 18572 29426 18624
rect 29638 18572 29644 18624
rect 29696 18572 29702 18624
rect 29914 18572 29920 18624
rect 29972 18612 29978 18624
rect 31588 18612 31616 18643
rect 32582 18640 32588 18652
rect 32640 18640 32646 18692
rect 33686 18640 33692 18692
rect 33744 18640 33750 18692
rect 34072 18680 34100 18788
rect 34146 18776 34152 18828
rect 34204 18776 34210 18828
rect 34241 18819 34299 18825
rect 34241 18785 34253 18819
rect 34287 18816 34299 18819
rect 34716 18816 34744 18847
rect 34974 18816 34980 18828
rect 34287 18788 34980 18816
rect 34287 18785 34299 18788
rect 34241 18779 34299 18785
rect 34974 18776 34980 18788
rect 35032 18776 35038 18828
rect 34333 18751 34391 18757
rect 34333 18717 34345 18751
rect 34379 18717 34391 18751
rect 34333 18711 34391 18717
rect 34517 18751 34575 18757
rect 34517 18717 34529 18751
rect 34563 18748 34575 18751
rect 35544 18748 35572 18856
rect 36170 18844 36176 18896
rect 36228 18844 36234 18896
rect 36817 18887 36875 18893
rect 36817 18853 36829 18887
rect 36863 18853 36875 18887
rect 36817 18847 36875 18853
rect 36354 18816 36360 18828
rect 35912 18788 36360 18816
rect 35912 18757 35940 18788
rect 36354 18776 36360 18788
rect 36412 18816 36418 18828
rect 36832 18816 36860 18847
rect 37274 18844 37280 18896
rect 37332 18884 37338 18896
rect 37734 18884 37740 18896
rect 37332 18856 37740 18884
rect 37332 18844 37338 18856
rect 37734 18844 37740 18856
rect 37792 18844 37798 18896
rect 36412 18788 36860 18816
rect 36412 18776 36418 18788
rect 36556 18757 36584 18788
rect 34563 18720 35572 18748
rect 35897 18751 35955 18757
rect 34563 18717 34575 18720
rect 34517 18711 34575 18717
rect 35897 18717 35909 18751
rect 35943 18717 35955 18751
rect 35897 18711 35955 18717
rect 36081 18751 36139 18757
rect 36081 18717 36093 18751
rect 36127 18748 36139 18751
rect 36541 18751 36599 18757
rect 36127 18720 36400 18748
rect 36127 18717 36139 18720
rect 36081 18711 36139 18717
rect 34348 18680 34376 18711
rect 34072 18652 34376 18680
rect 34422 18640 34428 18692
rect 34480 18680 34486 18692
rect 36372 18689 36400 18720
rect 36541 18717 36553 18751
rect 36587 18717 36599 18751
rect 36541 18711 36599 18717
rect 36630 18708 36636 18760
rect 36688 18748 36694 18760
rect 37458 18748 37464 18760
rect 36688 18720 37464 18748
rect 36688 18708 36694 18720
rect 37458 18708 37464 18720
rect 37516 18708 37522 18760
rect 34853 18683 34911 18689
rect 34853 18680 34865 18683
rect 34480 18652 34865 18680
rect 34480 18640 34486 18652
rect 34853 18649 34865 18652
rect 34899 18649 34911 18683
rect 34853 18643 34911 18649
rect 35069 18683 35127 18689
rect 35069 18649 35081 18683
rect 35115 18649 35127 18683
rect 35069 18643 35127 18649
rect 36357 18683 36415 18689
rect 36357 18649 36369 18683
rect 36403 18649 36415 18683
rect 36357 18643 36415 18649
rect 29972 18584 31616 18612
rect 33505 18615 33563 18621
rect 29972 18572 29978 18584
rect 33505 18581 33517 18615
rect 33551 18612 33563 18615
rect 33594 18612 33600 18624
rect 33551 18584 33600 18612
rect 33551 18581 33563 18584
rect 33505 18575 33563 18581
rect 33594 18572 33600 18584
rect 33652 18572 33658 18624
rect 33781 18615 33839 18621
rect 33781 18581 33793 18615
rect 33827 18612 33839 18615
rect 34606 18612 34612 18624
rect 33827 18584 34612 18612
rect 33827 18581 33839 18584
rect 33781 18575 33839 18581
rect 34606 18572 34612 18584
rect 34664 18572 34670 18624
rect 34698 18572 34704 18624
rect 34756 18612 34762 18624
rect 35084 18612 35112 18643
rect 34756 18584 35112 18612
rect 34756 18572 34762 18584
rect 35250 18572 35256 18624
rect 35308 18612 35314 18624
rect 36372 18612 36400 18643
rect 37090 18640 37096 18692
rect 37148 18640 37154 18692
rect 37274 18612 37280 18624
rect 35308 18584 37280 18612
rect 35308 18572 35314 18584
rect 37274 18572 37280 18584
rect 37332 18572 37338 18624
rect 1104 18522 38824 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 38824 18522
rect 1104 18448 38824 18470
rect 4522 18368 4528 18420
rect 4580 18368 4586 18420
rect 7837 18411 7895 18417
rect 7837 18377 7849 18411
rect 7883 18408 7895 18411
rect 7883 18380 8156 18408
rect 7883 18377 7895 18380
rect 7837 18371 7895 18377
rect 4706 18340 4712 18352
rect 3528 18312 4712 18340
rect 2866 18232 2872 18284
rect 2924 18232 2930 18284
rect 3528 18281 3556 18312
rect 4706 18300 4712 18312
rect 4764 18340 4770 18352
rect 7469 18343 7527 18349
rect 4764 18312 6040 18340
rect 4764 18300 4770 18312
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18241 3571 18275
rect 3513 18235 3571 18241
rect 3786 18232 3792 18284
rect 3844 18272 3850 18284
rect 3973 18275 4031 18281
rect 3973 18272 3985 18275
rect 3844 18244 3985 18272
rect 3844 18232 3850 18244
rect 3973 18241 3985 18244
rect 4019 18241 4031 18275
rect 3973 18235 4031 18241
rect 4341 18275 4399 18281
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 4430 18272 4436 18284
rect 4387 18244 4436 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 4430 18232 4436 18244
rect 4488 18232 4494 18284
rect 4890 18232 4896 18284
rect 4948 18232 4954 18284
rect 4982 18232 4988 18284
rect 5040 18232 5046 18284
rect 6012 18281 6040 18312
rect 7469 18309 7481 18343
rect 7515 18340 7527 18343
rect 7558 18340 7564 18352
rect 7515 18312 7564 18340
rect 7515 18309 7527 18312
rect 7469 18303 7527 18309
rect 7558 18300 7564 18312
rect 7616 18300 7622 18352
rect 7685 18343 7743 18349
rect 7685 18309 7697 18343
rect 7731 18340 7743 18343
rect 7926 18340 7932 18352
rect 7731 18312 7932 18340
rect 7731 18309 7743 18312
rect 7685 18303 7743 18309
rect 7926 18300 7932 18312
rect 7984 18300 7990 18352
rect 8128 18340 8156 18380
rect 8478 18368 8484 18420
rect 8536 18368 8542 18420
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 9125 18411 9183 18417
rect 9125 18408 9137 18411
rect 8720 18380 9137 18408
rect 8720 18368 8726 18380
rect 9125 18377 9137 18380
rect 9171 18377 9183 18411
rect 9125 18371 9183 18377
rect 9398 18368 9404 18420
rect 9456 18408 9462 18420
rect 10045 18411 10103 18417
rect 10045 18408 10057 18411
rect 9456 18380 10057 18408
rect 9456 18368 9462 18380
rect 10045 18377 10057 18380
rect 10091 18377 10103 18411
rect 10045 18371 10103 18377
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 10376 18380 10517 18408
rect 10376 18368 10382 18380
rect 10505 18377 10517 18380
rect 10551 18377 10563 18411
rect 10505 18371 10563 18377
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 13814 18408 13820 18420
rect 13771 18380 13820 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 14277 18411 14335 18417
rect 14277 18377 14289 18411
rect 14323 18408 14335 18411
rect 15194 18408 15200 18420
rect 14323 18380 15200 18408
rect 14323 18377 14335 18380
rect 14277 18371 14335 18377
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 16485 18411 16543 18417
rect 16485 18377 16497 18411
rect 16531 18408 16543 18411
rect 16758 18408 16764 18420
rect 16531 18380 16764 18408
rect 16531 18377 16543 18380
rect 16485 18371 16543 18377
rect 16758 18368 16764 18380
rect 16816 18368 16822 18420
rect 17586 18368 17592 18420
rect 17644 18408 17650 18420
rect 22557 18411 22615 18417
rect 17644 18380 19840 18408
rect 17644 18368 17650 18380
rect 8496 18340 8524 18368
rect 14918 18340 14924 18352
rect 8128 18312 9444 18340
rect 8128 18281 8156 18312
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18272 5227 18275
rect 5261 18275 5319 18281
rect 5261 18272 5273 18275
rect 5215 18244 5273 18272
rect 5215 18241 5227 18244
rect 5169 18235 5227 18241
rect 5261 18241 5273 18244
rect 5307 18241 5319 18275
rect 5261 18235 5319 18241
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18241 6239 18275
rect 6181 18235 6239 18241
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18241 8171 18275
rect 8113 18235 8171 18241
rect 1394 18164 1400 18216
rect 1452 18204 1458 18216
rect 1489 18207 1547 18213
rect 1489 18204 1501 18207
rect 1452 18176 1501 18204
rect 1452 18164 1458 18176
rect 1489 18173 1501 18176
rect 1535 18173 1547 18207
rect 1489 18167 1547 18173
rect 1762 18164 1768 18216
rect 1820 18164 1826 18216
rect 3234 18164 3240 18216
rect 3292 18204 3298 18216
rect 3697 18207 3755 18213
rect 3697 18204 3709 18207
rect 3292 18176 3709 18204
rect 3292 18164 3298 18176
rect 3697 18173 3709 18176
rect 3743 18173 3755 18207
rect 3697 18167 3755 18173
rect 2958 18096 2964 18148
rect 3016 18136 3022 18148
rect 3329 18139 3387 18145
rect 3329 18136 3341 18139
rect 3016 18108 3341 18136
rect 3016 18096 3022 18108
rect 3329 18105 3341 18108
rect 3375 18136 3387 18139
rect 3418 18136 3424 18148
rect 3375 18108 3424 18136
rect 3375 18105 3387 18108
rect 3329 18099 3387 18105
rect 3418 18096 3424 18108
rect 3476 18096 3482 18148
rect 3712 18136 3740 18167
rect 3878 18164 3884 18216
rect 3936 18164 3942 18216
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 5092 18176 5825 18204
rect 4062 18136 4068 18148
rect 3712 18108 4068 18136
rect 4062 18096 4068 18108
rect 4120 18096 4126 18148
rect 5092 18080 5120 18176
rect 5813 18173 5825 18176
rect 5859 18173 5871 18207
rect 5813 18167 5871 18173
rect 5169 18139 5227 18145
rect 5169 18105 5181 18139
rect 5215 18136 5227 18139
rect 6196 18136 6224 18235
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 8352 18244 8493 18272
rect 8352 18232 8358 18244
rect 8481 18241 8493 18244
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8754 18232 8760 18284
rect 8812 18272 8818 18284
rect 9416 18281 9444 18312
rect 12912 18312 14924 18340
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 8812 18244 9229 18272
rect 8812 18232 8818 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18241 9459 18275
rect 9401 18235 9459 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18272 10471 18275
rect 10870 18272 10876 18284
rect 10459 18244 10876 18272
rect 10459 18241 10471 18244
rect 10413 18235 10471 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 12618 18232 12624 18284
rect 12676 18232 12682 18284
rect 12912 18281 12940 18312
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 13262 18232 13268 18284
rect 13320 18232 13326 18284
rect 13354 18232 13360 18284
rect 13412 18272 13418 18284
rect 13541 18275 13599 18281
rect 13541 18272 13553 18275
rect 13412 18244 13553 18272
rect 13412 18232 13418 18244
rect 13541 18241 13553 18244
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 13814 18232 13820 18284
rect 13872 18232 13878 18284
rect 14108 18281 14136 18312
rect 14918 18300 14924 18312
rect 14976 18300 14982 18352
rect 15013 18343 15071 18349
rect 15013 18309 15025 18343
rect 15059 18340 15071 18343
rect 15286 18340 15292 18352
rect 15059 18312 15292 18340
rect 15059 18309 15071 18312
rect 15013 18303 15071 18309
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 17126 18300 17132 18352
rect 17184 18300 17190 18352
rect 17359 18343 17417 18349
rect 17359 18309 17371 18343
rect 17405 18340 17417 18343
rect 17678 18340 17684 18352
rect 17405 18312 17684 18340
rect 17405 18309 17417 18312
rect 17359 18303 17417 18309
rect 17678 18300 17684 18312
rect 17736 18300 17742 18352
rect 17862 18300 17868 18352
rect 17920 18340 17926 18352
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 17920 18312 18245 18340
rect 17920 18300 17926 18312
rect 18233 18309 18245 18312
rect 18279 18309 18291 18343
rect 19518 18340 19524 18352
rect 19458 18326 19524 18340
rect 18233 18303 18291 18309
rect 19444 18312 19524 18326
rect 14093 18275 14151 18281
rect 14093 18272 14105 18275
rect 13924 18244 14105 18272
rect 7466 18164 7472 18216
rect 7524 18204 7530 18216
rect 7929 18207 7987 18213
rect 7929 18204 7941 18207
rect 7524 18176 7941 18204
rect 7524 18164 7530 18176
rect 7929 18173 7941 18176
rect 7975 18173 7987 18207
rect 7929 18167 7987 18173
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 9180 18176 9321 18204
rect 9180 18164 9186 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 11882 18164 11888 18216
rect 11940 18204 11946 18216
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 11940 18176 12081 18204
rect 11940 18164 11946 18176
rect 12069 18173 12081 18176
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12584 18176 12817 18204
rect 12584 18164 12590 18176
rect 12805 18173 12817 18176
rect 12851 18204 12863 18207
rect 12851 18176 13584 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 5215 18108 6224 18136
rect 12713 18139 12771 18145
rect 5215 18105 5227 18108
rect 5169 18099 5227 18105
rect 12713 18105 12725 18139
rect 12759 18136 12771 18139
rect 12986 18136 12992 18148
rect 12759 18108 12992 18136
rect 12759 18105 12771 18108
rect 12713 18099 12771 18105
rect 12986 18096 12992 18108
rect 13044 18096 13050 18148
rect 13081 18139 13139 18145
rect 13081 18105 13093 18139
rect 13127 18136 13139 18139
rect 13357 18139 13415 18145
rect 13357 18136 13369 18139
rect 13127 18108 13369 18136
rect 13127 18105 13139 18108
rect 13081 18099 13139 18105
rect 13357 18105 13369 18108
rect 13403 18105 13415 18139
rect 13357 18099 13415 18105
rect 13446 18096 13452 18148
rect 13504 18096 13510 18148
rect 13556 18080 13584 18176
rect 13722 18164 13728 18216
rect 13780 18204 13786 18216
rect 13924 18204 13952 18244
rect 14093 18241 14105 18244
rect 14139 18241 14151 18275
rect 14093 18235 14151 18241
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 13780 18176 13952 18204
rect 13780 18164 13786 18176
rect 13998 18164 14004 18216
rect 14056 18164 14062 18216
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 14240 18176 14381 18204
rect 14240 18164 14246 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14660 18204 14688 18235
rect 14734 18232 14740 18284
rect 14792 18232 14798 18284
rect 16114 18232 16120 18284
rect 16172 18232 16178 18284
rect 17034 18232 17040 18284
rect 17092 18232 17098 18284
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 17770 18272 17776 18284
rect 17543 18244 17776 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 17954 18232 17960 18284
rect 18012 18232 18018 18284
rect 15010 18204 15016 18216
rect 14660 18176 15016 18204
rect 14369 18167 14427 18173
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 17310 18164 17316 18216
rect 17368 18204 17374 18216
rect 17865 18207 17923 18213
rect 17865 18204 17877 18207
rect 17368 18176 17877 18204
rect 17368 18164 17374 18176
rect 17865 18173 17877 18176
rect 17911 18204 17923 18207
rect 19444 18204 19472 18312
rect 19518 18300 19524 18312
rect 19576 18300 19582 18352
rect 19812 18272 19840 18380
rect 22557 18377 22569 18411
rect 22603 18408 22615 18411
rect 22922 18408 22928 18420
rect 22603 18380 22928 18408
rect 22603 18377 22615 18380
rect 22557 18371 22615 18377
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 24397 18411 24455 18417
rect 24397 18377 24409 18411
rect 24443 18408 24455 18411
rect 24854 18408 24860 18420
rect 24443 18380 24860 18408
rect 24443 18377 24455 18380
rect 24397 18371 24455 18377
rect 24854 18368 24860 18380
rect 24912 18368 24918 18420
rect 25314 18368 25320 18420
rect 25372 18408 25378 18420
rect 25409 18411 25467 18417
rect 25409 18408 25421 18411
rect 25372 18380 25421 18408
rect 25372 18368 25378 18380
rect 25409 18377 25421 18380
rect 25455 18377 25467 18411
rect 25409 18371 25467 18377
rect 28169 18411 28227 18417
rect 28169 18377 28181 18411
rect 28215 18408 28227 18411
rect 28258 18408 28264 18420
rect 28215 18380 28264 18408
rect 28215 18377 28227 18380
rect 28169 18371 28227 18377
rect 28258 18368 28264 18380
rect 28316 18368 28322 18420
rect 28445 18411 28503 18417
rect 28445 18377 28457 18411
rect 28491 18408 28503 18411
rect 28810 18408 28816 18420
rect 28491 18380 28816 18408
rect 28491 18377 28503 18380
rect 28445 18371 28503 18377
rect 28810 18368 28816 18380
rect 28868 18368 28874 18420
rect 31757 18411 31815 18417
rect 31757 18377 31769 18411
rect 31803 18408 31815 18411
rect 31803 18380 34376 18408
rect 31803 18377 31815 18380
rect 31757 18371 31815 18377
rect 23474 18300 23480 18352
rect 23532 18340 23538 18352
rect 23532 18312 24256 18340
rect 23532 18300 23538 18312
rect 19981 18275 20039 18281
rect 19981 18272 19993 18275
rect 19812 18244 19993 18272
rect 19981 18241 19993 18244
rect 20027 18272 20039 18275
rect 20070 18272 20076 18284
rect 20027 18244 20076 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22462 18272 22468 18284
rect 22235 18244 22468 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22462 18232 22468 18244
rect 22520 18232 22526 18284
rect 23566 18232 23572 18284
rect 23624 18232 23630 18284
rect 24228 18281 24256 18312
rect 27246 18300 27252 18352
rect 27304 18340 27310 18352
rect 27801 18343 27859 18349
rect 27801 18340 27813 18343
rect 27304 18312 27813 18340
rect 27304 18300 27310 18312
rect 27801 18309 27813 18312
rect 27847 18340 27859 18343
rect 27847 18312 28580 18340
rect 27847 18309 27859 18312
rect 27801 18303 27859 18309
rect 24213 18275 24271 18281
rect 24213 18241 24225 18275
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 24854 18232 24860 18284
rect 24912 18272 24918 18284
rect 24949 18275 25007 18281
rect 24949 18272 24961 18275
rect 24912 18244 24961 18272
rect 24912 18232 24918 18244
rect 24949 18241 24961 18244
rect 24995 18272 25007 18275
rect 25593 18275 25651 18281
rect 25593 18272 25605 18275
rect 24995 18244 25605 18272
rect 24995 18241 25007 18244
rect 24949 18235 25007 18241
rect 25593 18241 25605 18244
rect 25639 18241 25651 18275
rect 25593 18235 25651 18241
rect 25685 18275 25743 18281
rect 25685 18241 25697 18275
rect 25731 18272 25743 18275
rect 26142 18272 26148 18284
rect 25731 18244 26148 18272
rect 25731 18241 25743 18244
rect 25685 18235 25743 18241
rect 17911 18176 19472 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 21266 18164 21272 18216
rect 21324 18204 21330 18216
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 21324 18176 22293 18204
rect 21324 18164 21330 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 23934 18164 23940 18216
rect 23992 18164 23998 18216
rect 25041 18207 25099 18213
rect 25041 18173 25053 18207
rect 25087 18204 25099 18207
rect 25409 18207 25467 18213
rect 25409 18204 25421 18207
rect 25087 18176 25421 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 25409 18173 25421 18176
rect 25455 18204 25467 18207
rect 25498 18204 25504 18216
rect 25455 18176 25504 18204
rect 25455 18173 25467 18176
rect 25409 18167 25467 18173
rect 14461 18139 14519 18145
rect 14461 18105 14473 18139
rect 14507 18136 14519 18139
rect 14507 18108 14872 18136
rect 14507 18105 14519 18108
rect 14461 18099 14519 18105
rect 3970 18028 3976 18080
rect 4028 18068 4034 18080
rect 4249 18071 4307 18077
rect 4249 18068 4261 18071
rect 4028 18040 4261 18068
rect 4028 18028 4034 18040
rect 4249 18037 4261 18040
rect 4295 18037 4307 18071
rect 4249 18031 4307 18037
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 5074 18068 5080 18080
rect 4396 18040 5080 18068
rect 4396 18028 4402 18040
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 6181 18071 6239 18077
rect 6181 18037 6193 18071
rect 6227 18068 6239 18071
rect 6546 18068 6552 18080
rect 6227 18040 6552 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 7558 18028 7564 18080
rect 7616 18068 7622 18080
rect 7653 18071 7711 18077
rect 7653 18068 7665 18071
rect 7616 18040 7665 18068
rect 7616 18028 7622 18040
rect 7653 18037 7665 18040
rect 7699 18037 7711 18071
rect 7653 18031 7711 18037
rect 11517 18071 11575 18077
rect 11517 18037 11529 18071
rect 11563 18068 11575 18071
rect 11974 18068 11980 18080
rect 11563 18040 11980 18068
rect 11563 18037 11575 18040
rect 11517 18031 11575 18037
rect 11974 18028 11980 18040
rect 12032 18028 12038 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 13817 18071 13875 18077
rect 13817 18068 13829 18071
rect 13596 18040 13829 18068
rect 13596 18028 13602 18040
rect 13817 18037 13829 18040
rect 13863 18037 13875 18071
rect 13817 18031 13875 18037
rect 14550 18028 14556 18080
rect 14608 18028 14614 18080
rect 14844 18068 14872 18108
rect 17678 18096 17684 18148
rect 17736 18136 17742 18148
rect 17736 18108 18092 18136
rect 17736 18096 17742 18108
rect 16022 18068 16028 18080
rect 14844 18040 16028 18068
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 16853 18071 16911 18077
rect 16853 18037 16865 18071
rect 16899 18068 16911 18071
rect 16942 18068 16948 18080
rect 16899 18040 16948 18068
rect 16899 18037 16911 18040
rect 16853 18031 16911 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 18064 18068 18092 18108
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 25056 18136 25084 18167
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 25700 18136 25728 18235
rect 26142 18232 26148 18244
rect 26200 18232 26206 18284
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18241 27675 18275
rect 27617 18235 27675 18241
rect 28077 18275 28135 18281
rect 28077 18241 28089 18275
rect 28123 18272 28135 18275
rect 28166 18272 28172 18284
rect 28123 18244 28172 18272
rect 28123 18241 28135 18244
rect 28077 18235 28135 18241
rect 27632 18204 27660 18235
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 28258 18232 28264 18284
rect 28316 18272 28322 18284
rect 28552 18281 28580 18312
rect 29178 18300 29184 18352
rect 29236 18340 29242 18352
rect 30650 18340 30656 18352
rect 29236 18312 29960 18340
rect 29236 18300 29242 18312
rect 28353 18275 28411 18281
rect 28353 18272 28365 18275
rect 28316 18244 28365 18272
rect 28316 18232 28322 18244
rect 28353 18241 28365 18244
rect 28399 18241 28411 18275
rect 28353 18235 28411 18241
rect 28537 18275 28595 18281
rect 28537 18241 28549 18275
rect 28583 18241 28595 18275
rect 28537 18235 28595 18241
rect 27706 18204 27712 18216
rect 27632 18176 27712 18204
rect 27706 18164 27712 18176
rect 27764 18204 27770 18216
rect 28442 18204 28448 18216
rect 27764 18176 28448 18204
rect 27764 18164 27770 18176
rect 28442 18164 28448 18176
rect 28500 18164 28506 18216
rect 23808 18108 25084 18136
rect 25148 18108 25728 18136
rect 28552 18136 28580 18235
rect 28994 18232 29000 18284
rect 29052 18232 29058 18284
rect 29362 18232 29368 18284
rect 29420 18272 29426 18284
rect 29825 18275 29883 18281
rect 29825 18272 29837 18275
rect 29420 18244 29837 18272
rect 29420 18232 29426 18244
rect 29825 18241 29837 18244
rect 29871 18241 29883 18275
rect 29932 18272 29960 18312
rect 30208 18312 30656 18340
rect 30208 18281 30236 18312
rect 30650 18300 30656 18312
rect 30708 18340 30714 18352
rect 31386 18340 31392 18352
rect 30708 18312 31392 18340
rect 30708 18300 30714 18312
rect 31386 18300 31392 18312
rect 31444 18300 31450 18352
rect 32122 18300 32128 18352
rect 32180 18340 32186 18352
rect 32180 18312 33916 18340
rect 32180 18300 32186 18312
rect 30009 18275 30067 18281
rect 30009 18272 30021 18275
rect 29932 18244 30021 18272
rect 29825 18235 29883 18241
rect 30009 18241 30021 18244
rect 30055 18241 30067 18275
rect 30009 18235 30067 18241
rect 30193 18275 30251 18281
rect 30193 18241 30205 18275
rect 30239 18241 30251 18275
rect 30193 18235 30251 18241
rect 30377 18275 30435 18281
rect 30377 18241 30389 18275
rect 30423 18241 30435 18275
rect 30377 18235 30435 18241
rect 30561 18275 30619 18281
rect 30561 18241 30573 18275
rect 30607 18272 30619 18275
rect 31113 18275 31171 18281
rect 31113 18272 31125 18275
rect 30607 18244 31125 18272
rect 30607 18241 30619 18244
rect 30561 18235 30619 18241
rect 31113 18241 31125 18244
rect 31159 18241 31171 18275
rect 31113 18235 31171 18241
rect 31206 18275 31264 18281
rect 31206 18241 31218 18275
rect 31252 18241 31264 18275
rect 31206 18235 31264 18241
rect 31481 18275 31539 18281
rect 31481 18241 31493 18275
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 31619 18275 31677 18281
rect 31619 18241 31631 18275
rect 31665 18272 31677 18275
rect 32030 18272 32036 18284
rect 31665 18244 32036 18272
rect 31665 18241 31677 18244
rect 31619 18235 31677 18241
rect 29086 18164 29092 18216
rect 29144 18204 29150 18216
rect 30101 18207 30159 18213
rect 30101 18204 30113 18207
rect 29144 18176 30113 18204
rect 29144 18164 29150 18176
rect 30101 18173 30113 18176
rect 30147 18173 30159 18207
rect 30392 18204 30420 18235
rect 30926 18204 30932 18216
rect 30392 18176 30932 18204
rect 30101 18167 30159 18173
rect 30926 18164 30932 18176
rect 30984 18204 30990 18216
rect 31220 18204 31248 18235
rect 30984 18176 31248 18204
rect 30984 18164 30990 18176
rect 31496 18136 31524 18235
rect 32030 18232 32036 18244
rect 32088 18272 32094 18284
rect 33042 18272 33048 18284
rect 32088 18244 33048 18272
rect 32088 18232 32094 18244
rect 33042 18232 33048 18244
rect 33100 18232 33106 18284
rect 33410 18232 33416 18284
rect 33468 18232 33474 18284
rect 33505 18275 33563 18281
rect 33505 18241 33517 18275
rect 33551 18241 33563 18275
rect 33505 18235 33563 18241
rect 33226 18204 33232 18216
rect 33152 18176 33232 18204
rect 28552 18108 31524 18136
rect 23808 18096 23814 18108
rect 19610 18068 19616 18080
rect 18064 18040 19616 18068
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 21910 18028 21916 18080
rect 21968 18068 21974 18080
rect 25148 18077 25176 18108
rect 22189 18071 22247 18077
rect 22189 18068 22201 18071
rect 21968 18040 22201 18068
rect 21968 18028 21974 18040
rect 22189 18037 22201 18040
rect 22235 18037 22247 18071
rect 22189 18031 22247 18037
rect 23661 18071 23719 18077
rect 23661 18037 23673 18071
rect 23707 18068 23719 18071
rect 24029 18071 24087 18077
rect 24029 18068 24041 18071
rect 23707 18040 24041 18068
rect 23707 18037 23719 18040
rect 23661 18031 23719 18037
rect 24029 18037 24041 18040
rect 24075 18037 24087 18071
rect 24029 18031 24087 18037
rect 25133 18071 25191 18077
rect 25133 18037 25145 18071
rect 25179 18037 25191 18071
rect 25133 18031 25191 18037
rect 25317 18071 25375 18077
rect 25317 18037 25329 18071
rect 25363 18068 25375 18071
rect 25406 18068 25412 18080
rect 25363 18040 25412 18068
rect 25363 18037 25375 18040
rect 25317 18031 25375 18037
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 27985 18071 28043 18077
rect 27985 18037 27997 18071
rect 28031 18068 28043 18071
rect 28718 18068 28724 18080
rect 28031 18040 28724 18068
rect 28031 18037 28043 18040
rect 27985 18031 28043 18037
rect 28718 18028 28724 18040
rect 28776 18028 28782 18080
rect 31496 18068 31524 18108
rect 31662 18096 31668 18148
rect 31720 18136 31726 18148
rect 33152 18136 33180 18176
rect 33226 18164 33232 18176
rect 33284 18164 33290 18216
rect 33520 18204 33548 18235
rect 33594 18204 33600 18216
rect 33520 18176 33600 18204
rect 33594 18164 33600 18176
rect 33652 18164 33658 18216
rect 33888 18145 33916 18312
rect 34348 18281 34376 18380
rect 34422 18368 34428 18420
rect 34480 18408 34486 18420
rect 37366 18408 37372 18420
rect 34480 18380 37372 18408
rect 34480 18368 34486 18380
rect 37366 18368 37372 18380
rect 37424 18368 37430 18420
rect 34514 18300 34520 18352
rect 34572 18340 34578 18352
rect 35069 18343 35127 18349
rect 35069 18340 35081 18343
rect 34572 18312 35081 18340
rect 34572 18300 34578 18312
rect 35069 18309 35081 18312
rect 35115 18309 35127 18343
rect 35069 18303 35127 18309
rect 34333 18275 34391 18281
rect 34333 18241 34345 18275
rect 34379 18241 34391 18275
rect 34333 18235 34391 18241
rect 34606 18232 34612 18284
rect 34664 18232 34670 18284
rect 34698 18232 34704 18284
rect 34756 18272 34762 18284
rect 34974 18272 34980 18284
rect 34756 18244 34980 18272
rect 34756 18232 34762 18244
rect 34974 18232 34980 18244
rect 35032 18232 35038 18284
rect 35250 18232 35256 18284
rect 35308 18232 35314 18284
rect 34422 18164 34428 18216
rect 34480 18204 34486 18216
rect 35268 18204 35296 18232
rect 34480 18176 35296 18204
rect 34480 18164 34486 18176
rect 31720 18108 33180 18136
rect 33321 18139 33379 18145
rect 31720 18096 31726 18108
rect 33321 18105 33333 18139
rect 33367 18136 33379 18139
rect 33873 18139 33931 18145
rect 33367 18108 33824 18136
rect 33367 18105 33379 18108
rect 33321 18099 33379 18105
rect 33502 18068 33508 18080
rect 31496 18040 33508 18068
rect 33502 18028 33508 18040
rect 33560 18028 33566 18080
rect 33796 18068 33824 18108
rect 33873 18105 33885 18139
rect 33919 18105 33931 18139
rect 33873 18099 33931 18105
rect 34238 18068 34244 18080
rect 33796 18040 34244 18068
rect 34238 18028 34244 18040
rect 34296 18028 34302 18080
rect 35437 18071 35495 18077
rect 35437 18037 35449 18071
rect 35483 18068 35495 18071
rect 35802 18068 35808 18080
rect 35483 18040 35808 18068
rect 35483 18037 35495 18040
rect 35437 18031 35495 18037
rect 35802 18028 35808 18040
rect 35860 18028 35866 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2409 17867 2467 17873
rect 2409 17864 2421 17867
rect 1820 17836 2421 17864
rect 1820 17824 1826 17836
rect 2409 17833 2421 17836
rect 2455 17833 2467 17867
rect 2409 17827 2467 17833
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 4617 17867 4675 17873
rect 4617 17864 4629 17867
rect 2823 17836 4629 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 4617 17833 4629 17836
rect 4663 17864 4675 17867
rect 4706 17864 4712 17876
rect 4663 17836 4712 17864
rect 4663 17833 4675 17836
rect 4617 17827 4675 17833
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 4801 17867 4859 17873
rect 4801 17833 4813 17867
rect 4847 17864 4859 17867
rect 4982 17864 4988 17876
rect 4847 17836 4988 17864
rect 4847 17833 4859 17836
rect 4801 17827 4859 17833
rect 4982 17824 4988 17836
rect 5040 17864 5046 17876
rect 5350 17864 5356 17876
rect 5040 17836 5356 17864
rect 5040 17824 5046 17836
rect 5350 17824 5356 17836
rect 5408 17824 5414 17876
rect 8754 17824 8760 17876
rect 8812 17824 8818 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 11882 17864 11888 17876
rect 10827 17836 11888 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 11882 17824 11888 17836
rect 11940 17864 11946 17876
rect 11940 17836 12434 17864
rect 11940 17824 11946 17836
rect 5074 17756 5080 17808
rect 5132 17756 5138 17808
rect 7285 17799 7343 17805
rect 7285 17765 7297 17799
rect 7331 17796 7343 17799
rect 12406 17796 12434 17836
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12805 17867 12863 17873
rect 12805 17864 12817 17867
rect 12676 17836 12817 17864
rect 12676 17824 12682 17836
rect 12805 17833 12817 17836
rect 12851 17833 12863 17867
rect 12805 17827 12863 17833
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 13814 17864 13820 17876
rect 12952 17836 13820 17864
rect 12952 17824 12958 17836
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 14918 17824 14924 17876
rect 14976 17864 14982 17876
rect 15746 17864 15752 17876
rect 14976 17836 15752 17864
rect 14976 17824 14982 17836
rect 15746 17824 15752 17836
rect 15804 17864 15810 17876
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 15804 17836 15853 17864
rect 15804 17824 15810 17836
rect 15841 17833 15853 17836
rect 15887 17833 15899 17867
rect 15841 17827 15899 17833
rect 18414 17824 18420 17876
rect 18472 17824 18478 17876
rect 19794 17824 19800 17876
rect 19852 17824 19858 17876
rect 24489 17867 24547 17873
rect 24489 17833 24501 17867
rect 24535 17864 24547 17867
rect 24854 17864 24860 17876
rect 24535 17836 24860 17864
rect 24535 17833 24547 17836
rect 24489 17827 24547 17833
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 27246 17824 27252 17876
rect 27304 17824 27310 17876
rect 27982 17824 27988 17876
rect 28040 17864 28046 17876
rect 30190 17864 30196 17876
rect 28040 17836 30196 17864
rect 28040 17824 28046 17836
rect 30190 17824 30196 17836
rect 30248 17864 30254 17876
rect 30834 17864 30840 17876
rect 30248 17836 30840 17864
rect 30248 17824 30254 17836
rect 30834 17824 30840 17836
rect 30892 17824 30898 17876
rect 30926 17824 30932 17876
rect 30984 17824 30990 17876
rect 31726 17836 33180 17864
rect 26786 17796 26792 17808
rect 7331 17768 8156 17796
rect 12406 17768 13032 17796
rect 7331 17765 7343 17768
rect 7285 17759 7343 17765
rect 3053 17731 3111 17737
rect 3053 17728 3065 17731
rect 2608 17700 3065 17728
rect 2608 17669 2636 17700
rect 3053 17697 3065 17700
rect 3099 17697 3111 17731
rect 3053 17691 3111 17697
rect 6546 17688 6552 17740
rect 6604 17688 6610 17740
rect 6822 17688 6828 17740
rect 6880 17688 6886 17740
rect 7926 17688 7932 17740
rect 7984 17688 7990 17740
rect 8128 17737 8156 17768
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17697 8171 17731
rect 10873 17731 10931 17737
rect 10873 17728 10885 17731
rect 8113 17691 8171 17697
rect 9048 17700 10885 17728
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17629 2651 17663
rect 2593 17623 2651 17629
rect 2869 17663 2927 17669
rect 2869 17629 2881 17663
rect 2915 17629 2927 17663
rect 2869 17623 2927 17629
rect 2884 17592 2912 17623
rect 2958 17620 2964 17672
rect 3016 17620 3022 17672
rect 3142 17620 3148 17672
rect 3200 17620 3206 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4430 17660 4436 17672
rect 4212 17632 4436 17660
rect 4212 17620 4218 17632
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 7009 17663 7067 17669
rect 7009 17629 7021 17663
rect 7055 17660 7067 17663
rect 7558 17660 7564 17672
rect 7055 17632 7564 17660
rect 7055 17629 7067 17632
rect 7009 17623 7067 17629
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 9048 17669 9076 17700
rect 10873 17697 10885 17700
rect 10919 17697 10931 17731
rect 10873 17691 10931 17697
rect 12526 17688 12532 17740
rect 12584 17728 12590 17740
rect 12621 17731 12679 17737
rect 12621 17728 12633 17731
rect 12584 17700 12633 17728
rect 12584 17688 12590 17700
rect 12621 17697 12633 17700
rect 12667 17697 12679 17731
rect 12621 17691 12679 17697
rect 9033 17663 9091 17669
rect 9033 17629 9045 17663
rect 9079 17629 9091 17663
rect 9033 17623 9091 17629
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 2884 17564 3801 17592
rect 3789 17561 3801 17564
rect 3835 17561 3847 17595
rect 3789 17555 3847 17561
rect 4522 17552 4528 17604
rect 4580 17592 4586 17604
rect 4985 17595 5043 17601
rect 4985 17592 4997 17595
rect 4580 17564 4997 17592
rect 4580 17552 4586 17564
rect 4985 17561 4997 17564
rect 5031 17592 5043 17595
rect 5074 17592 5080 17604
rect 5031 17564 5080 17592
rect 5031 17561 5043 17564
rect 4985 17555 5043 17561
rect 5074 17552 5080 17564
rect 5132 17552 5138 17604
rect 5902 17552 5908 17604
rect 5960 17552 5966 17604
rect 7285 17595 7343 17601
rect 7285 17561 7297 17595
rect 7331 17592 7343 17595
rect 7377 17595 7435 17601
rect 7377 17592 7389 17595
rect 7331 17564 7389 17592
rect 7331 17561 7343 17564
rect 7285 17555 7343 17561
rect 7377 17561 7389 17564
rect 7423 17561 7435 17595
rect 9048 17592 9076 17623
rect 10410 17620 10416 17672
rect 10468 17620 10474 17672
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17660 12863 17663
rect 12894 17660 12900 17672
rect 12851 17632 12900 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 9214 17592 9220 17604
rect 9048 17564 9220 17592
rect 7377 17555 7435 17561
rect 9214 17552 9220 17564
rect 9272 17552 9278 17604
rect 9306 17552 9312 17604
rect 9364 17552 9370 17604
rect 4785 17527 4843 17533
rect 4785 17493 4797 17527
rect 4831 17524 4843 17527
rect 4890 17524 4896 17536
rect 4831 17496 4896 17524
rect 4831 17493 4843 17496
rect 4785 17487 4843 17493
rect 4890 17484 4896 17496
rect 4948 17524 4954 17536
rect 5258 17524 5264 17536
rect 4948 17496 5264 17524
rect 4948 17484 4954 17496
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 7064 17496 7113 17524
rect 7064 17484 7070 17496
rect 7101 17493 7113 17496
rect 7147 17524 7159 17527
rect 7650 17524 7656 17536
rect 7147 17496 7656 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 10428 17524 10456 17620
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 11790 17552 11796 17604
rect 11848 17552 11854 17604
rect 8168 17496 10456 17524
rect 8168 17484 8174 17496
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 12820 17524 12848 17623
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 13004 17669 13032 17768
rect 25608 17768 26792 17796
rect 25608 17740 25636 17768
rect 26786 17756 26792 17768
rect 26844 17756 26850 17808
rect 28258 17756 28264 17808
rect 28316 17796 28322 17808
rect 30282 17796 30288 17808
rect 28316 17768 30288 17796
rect 28316 17756 28322 17768
rect 30282 17756 30288 17768
rect 30340 17756 30346 17808
rect 31726 17796 31754 17836
rect 30392 17768 31754 17796
rect 33152 17796 33180 17836
rect 33226 17824 33232 17876
rect 33284 17824 33290 17876
rect 33318 17824 33324 17876
rect 33376 17864 33382 17876
rect 33505 17867 33563 17873
rect 33505 17864 33517 17867
rect 33376 17836 33517 17864
rect 33376 17824 33382 17836
rect 33505 17833 33517 17836
rect 33551 17833 33563 17867
rect 33505 17827 33563 17833
rect 33594 17824 33600 17876
rect 33652 17864 33658 17876
rect 34149 17867 34207 17873
rect 34149 17864 34161 17867
rect 33652 17836 34161 17864
rect 33652 17824 33658 17836
rect 34149 17833 34161 17836
rect 34195 17833 34207 17867
rect 34149 17827 34207 17833
rect 37090 17824 37096 17876
rect 37148 17864 37154 17876
rect 37231 17867 37289 17873
rect 37231 17864 37243 17867
rect 37148 17836 37243 17864
rect 37148 17824 37154 17836
rect 37231 17833 37243 17836
rect 37277 17833 37289 17867
rect 37231 17827 37289 17833
rect 34514 17796 34520 17808
rect 33152 17768 34520 17796
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17728 13415 17731
rect 13814 17728 13820 17740
rect 13403 17700 13820 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 14093 17731 14151 17737
rect 14093 17697 14105 17731
rect 14139 17728 14151 17731
rect 14734 17728 14740 17740
rect 14139 17700 14740 17728
rect 14139 17697 14151 17700
rect 14093 17691 14151 17697
rect 14734 17688 14740 17700
rect 14792 17728 14798 17740
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 14792 17700 16681 17728
rect 14792 17688 14798 17700
rect 16669 17697 16681 17700
rect 16715 17728 16727 17731
rect 17954 17728 17960 17740
rect 16715 17700 17960 17728
rect 16715 17697 16727 17700
rect 16669 17691 16727 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 19484 17700 21281 17728
rect 19484 17688 19490 17700
rect 21269 17697 21281 17700
rect 21315 17697 21327 17731
rect 21269 17691 21327 17697
rect 23017 17731 23075 17737
rect 23017 17697 23029 17731
rect 23063 17728 23075 17731
rect 23566 17728 23572 17740
rect 23063 17700 23572 17728
rect 23063 17697 23075 17700
rect 23017 17691 23075 17697
rect 23566 17688 23572 17700
rect 23624 17728 23630 17740
rect 23661 17731 23719 17737
rect 23661 17728 23673 17731
rect 23624 17700 23673 17728
rect 23624 17688 23630 17700
rect 23661 17697 23673 17700
rect 23707 17697 23719 17731
rect 25590 17728 25596 17740
rect 23661 17691 23719 17697
rect 24136 17700 25596 17728
rect 24136 17672 24164 17700
rect 25590 17688 25596 17700
rect 25648 17688 25654 17740
rect 30392 17728 30420 17768
rect 34514 17756 34520 17768
rect 34572 17756 34578 17808
rect 32122 17728 32128 17740
rect 26621 17700 27292 17728
rect 26621 17672 26649 17700
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17629 13047 17663
rect 12989 17623 13047 17629
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17660 13507 17663
rect 13538 17660 13544 17672
rect 13495 17632 13544 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 13004 17592 13032 17623
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18748 17632 19257 17660
rect 18748 17620 18754 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19610 17620 19616 17672
rect 19668 17620 19674 17672
rect 23934 17620 23940 17672
rect 23992 17620 23998 17672
rect 24029 17663 24087 17669
rect 24029 17629 24041 17663
rect 24075 17660 24087 17663
rect 24118 17660 24124 17672
rect 24075 17632 24124 17660
rect 24075 17629 24087 17632
rect 24029 17623 24087 17629
rect 24118 17620 24124 17632
rect 24176 17620 24182 17672
rect 24762 17620 24768 17672
rect 24820 17620 24826 17672
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17629 24915 17663
rect 24857 17623 24915 17629
rect 24949 17663 25007 17669
rect 24949 17629 24961 17663
rect 24995 17629 25007 17663
rect 24949 17623 25007 17629
rect 25133 17663 25191 17669
rect 25133 17629 25145 17663
rect 25179 17660 25191 17663
rect 25222 17660 25228 17672
rect 25179 17632 25228 17660
rect 25179 17629 25191 17632
rect 25133 17623 25191 17629
rect 13078 17592 13084 17604
rect 13004 17564 13084 17592
rect 13078 17552 13084 17564
rect 13136 17592 13142 17604
rect 13998 17592 14004 17604
rect 13136 17564 14004 17592
rect 13136 17552 13142 17564
rect 13998 17552 14004 17564
rect 14056 17552 14062 17604
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17561 14427 17595
rect 14369 17555 14427 17561
rect 10928 17496 12848 17524
rect 13541 17527 13599 17533
rect 10928 17484 10934 17496
rect 13541 17493 13553 17527
rect 13587 17524 13599 17527
rect 13722 17524 13728 17536
rect 13587 17496 13728 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 13909 17527 13967 17533
rect 13909 17493 13921 17527
rect 13955 17524 13967 17527
rect 14384 17524 14412 17555
rect 16942 17552 16948 17604
rect 17000 17552 17006 17604
rect 17236 17564 17434 17592
rect 13955 17496 14412 17524
rect 13955 17493 13967 17496
rect 13909 17487 13967 17493
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 17236 17524 17264 17564
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19429 17595 19487 17601
rect 19429 17592 19441 17595
rect 19392 17564 19441 17592
rect 19392 17552 19398 17564
rect 19429 17561 19441 17564
rect 19475 17561 19487 17595
rect 19429 17555 19487 17561
rect 19521 17595 19579 17601
rect 19521 17561 19533 17595
rect 19567 17592 19579 17595
rect 21266 17592 21272 17604
rect 19567 17564 21272 17592
rect 19567 17561 19579 17564
rect 19521 17555 19579 17561
rect 21266 17552 21272 17564
rect 21324 17552 21330 17604
rect 21542 17552 21548 17604
rect 21600 17552 21606 17604
rect 22094 17552 22100 17604
rect 22152 17552 22158 17604
rect 22830 17552 22836 17604
rect 22888 17592 22894 17604
rect 23109 17595 23167 17601
rect 23109 17592 23121 17595
rect 22888 17564 23121 17592
rect 22888 17552 22894 17564
rect 23109 17561 23121 17564
rect 23155 17561 23167 17595
rect 23109 17555 23167 17561
rect 23842 17552 23848 17604
rect 23900 17592 23906 17604
rect 24213 17595 24271 17601
rect 24213 17592 24225 17595
rect 23900 17564 24225 17592
rect 23900 17552 23906 17564
rect 24213 17561 24225 17564
rect 24259 17592 24271 17595
rect 24486 17592 24492 17604
rect 24259 17564 24492 17592
rect 24259 17561 24271 17564
rect 24213 17555 24271 17561
rect 24486 17552 24492 17564
rect 24544 17592 24550 17604
rect 24872 17592 24900 17623
rect 24544 17564 24900 17592
rect 24544 17552 24550 17564
rect 17954 17524 17960 17536
rect 16172 17496 17960 17524
rect 16172 17484 16178 17496
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 23750 17484 23756 17536
rect 23808 17524 23814 17536
rect 24118 17524 24124 17536
rect 23808 17496 24124 17524
rect 23808 17484 23814 17496
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 24964 17524 24992 17623
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 25498 17620 25504 17672
rect 25556 17660 25562 17672
rect 25961 17663 26019 17669
rect 25961 17660 25973 17663
rect 25556 17632 25973 17660
rect 25556 17620 25562 17632
rect 25961 17629 25973 17632
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 26142 17620 26148 17672
rect 26200 17620 26206 17672
rect 26602 17620 26608 17672
rect 26660 17620 26666 17672
rect 26786 17620 26792 17672
rect 26844 17660 26850 17672
rect 27264 17669 27292 17700
rect 28184 17700 29040 17728
rect 28184 17672 28212 17700
rect 29012 17672 29040 17700
rect 30024 17700 30420 17728
rect 30484 17700 32128 17728
rect 30024 17672 30052 17700
rect 27065 17663 27123 17669
rect 27065 17660 27077 17663
rect 26844 17632 27077 17660
rect 26844 17620 26850 17632
rect 27065 17629 27077 17632
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 27249 17663 27307 17669
rect 27249 17629 27261 17663
rect 27295 17629 27307 17663
rect 27249 17623 27307 17629
rect 27798 17620 27804 17672
rect 27856 17660 27862 17672
rect 27893 17663 27951 17669
rect 27893 17660 27905 17663
rect 27856 17632 27905 17660
rect 27856 17620 27862 17632
rect 27893 17629 27905 17632
rect 27939 17629 27951 17663
rect 27893 17623 27951 17629
rect 27982 17620 27988 17672
rect 28040 17660 28046 17672
rect 28077 17663 28135 17669
rect 28077 17660 28089 17663
rect 28040 17632 28089 17660
rect 28040 17620 28046 17632
rect 28077 17629 28089 17632
rect 28123 17629 28135 17663
rect 28077 17623 28135 17629
rect 28166 17620 28172 17672
rect 28224 17620 28230 17672
rect 28258 17620 28264 17672
rect 28316 17620 28322 17672
rect 28445 17663 28503 17669
rect 28445 17629 28457 17663
rect 28491 17629 28503 17663
rect 28445 17623 28503 17629
rect 26421 17595 26479 17601
rect 26421 17561 26433 17595
rect 26467 17561 26479 17595
rect 26421 17555 26479 17561
rect 26513 17595 26571 17601
rect 26513 17561 26525 17595
rect 26559 17592 26571 17595
rect 26973 17595 27031 17601
rect 26973 17592 26985 17595
rect 26559 17564 26985 17592
rect 26559 17561 26571 17564
rect 26513 17555 26571 17561
rect 26973 17561 26985 17564
rect 27019 17592 27031 17595
rect 28350 17592 28356 17604
rect 27019 17564 28356 17592
rect 27019 17561 27031 17564
rect 26973 17555 27031 17561
rect 24912 17496 24992 17524
rect 26436 17524 26464 17555
rect 28350 17552 28356 17564
rect 28408 17552 28414 17604
rect 28460 17592 28488 17623
rect 28718 17620 28724 17672
rect 28776 17620 28782 17672
rect 28902 17620 28908 17672
rect 28960 17620 28966 17672
rect 28994 17620 29000 17672
rect 29052 17620 29058 17672
rect 29086 17620 29092 17672
rect 29144 17660 29150 17672
rect 29638 17660 29644 17672
rect 29144 17632 29644 17660
rect 29144 17620 29150 17632
rect 29638 17620 29644 17632
rect 29696 17620 29702 17672
rect 30006 17620 30012 17672
rect 30064 17620 30070 17672
rect 30190 17620 30196 17672
rect 30248 17620 30254 17672
rect 30285 17663 30343 17669
rect 30285 17629 30297 17663
rect 30331 17629 30343 17663
rect 30285 17623 30343 17629
rect 29178 17592 29184 17604
rect 28460 17564 29184 17592
rect 29178 17552 29184 17564
rect 29236 17552 29242 17604
rect 30300 17592 30328 17623
rect 30374 17620 30380 17672
rect 30432 17660 30438 17672
rect 30484 17660 30512 17700
rect 32122 17688 32128 17700
rect 32180 17688 32186 17740
rect 32214 17688 32220 17740
rect 32272 17688 32278 17740
rect 32306 17688 32312 17740
rect 32364 17728 32370 17740
rect 34790 17728 34796 17740
rect 32364 17700 34796 17728
rect 32364 17688 32370 17700
rect 34790 17688 34796 17700
rect 34848 17688 34854 17740
rect 35802 17688 35808 17740
rect 35860 17688 35866 17740
rect 30432 17632 30512 17660
rect 30561 17663 30619 17669
rect 30432 17620 30438 17632
rect 30561 17629 30573 17663
rect 30607 17660 30619 17663
rect 30650 17660 30656 17672
rect 30607 17632 30656 17660
rect 30607 17629 30619 17632
rect 30561 17623 30619 17629
rect 30650 17620 30656 17632
rect 30708 17620 30714 17672
rect 30837 17663 30895 17669
rect 30837 17629 30849 17663
rect 30883 17629 30895 17663
rect 30837 17623 30895 17629
rect 30852 17592 30880 17623
rect 30926 17620 30932 17672
rect 30984 17660 30990 17672
rect 31662 17660 31668 17672
rect 30984 17632 31668 17660
rect 30984 17620 30990 17632
rect 31662 17620 31668 17632
rect 31720 17660 31726 17672
rect 31849 17663 31907 17669
rect 31849 17660 31861 17663
rect 31720 17632 31861 17660
rect 31720 17620 31726 17632
rect 31849 17629 31861 17632
rect 31895 17629 31907 17663
rect 31849 17623 31907 17629
rect 32030 17620 32036 17672
rect 32088 17620 32094 17672
rect 30208 17564 30880 17592
rect 30208 17536 30236 17564
rect 31018 17552 31024 17604
rect 31076 17592 31082 17604
rect 32232 17592 32260 17688
rect 32398 17620 32404 17672
rect 32456 17620 32462 17672
rect 32490 17620 32496 17672
rect 32548 17660 32554 17672
rect 32802 17663 32860 17669
rect 32802 17660 32814 17663
rect 32548 17632 32814 17660
rect 32548 17620 32554 17632
rect 32802 17629 32814 17632
rect 32848 17629 32860 17663
rect 32802 17623 32860 17629
rect 33318 17620 33324 17672
rect 33376 17620 33382 17672
rect 33689 17663 33747 17669
rect 33689 17629 33701 17663
rect 33735 17629 33747 17663
rect 33689 17623 33747 17629
rect 34333 17663 34391 17669
rect 34333 17629 34345 17663
rect 34379 17660 34391 17663
rect 34422 17660 34428 17672
rect 34379 17632 34428 17660
rect 34379 17629 34391 17632
rect 34333 17623 34391 17629
rect 31076 17564 32260 17592
rect 32585 17595 32643 17601
rect 31076 17552 31082 17564
rect 32585 17561 32597 17595
rect 32631 17592 32643 17595
rect 32631 17564 32904 17592
rect 32631 17561 32643 17564
rect 32585 17555 32643 17561
rect 26878 17524 26884 17536
rect 26436 17496 26884 17524
rect 24912 17484 24918 17496
rect 26878 17484 26884 17496
rect 26936 17484 26942 17536
rect 28258 17484 28264 17536
rect 28316 17524 28322 17536
rect 28629 17527 28687 17533
rect 28629 17524 28641 17527
rect 28316 17496 28641 17524
rect 28316 17484 28322 17496
rect 28629 17493 28641 17496
rect 28675 17493 28687 17527
rect 28629 17487 28687 17493
rect 29273 17527 29331 17533
rect 29273 17493 29285 17527
rect 29319 17524 29331 17527
rect 29454 17524 29460 17536
rect 29319 17496 29460 17524
rect 29319 17493 29331 17496
rect 29273 17487 29331 17493
rect 29454 17484 29460 17496
rect 29512 17484 29518 17536
rect 30190 17484 30196 17536
rect 30248 17484 30254 17536
rect 30558 17484 30564 17536
rect 30616 17524 30622 17536
rect 30745 17527 30803 17533
rect 30745 17524 30757 17527
rect 30616 17496 30757 17524
rect 30616 17484 30622 17496
rect 30745 17493 30757 17496
rect 30791 17493 30803 17527
rect 30745 17487 30803 17493
rect 32674 17484 32680 17536
rect 32732 17484 32738 17536
rect 32876 17533 32904 17564
rect 32861 17527 32919 17533
rect 32861 17493 32873 17527
rect 32907 17493 32919 17527
rect 33704 17524 33732 17623
rect 34422 17620 34428 17632
rect 34480 17620 34486 17672
rect 34606 17620 34612 17672
rect 34664 17660 34670 17672
rect 35437 17663 35495 17669
rect 35437 17660 35449 17663
rect 34664 17632 35449 17660
rect 34664 17620 34670 17632
rect 35437 17629 35449 17632
rect 35483 17629 35495 17663
rect 35437 17623 35495 17629
rect 34517 17595 34575 17601
rect 34517 17561 34529 17595
rect 34563 17592 34575 17595
rect 34698 17592 34704 17604
rect 34563 17564 34704 17592
rect 34563 17561 34575 17564
rect 34517 17555 34575 17561
rect 34698 17552 34704 17564
rect 34756 17552 34762 17604
rect 36170 17552 36176 17604
rect 36228 17552 36234 17604
rect 34790 17524 34796 17536
rect 33704 17496 34796 17524
rect 32861 17487 32919 17493
rect 34790 17484 34796 17496
rect 34848 17524 34854 17536
rect 37642 17524 37648 17536
rect 34848 17496 37648 17524
rect 34848 17484 34854 17496
rect 37642 17484 37648 17496
rect 37700 17484 37706 17536
rect 1104 17434 38824 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 38824 17434
rect 1104 17360 38824 17382
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5442 17320 5448 17332
rect 5316 17292 5448 17320
rect 5316 17280 5322 17292
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 7834 17320 7840 17332
rect 7699 17292 7840 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 9364 17292 10425 17320
rect 9364 17280 9370 17292
rect 10413 17289 10425 17292
rect 10459 17289 10471 17323
rect 10413 17283 10471 17289
rect 10870 17280 10876 17332
rect 10928 17280 10934 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 11204 17292 11529 17320
rect 11204 17280 11210 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 11974 17280 11980 17332
rect 12032 17280 12038 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 13630 17320 13636 17332
rect 13219 17292 13636 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 13814 17280 13820 17332
rect 13872 17280 13878 17332
rect 14550 17280 14556 17332
rect 14608 17320 14614 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14608 17292 15117 17320
rect 14608 17280 14614 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 15105 17283 15163 17289
rect 21542 17280 21548 17332
rect 21600 17320 21606 17332
rect 22005 17323 22063 17329
rect 22005 17320 22017 17323
rect 21600 17292 22017 17320
rect 21600 17280 21606 17292
rect 22005 17289 22017 17292
rect 22051 17289 22063 17323
rect 22005 17283 22063 17289
rect 22373 17323 22431 17329
rect 22373 17289 22385 17323
rect 22419 17320 22431 17323
rect 22830 17320 22836 17332
rect 22419 17292 22836 17320
rect 22419 17289 22431 17292
rect 22373 17283 22431 17289
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 23661 17323 23719 17329
rect 23661 17289 23673 17323
rect 23707 17320 23719 17323
rect 24854 17320 24860 17332
rect 23707 17292 24860 17320
rect 23707 17289 23719 17292
rect 23661 17283 23719 17289
rect 24854 17280 24860 17292
rect 24912 17280 24918 17332
rect 24946 17280 24952 17332
rect 25004 17280 25010 17332
rect 25869 17323 25927 17329
rect 25869 17289 25881 17323
rect 25915 17320 25927 17323
rect 26602 17320 26608 17332
rect 25915 17292 26608 17320
rect 25915 17289 25927 17292
rect 25869 17283 25927 17289
rect 26602 17280 26608 17292
rect 26660 17280 26666 17332
rect 27709 17323 27767 17329
rect 27709 17289 27721 17323
rect 27755 17320 27767 17323
rect 28166 17320 28172 17332
rect 27755 17292 28172 17320
rect 27755 17289 27767 17292
rect 27709 17283 27767 17289
rect 28166 17280 28172 17292
rect 28224 17280 28230 17332
rect 28350 17280 28356 17332
rect 28408 17320 28414 17332
rect 29914 17320 29920 17332
rect 28408 17292 29920 17320
rect 28408 17280 28414 17292
rect 29914 17280 29920 17292
rect 29972 17280 29978 17332
rect 30116 17292 32352 17320
rect 2777 17255 2835 17261
rect 2777 17221 2789 17255
rect 2823 17252 2835 17255
rect 3234 17252 3240 17264
rect 2823 17224 3240 17252
rect 2823 17221 2835 17224
rect 2777 17215 2835 17221
rect 3234 17212 3240 17224
rect 3292 17252 3298 17264
rect 3878 17252 3884 17264
rect 3292 17224 3884 17252
rect 3292 17212 3298 17224
rect 3878 17212 3884 17224
rect 3936 17212 3942 17264
rect 4430 17212 4436 17264
rect 4488 17212 4494 17264
rect 8110 17212 8116 17264
rect 8168 17212 8174 17264
rect 9122 17212 9128 17264
rect 9180 17212 9186 17264
rect 9214 17212 9220 17264
rect 9272 17252 9278 17264
rect 10781 17255 10839 17261
rect 9272 17224 9444 17252
rect 9272 17212 9278 17224
rect 2225 17187 2283 17193
rect 2225 17153 2237 17187
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17184 2467 17187
rect 2498 17184 2504 17196
rect 2455 17156 2504 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 2240 17116 2268 17147
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17184 2651 17187
rect 2639 17156 2774 17184
rect 2639 17153 2651 17156
rect 2593 17147 2651 17153
rect 2608 17116 2636 17147
rect 2240 17088 2636 17116
rect 2746 17116 2774 17156
rect 4062 17144 4068 17196
rect 4120 17144 4126 17196
rect 4893 17187 4951 17193
rect 4893 17153 4905 17187
rect 4939 17184 4951 17187
rect 5718 17184 5724 17196
rect 4939 17156 5724 17184
rect 4939 17153 4951 17156
rect 4893 17147 4951 17153
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 9416 17193 9444 17224
rect 10781 17221 10793 17255
rect 10827 17252 10839 17255
rect 11992 17252 12020 17280
rect 10827 17224 12020 17252
rect 10827 17221 10839 17224
rect 10781 17215 10839 17221
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 9401 17187 9459 17193
rect 6871 17156 6960 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 3142 17116 3148 17128
rect 2746 17088 3148 17116
rect 3142 17076 3148 17088
rect 3200 17116 3206 17128
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 3200 17088 3433 17116
rect 3200 17076 3206 17088
rect 3421 17085 3433 17088
rect 3467 17116 3479 17119
rect 3786 17116 3792 17128
rect 3467 17088 3792 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 3786 17076 3792 17088
rect 3844 17076 3850 17128
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 5350 17116 5356 17128
rect 4847 17088 5356 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 5902 17116 5908 17128
rect 5460 17088 5908 17116
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 5460 17048 5488 17088
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 3016 17020 5488 17048
rect 3016 17008 3022 17020
rect 2406 16940 2412 16992
rect 2464 16940 2470 16992
rect 2774 16940 2780 16992
rect 2832 16940 2838 16992
rect 2866 16940 2872 16992
rect 2924 16940 2930 16992
rect 4522 16940 4528 16992
rect 4580 16940 4586 16992
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 5077 16983 5135 16989
rect 5077 16980 5089 16983
rect 4764 16952 5089 16980
rect 4764 16940 4770 16952
rect 5077 16949 5089 16952
rect 5123 16949 5135 16983
rect 5077 16943 5135 16949
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 5592 16952 5917 16980
rect 5592 16940 5598 16952
rect 5905 16949 5917 16952
rect 5951 16949 5963 16983
rect 5905 16943 5963 16949
rect 6730 16940 6736 16992
rect 6788 16940 6794 16992
rect 6932 16989 6960 17156
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17184 11943 17187
rect 12526 17184 12532 17196
rect 11931 17156 12532 17184
rect 11931 17153 11943 17156
rect 11885 17147 11943 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12710 17144 12716 17196
rect 12768 17144 12774 17196
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17184 13047 17187
rect 13078 17184 13084 17196
rect 13035 17156 13084 17184
rect 13035 17153 13047 17156
rect 12989 17147 13047 17153
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 7558 17076 7564 17128
rect 7616 17076 7622 17128
rect 7650 17076 7656 17128
rect 7708 17116 7714 17128
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 7708 17088 9505 17116
rect 7708 17076 7714 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 10686 17116 10692 17128
rect 9732 17088 10692 17116
rect 9732 17076 9738 17088
rect 10686 17076 10692 17088
rect 10744 17116 10750 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10744 17088 10977 17116
rect 10744 17076 10750 17088
rect 10965 17085 10977 17088
rect 11011 17116 11023 17119
rect 12069 17119 12127 17125
rect 12069 17116 12081 17119
rect 11011 17088 12081 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 12069 17085 12081 17088
rect 12115 17116 12127 17119
rect 13832 17116 13860 17280
rect 14093 17255 14151 17261
rect 14093 17221 14105 17255
rect 14139 17252 14151 17255
rect 15930 17252 15936 17264
rect 14139 17224 15936 17252
rect 14139 17221 14151 17224
rect 14093 17215 14151 17221
rect 15930 17212 15936 17224
rect 15988 17212 15994 17264
rect 18782 17212 18788 17264
rect 18840 17212 18846 17264
rect 18966 17212 18972 17264
rect 19024 17261 19030 17264
rect 19024 17255 19043 17261
rect 19031 17221 19043 17255
rect 19024 17215 19043 17221
rect 19024 17212 19030 17215
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 18414 17144 18420 17196
rect 18472 17144 18478 17196
rect 19886 17144 19892 17196
rect 19944 17144 19950 17196
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17184 22523 17187
rect 23293 17187 23351 17193
rect 23293 17184 23305 17187
rect 22511 17156 23305 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 23293 17153 23305 17156
rect 23339 17184 23351 17187
rect 23474 17184 23480 17196
rect 23339 17156 23480 17184
rect 23339 17153 23351 17156
rect 23293 17147 23351 17153
rect 23474 17144 23480 17156
rect 23532 17184 23538 17196
rect 23532 17156 23796 17184
rect 23532 17144 23538 17156
rect 12115 17088 13860 17116
rect 12115 17085 12127 17088
rect 12069 17079 12127 17085
rect 19518 17076 19524 17128
rect 19576 17076 19582 17128
rect 20162 17076 20168 17128
rect 20220 17116 20226 17128
rect 20625 17119 20683 17125
rect 20625 17116 20637 17119
rect 20220 17088 20637 17116
rect 20220 17076 20226 17088
rect 20625 17085 20637 17088
rect 20671 17085 20683 17119
rect 20625 17079 20683 17085
rect 21082 17076 21088 17128
rect 21140 17116 21146 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 21140 17088 21189 17116
rect 21140 17076 21146 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 22649 17119 22707 17125
rect 22649 17085 22661 17119
rect 22695 17116 22707 17119
rect 23198 17116 23204 17128
rect 22695 17088 23204 17116
rect 22695 17085 22707 17088
rect 22649 17079 22707 17085
rect 23198 17076 23204 17088
rect 23256 17076 23262 17128
rect 23566 17076 23572 17128
rect 23624 17116 23630 17128
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23624 17088 23673 17116
rect 23624 17076 23630 17088
rect 23661 17085 23673 17088
rect 23707 17085 23719 17119
rect 23768 17116 23796 17156
rect 23934 17144 23940 17196
rect 23992 17144 23998 17196
rect 24029 17187 24087 17193
rect 24029 17153 24041 17187
rect 24075 17153 24087 17187
rect 24029 17147 24087 17153
rect 24044 17116 24072 17147
rect 24118 17144 24124 17196
rect 24176 17184 24182 17196
rect 24213 17187 24271 17193
rect 24213 17184 24225 17187
rect 24176 17156 24225 17184
rect 24176 17144 24182 17156
rect 24213 17153 24225 17156
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 24486 17144 24492 17196
rect 24544 17144 24550 17196
rect 24762 17144 24768 17196
rect 24820 17144 24826 17196
rect 24872 17184 24900 17280
rect 24964 17252 24992 17280
rect 26620 17252 26648 17280
rect 24964 17224 26280 17252
rect 26620 17224 27568 17252
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 24872 17156 24961 17184
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 25222 17144 25228 17196
rect 25280 17144 25286 17196
rect 25406 17144 25412 17196
rect 25464 17144 25470 17196
rect 25590 17144 25596 17196
rect 25648 17144 25654 17196
rect 26252 17193 26280 17224
rect 25777 17187 25835 17193
rect 25777 17153 25789 17187
rect 25823 17153 25835 17187
rect 25777 17147 25835 17153
rect 25961 17187 26019 17193
rect 25961 17153 25973 17187
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 26237 17187 26295 17193
rect 26237 17153 26249 17187
rect 26283 17184 26295 17187
rect 26786 17184 26792 17196
rect 26283 17156 26792 17184
rect 26283 17153 26295 17156
rect 26237 17147 26295 17153
rect 23768 17088 24072 17116
rect 24780 17116 24808 17144
rect 25501 17119 25559 17125
rect 25501 17116 25513 17119
rect 24780 17088 25513 17116
rect 23661 17079 23719 17085
rect 25501 17085 25513 17088
rect 25547 17116 25559 17119
rect 25792 17116 25820 17147
rect 25547 17088 25820 17116
rect 25547 17085 25559 17088
rect 25501 17079 25559 17085
rect 10137 17051 10195 17057
rect 10137 17017 10149 17051
rect 10183 17048 10195 17051
rect 11330 17048 11336 17060
rect 10183 17020 11336 17048
rect 10183 17017 10195 17020
rect 10137 17011 10195 17017
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 19337 17051 19395 17057
rect 19337 17017 19349 17051
rect 19383 17048 19395 17051
rect 19536 17048 19564 17076
rect 19978 17048 19984 17060
rect 19383 17020 19984 17048
rect 19383 17017 19395 17020
rect 19337 17011 19395 17017
rect 19978 17008 19984 17020
rect 20036 17008 20042 17060
rect 23385 17051 23443 17057
rect 23385 17017 23397 17051
rect 23431 17048 23443 17051
rect 23845 17051 23903 17057
rect 23845 17048 23857 17051
rect 23431 17020 23857 17048
rect 23431 17017 23443 17020
rect 23385 17011 23443 17017
rect 23845 17017 23857 17020
rect 23891 17017 23903 17051
rect 23845 17011 23903 17017
rect 24581 17051 24639 17057
rect 24581 17017 24593 17051
rect 24627 17048 24639 17051
rect 25976 17048 26004 17147
rect 26786 17144 26792 17156
rect 26844 17144 26850 17196
rect 26878 17144 26884 17196
rect 26936 17184 26942 17196
rect 27540 17193 27568 17224
rect 27249 17187 27307 17193
rect 27249 17184 27261 17187
rect 26936 17156 27261 17184
rect 26936 17144 26942 17156
rect 27249 17153 27261 17156
rect 27295 17153 27307 17187
rect 27249 17147 27307 17153
rect 27525 17187 27583 17193
rect 27525 17153 27537 17187
rect 27571 17153 27583 17187
rect 27525 17147 27583 17153
rect 27709 17187 27767 17193
rect 27709 17153 27721 17187
rect 27755 17153 27767 17187
rect 28184 17184 28212 17280
rect 30116 17261 30144 17292
rect 28721 17255 28779 17261
rect 28721 17221 28733 17255
rect 28767 17252 28779 17255
rect 30101 17255 30159 17261
rect 28767 17224 29868 17252
rect 28767 17221 28779 17224
rect 28721 17215 28779 17221
rect 28905 17187 28963 17193
rect 28905 17184 28917 17187
rect 28184 17156 28917 17184
rect 27709 17147 27767 17153
rect 28905 17153 28917 17156
rect 28951 17153 28963 17187
rect 28905 17147 28963 17153
rect 26050 17076 26056 17128
rect 26108 17116 26114 17128
rect 26973 17119 27031 17125
rect 26973 17116 26985 17119
rect 26108 17088 26985 17116
rect 26108 17076 26114 17088
rect 26973 17085 26985 17088
rect 27019 17116 27031 17119
rect 27724 17116 27752 17147
rect 29086 17144 29092 17196
rect 29144 17144 29150 17196
rect 29273 17187 29331 17193
rect 29273 17153 29285 17187
rect 29319 17153 29331 17187
rect 29273 17147 29331 17153
rect 27019 17088 27752 17116
rect 27019 17085 27031 17088
rect 26973 17079 27031 17085
rect 29178 17076 29184 17128
rect 29236 17076 29242 17128
rect 29288 17116 29316 17147
rect 29454 17144 29460 17196
rect 29512 17144 29518 17196
rect 29840 17193 29868 17224
rect 30101 17221 30113 17255
rect 30147 17221 30159 17255
rect 30101 17215 30159 17221
rect 30561 17255 30619 17261
rect 30561 17221 30573 17255
rect 30607 17252 30619 17255
rect 31018 17252 31024 17264
rect 30607 17224 31024 17252
rect 30607 17221 30619 17224
rect 30561 17215 30619 17221
rect 31018 17212 31024 17224
rect 31076 17212 31082 17264
rect 32125 17255 32183 17261
rect 32125 17252 32137 17255
rect 31726 17224 32137 17252
rect 29825 17187 29883 17193
rect 29825 17153 29837 17187
rect 29871 17153 29883 17187
rect 29825 17147 29883 17153
rect 29914 17144 29920 17196
rect 29972 17184 29978 17196
rect 29972 17156 30017 17184
rect 29972 17144 29978 17156
rect 30190 17144 30196 17196
rect 30248 17144 30254 17196
rect 30282 17144 30288 17196
rect 30340 17193 30346 17196
rect 30340 17184 30348 17193
rect 30340 17156 30385 17184
rect 30340 17147 30348 17156
rect 30340 17144 30346 17147
rect 30650 17144 30656 17196
rect 30708 17144 30714 17196
rect 30929 17187 30987 17193
rect 30929 17153 30941 17187
rect 30975 17184 30987 17187
rect 31205 17187 31263 17193
rect 30975 17156 31156 17184
rect 30975 17153 30987 17156
rect 30929 17147 30987 17153
rect 30208 17116 30236 17144
rect 31021 17119 31079 17125
rect 31021 17116 31033 17119
rect 29288 17088 30236 17116
rect 30484 17088 31033 17116
rect 26142 17048 26148 17060
rect 24627 17020 26148 17048
rect 24627 17017 24639 17020
rect 24581 17011 24639 17017
rect 26142 17008 26148 17020
rect 26200 17048 26206 17060
rect 27065 17051 27123 17057
rect 27065 17048 27077 17051
rect 26200 17020 27077 17048
rect 26200 17008 26206 17020
rect 27065 17017 27077 17020
rect 27111 17017 27123 17051
rect 27065 17011 27123 17017
rect 27433 17051 27491 17057
rect 27433 17017 27445 17051
rect 27479 17048 27491 17051
rect 29288 17048 29316 17088
rect 30484 17057 30512 17088
rect 31021 17085 31033 17088
rect 31067 17085 31079 17119
rect 31128 17116 31156 17156
rect 31205 17153 31217 17187
rect 31251 17184 31263 17187
rect 31726 17184 31754 17224
rect 32125 17221 32137 17224
rect 32171 17221 32183 17255
rect 32324 17252 32352 17292
rect 32398 17280 32404 17332
rect 32456 17320 32462 17332
rect 32953 17323 33011 17329
rect 32953 17320 32965 17323
rect 32456 17292 32965 17320
rect 32456 17280 32462 17292
rect 32953 17289 32965 17292
rect 32999 17289 33011 17323
rect 36357 17323 36415 17329
rect 32953 17283 33011 17289
rect 33152 17292 33824 17320
rect 32490 17252 32496 17264
rect 32324 17224 32496 17252
rect 32125 17215 32183 17221
rect 32490 17212 32496 17224
rect 32548 17252 32554 17264
rect 33152 17252 33180 17292
rect 33796 17261 33824 17292
rect 36357 17289 36369 17323
rect 36403 17320 36415 17323
rect 36630 17320 36636 17332
rect 36403 17292 36636 17320
rect 36403 17289 36415 17292
rect 36357 17283 36415 17289
rect 36630 17280 36636 17292
rect 36688 17280 36694 17332
rect 32548 17224 32720 17252
rect 32548 17212 32554 17224
rect 31251 17156 31754 17184
rect 31941 17187 31999 17193
rect 31251 17153 31263 17156
rect 31205 17147 31263 17153
rect 31941 17153 31953 17187
rect 31987 17184 31999 17187
rect 32214 17184 32220 17196
rect 31987 17156 32220 17184
rect 31987 17153 31999 17156
rect 31941 17147 31999 17153
rect 32214 17144 32220 17156
rect 32272 17144 32278 17196
rect 32309 17187 32367 17193
rect 32309 17153 32321 17187
rect 32355 17184 32367 17187
rect 32355 17156 32444 17184
rect 32355 17153 32367 17156
rect 32309 17147 32367 17153
rect 31128 17088 31432 17116
rect 31021 17079 31079 17085
rect 27479 17020 29316 17048
rect 30469 17051 30527 17057
rect 27479 17017 27491 17020
rect 27433 17011 27491 17017
rect 30469 17017 30481 17051
rect 30515 17017 30527 17051
rect 30469 17011 30527 17017
rect 31404 16992 31432 17088
rect 6917 16983 6975 16989
rect 6917 16949 6929 16983
rect 6963 16980 6975 16983
rect 9766 16980 9772 16992
rect 6963 16952 9772 16980
rect 6963 16949 6975 16952
rect 6917 16943 6975 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 18230 16980 18236 16992
rect 15988 16952 18236 16980
rect 15988 16940 15994 16952
rect 18230 16940 18236 16952
rect 18288 16980 18294 16992
rect 18601 16983 18659 16989
rect 18601 16980 18613 16983
rect 18288 16952 18613 16980
rect 18288 16940 18294 16952
rect 18601 16949 18613 16952
rect 18647 16949 18659 16983
rect 18601 16943 18659 16949
rect 18690 16940 18696 16992
rect 18748 16980 18754 16992
rect 18969 16983 19027 16989
rect 18969 16980 18981 16983
rect 18748 16952 18981 16980
rect 18748 16940 18754 16952
rect 18969 16949 18981 16952
rect 19015 16949 19027 16983
rect 18969 16943 19027 16949
rect 19150 16940 19156 16992
rect 19208 16940 19214 16992
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 19705 16983 19763 16989
rect 19705 16980 19717 16983
rect 19576 16952 19717 16980
rect 19576 16940 19582 16952
rect 19705 16949 19717 16952
rect 19751 16949 19763 16983
rect 19705 16943 19763 16949
rect 20073 16983 20131 16989
rect 20073 16949 20085 16983
rect 20119 16980 20131 16983
rect 20254 16980 20260 16992
rect 20119 16952 20260 16980
rect 20119 16949 20131 16952
rect 20073 16943 20131 16949
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 24397 16983 24455 16989
rect 24397 16949 24409 16983
rect 24443 16980 24455 16983
rect 24854 16980 24860 16992
rect 24443 16952 24860 16980
rect 24443 16949 24455 16952
rect 24397 16943 24455 16949
rect 24854 16940 24860 16952
rect 24912 16940 24918 16992
rect 25866 16940 25872 16992
rect 25924 16980 25930 16992
rect 30006 16980 30012 16992
rect 25924 16952 30012 16980
rect 25924 16940 25930 16952
rect 30006 16940 30012 16952
rect 30064 16940 30070 16992
rect 30098 16940 30104 16992
rect 30156 16980 30162 16992
rect 31294 16980 31300 16992
rect 30156 16952 31300 16980
rect 30156 16940 30162 16952
rect 31294 16940 31300 16952
rect 31352 16940 31358 16992
rect 31386 16940 31392 16992
rect 31444 16940 31450 16992
rect 31754 16940 31760 16992
rect 31812 16940 31818 16992
rect 32416 16980 32444 17156
rect 32582 17144 32588 17196
rect 32640 17144 32646 17196
rect 32692 17193 32720 17224
rect 32876 17224 33180 17252
rect 33781 17255 33839 17261
rect 32876 17193 32904 17224
rect 33551 17221 33609 17227
rect 32677 17187 32735 17193
rect 32677 17153 32689 17187
rect 32723 17153 32735 17187
rect 32677 17147 32735 17153
rect 32861 17187 32919 17193
rect 32861 17153 32873 17187
rect 32907 17153 32919 17187
rect 32861 17147 32919 17153
rect 33134 17144 33140 17196
rect 33192 17144 33198 17196
rect 33551 17187 33563 17221
rect 33597 17187 33609 17221
rect 33781 17221 33793 17255
rect 33827 17252 33839 17255
rect 34422 17252 34428 17264
rect 33827 17224 34428 17252
rect 33827 17221 33839 17224
rect 33781 17215 33839 17221
rect 34422 17212 34428 17224
rect 34480 17212 34486 17264
rect 34517 17255 34575 17261
rect 34517 17221 34529 17255
rect 34563 17252 34575 17255
rect 34885 17255 34943 17261
rect 34885 17252 34897 17255
rect 34563 17224 34897 17252
rect 34563 17221 34575 17224
rect 34517 17215 34575 17221
rect 34885 17221 34897 17224
rect 34931 17221 34943 17255
rect 34885 17215 34943 17221
rect 33551 17184 33609 17187
rect 33336 17181 33609 17184
rect 33336 17156 33608 17181
rect 32493 17119 32551 17125
rect 32493 17085 32505 17119
rect 32539 17116 32551 17119
rect 32950 17116 32956 17128
rect 32539 17088 32956 17116
rect 32539 17085 32551 17088
rect 32493 17079 32551 17085
rect 32950 17076 32956 17088
rect 33008 17116 33014 17128
rect 33336 17125 33364 17156
rect 33686 17144 33692 17196
rect 33744 17184 33750 17196
rect 33965 17187 34023 17193
rect 33965 17184 33977 17187
rect 33744 17156 33977 17184
rect 33744 17144 33750 17156
rect 33965 17153 33977 17156
rect 34011 17153 34023 17187
rect 33965 17147 34023 17153
rect 34238 17144 34244 17196
rect 34296 17144 34302 17196
rect 34333 17187 34391 17193
rect 34333 17153 34345 17187
rect 34379 17153 34391 17187
rect 34333 17147 34391 17153
rect 33321 17119 33379 17125
rect 33321 17116 33333 17119
rect 33008 17088 33333 17116
rect 33008 17076 33014 17088
rect 33321 17085 33333 17088
rect 33367 17085 33379 17119
rect 34348 17116 34376 17147
rect 35986 17144 35992 17196
rect 36044 17144 36050 17196
rect 33321 17079 33379 17085
rect 33428 17088 34376 17116
rect 33428 17060 33456 17088
rect 34606 17076 34612 17128
rect 34664 17076 34670 17128
rect 33410 17008 33416 17060
rect 33468 17008 33474 17060
rect 34057 17051 34115 17057
rect 34057 17017 34069 17051
rect 34103 17048 34115 17051
rect 34514 17048 34520 17060
rect 34103 17020 34520 17048
rect 34103 17017 34115 17020
rect 34057 17011 34115 17017
rect 34514 17008 34520 17020
rect 34572 17008 34578 17060
rect 33597 16983 33655 16989
rect 33597 16980 33609 16983
rect 32416 16952 33609 16980
rect 33597 16949 33609 16952
rect 33643 16980 33655 16983
rect 33686 16980 33692 16992
rect 33643 16952 33692 16980
rect 33643 16949 33655 16952
rect 33597 16943 33655 16949
rect 33686 16940 33692 16952
rect 33744 16940 33750 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 3142 16736 3148 16788
rect 3200 16776 3206 16788
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 3200 16748 3433 16776
rect 3200 16736 3206 16748
rect 3421 16745 3433 16748
rect 3467 16745 3479 16779
rect 3421 16739 3479 16745
rect 7006 16736 7012 16788
rect 7064 16736 7070 16788
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 12805 16779 12863 16785
rect 12805 16776 12817 16779
rect 12768 16748 12817 16776
rect 12768 16736 12774 16748
rect 12805 16745 12817 16748
rect 12851 16745 12863 16779
rect 12805 16739 12863 16745
rect 15010 16736 15016 16788
rect 15068 16776 15074 16788
rect 15105 16779 15163 16785
rect 15105 16776 15117 16779
rect 15068 16748 15117 16776
rect 15068 16736 15074 16748
rect 15105 16745 15117 16748
rect 15151 16745 15163 16779
rect 15105 16739 15163 16745
rect 16209 16779 16267 16785
rect 16209 16745 16221 16779
rect 16255 16776 16267 16779
rect 17218 16776 17224 16788
rect 16255 16748 17224 16776
rect 16255 16745 16267 16748
rect 16209 16739 16267 16745
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17484 16779 17542 16785
rect 17484 16745 17496 16779
rect 17530 16776 17542 16779
rect 18598 16776 18604 16788
rect 17530 16748 18604 16776
rect 17530 16745 17542 16748
rect 17484 16739 17542 16745
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 18782 16736 18788 16788
rect 18840 16776 18846 16788
rect 18969 16779 19027 16785
rect 18969 16776 18981 16779
rect 18840 16748 18981 16776
rect 18840 16736 18846 16748
rect 18969 16745 18981 16748
rect 19015 16745 19027 16779
rect 18969 16739 19027 16745
rect 25133 16779 25191 16785
rect 25133 16745 25145 16779
rect 25179 16776 25191 16779
rect 25222 16776 25228 16788
rect 25179 16748 25228 16776
rect 25179 16745 25191 16748
rect 25133 16739 25191 16745
rect 25222 16736 25228 16748
rect 25280 16736 25286 16788
rect 29178 16736 29184 16788
rect 29236 16776 29242 16788
rect 29733 16779 29791 16785
rect 29733 16776 29745 16779
rect 29236 16748 29745 16776
rect 29236 16736 29242 16748
rect 29733 16745 29745 16748
rect 29779 16776 29791 16779
rect 30282 16776 30288 16788
rect 29779 16748 30288 16776
rect 29779 16745 29791 16748
rect 29733 16739 29791 16745
rect 30282 16736 30288 16748
rect 30340 16776 30346 16788
rect 32217 16779 32275 16785
rect 30340 16748 31156 16776
rect 30340 16736 30346 16748
rect 5169 16711 5227 16717
rect 5169 16677 5181 16711
rect 5215 16708 5227 16711
rect 5350 16708 5356 16720
rect 5215 16680 5356 16708
rect 5215 16677 5227 16680
rect 5169 16671 5227 16677
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 10965 16711 11023 16717
rect 10965 16708 10977 16711
rect 9600 16680 10977 16708
rect 1394 16600 1400 16652
rect 1452 16640 1458 16652
rect 4062 16640 4068 16652
rect 1452 16612 4068 16640
rect 1452 16600 1458 16612
rect 4062 16600 4068 16612
rect 4120 16640 4126 16652
rect 4249 16643 4307 16649
rect 4249 16640 4261 16643
rect 4120 16612 4261 16640
rect 4120 16600 4126 16612
rect 4249 16609 4261 16612
rect 4295 16640 4307 16643
rect 6914 16640 6920 16652
rect 4295 16612 6920 16640
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 6914 16600 6920 16612
rect 6972 16600 6978 16652
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 9600 16640 9628 16680
rect 10965 16677 10977 16680
rect 11011 16677 11023 16711
rect 15746 16708 15752 16720
rect 10965 16671 11023 16677
rect 15304 16680 15752 16708
rect 8527 16612 9628 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 9674 16600 9680 16652
rect 9732 16600 9738 16652
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 11241 16643 11299 16649
rect 11241 16640 11253 16643
rect 9824 16612 11253 16640
rect 9824 16600 9830 16612
rect 11241 16609 11253 16612
rect 11287 16609 11299 16643
rect 13722 16640 13728 16652
rect 11241 16603 11299 16609
rect 13004 16612 13728 16640
rect 8757 16575 8815 16581
rect 3068 16544 3372 16572
rect 1670 16464 1676 16516
rect 1728 16464 1734 16516
rect 2682 16464 2688 16516
rect 2740 16464 2746 16516
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 3068 16436 3096 16544
rect 3234 16464 3240 16516
rect 3292 16464 3298 16516
rect 3344 16504 3372 16544
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 9214 16572 9220 16584
rect 8803 16544 9220 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 9214 16532 9220 16544
rect 9272 16572 9278 16584
rect 10689 16575 10747 16581
rect 10689 16572 10701 16575
rect 9272 16544 10701 16572
rect 9272 16532 9278 16544
rect 10689 16541 10701 16544
rect 10735 16541 10747 16575
rect 10689 16535 10747 16541
rect 11330 16532 11336 16584
rect 11388 16532 11394 16584
rect 13004 16581 13032 16612
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 15304 16584 15332 16680
rect 15746 16668 15752 16680
rect 15804 16708 15810 16720
rect 16117 16711 16175 16717
rect 16117 16708 16129 16711
rect 15804 16680 16129 16708
rect 15804 16668 15810 16680
rect 16117 16677 16129 16680
rect 16163 16677 16175 16711
rect 16117 16671 16175 16677
rect 24854 16668 24860 16720
rect 24912 16708 24918 16720
rect 25682 16708 25688 16720
rect 24912 16680 25688 16708
rect 24912 16668 24918 16680
rect 25682 16668 25688 16680
rect 25740 16708 25746 16720
rect 26050 16708 26056 16720
rect 25740 16680 26056 16708
rect 25740 16668 25746 16680
rect 26050 16668 26056 16680
rect 26108 16668 26114 16720
rect 28626 16668 28632 16720
rect 28684 16708 28690 16720
rect 30926 16708 30932 16720
rect 28684 16680 30932 16708
rect 28684 16668 28690 16680
rect 30926 16668 30932 16680
rect 30984 16668 30990 16720
rect 15979 16643 16037 16649
rect 15979 16609 15991 16643
rect 16025 16609 16037 16643
rect 15979 16603 16037 16609
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16640 17279 16643
rect 17267 16612 19104 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 13262 16532 13268 16584
rect 13320 16532 13326 16584
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13814 16572 13820 16584
rect 13495 16544 13820 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 15286 16532 15292 16584
rect 15344 16532 15350 16584
rect 15562 16532 15568 16584
rect 15620 16532 15626 16584
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 3437 16507 3495 16513
rect 3437 16504 3449 16507
rect 3344 16476 3449 16504
rect 3437 16473 3449 16476
rect 3483 16473 3495 16507
rect 3437 16467 3495 16473
rect 4985 16507 5043 16513
rect 4985 16473 4997 16507
rect 5031 16504 5043 16507
rect 5258 16504 5264 16516
rect 5031 16476 5264 16504
rect 5031 16473 5043 16476
rect 4985 16467 5043 16473
rect 5258 16464 5264 16476
rect 5316 16464 5322 16516
rect 5902 16464 5908 16516
rect 5960 16464 5966 16516
rect 6362 16464 6368 16516
rect 6420 16504 6426 16516
rect 6641 16507 6699 16513
rect 6641 16504 6653 16507
rect 6420 16476 6653 16504
rect 6420 16464 6426 16476
rect 6641 16473 6653 16476
rect 6687 16473 6699 16507
rect 6641 16467 6699 16473
rect 6932 16476 7236 16504
rect 2556 16408 3096 16436
rect 2556 16396 2562 16408
rect 3142 16396 3148 16448
rect 3200 16396 3206 16448
rect 3605 16439 3663 16445
rect 3605 16405 3617 16439
rect 3651 16436 3663 16439
rect 4154 16436 4160 16448
rect 3651 16408 4160 16436
rect 3651 16405 3663 16408
rect 3605 16399 3663 16405
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 5276 16436 5304 16464
rect 6932 16436 6960 16476
rect 5276 16408 6960 16436
rect 7208 16436 7236 16476
rect 8018 16464 8024 16516
rect 8076 16464 8082 16516
rect 9953 16507 10011 16513
rect 9953 16504 9965 16507
rect 9048 16476 9965 16504
rect 9048 16436 9076 16476
rect 9953 16473 9965 16476
rect 9999 16473 10011 16507
rect 15764 16504 15792 16535
rect 15838 16532 15844 16584
rect 15896 16532 15902 16584
rect 15994 16504 16022 16603
rect 19076 16584 19104 16612
rect 19518 16600 19524 16652
rect 19576 16600 19582 16652
rect 20254 16600 20260 16652
rect 20312 16640 20318 16652
rect 23014 16640 23020 16652
rect 20312 16612 21128 16640
rect 20312 16600 20318 16612
rect 16298 16532 16304 16584
rect 16356 16532 16362 16584
rect 19058 16532 19064 16584
rect 19116 16572 19122 16584
rect 21100 16581 21128 16612
rect 22020 16612 23020 16640
rect 22020 16584 22048 16612
rect 23014 16600 23020 16612
rect 23072 16600 23078 16652
rect 24026 16600 24032 16652
rect 24084 16640 24090 16652
rect 25406 16640 25412 16652
rect 24084 16612 25412 16640
rect 24084 16600 24090 16612
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 19116 16544 19257 16572
rect 19116 16532 19122 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 21085 16575 21143 16581
rect 21085 16541 21097 16575
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 15764 16476 16022 16504
rect 9953 16467 10011 16473
rect 7208 16408 9076 16436
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 9493 16439 9551 16445
rect 9493 16436 9505 16439
rect 9456 16408 9505 16436
rect 9456 16396 9462 16408
rect 9493 16405 9505 16408
rect 9539 16405 9551 16439
rect 9493 16399 9551 16405
rect 9585 16439 9643 16445
rect 9585 16405 9597 16439
rect 9631 16436 9643 16439
rect 9858 16436 9864 16448
rect 9631 16408 9864 16436
rect 9631 16405 9643 16408
rect 9585 16399 9643 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 9968 16436 9996 16467
rect 15948 16448 15976 16476
rect 17954 16464 17960 16516
rect 18012 16464 18018 16516
rect 19260 16504 19288 16535
rect 22002 16532 22008 16584
rect 22060 16532 22066 16584
rect 22094 16532 22100 16584
rect 22152 16572 22158 16584
rect 22281 16575 22339 16581
rect 22281 16572 22293 16575
rect 22152 16544 22293 16572
rect 22152 16532 22158 16544
rect 22281 16541 22293 16544
rect 22327 16541 22339 16575
rect 22281 16535 22339 16541
rect 25130 16532 25136 16584
rect 25188 16532 25194 16584
rect 25332 16581 25360 16612
rect 25406 16600 25412 16612
rect 25464 16600 25470 16652
rect 26786 16600 26792 16652
rect 26844 16640 26850 16652
rect 27249 16643 27307 16649
rect 27249 16640 27261 16643
rect 26844 16612 27261 16640
rect 26844 16600 26850 16612
rect 27249 16609 27261 16612
rect 27295 16609 27307 16643
rect 27249 16603 27307 16609
rect 27525 16643 27583 16649
rect 27525 16609 27537 16643
rect 27571 16640 27583 16643
rect 28074 16640 28080 16652
rect 27571 16612 28080 16640
rect 27571 16609 27583 16612
rect 27525 16603 27583 16609
rect 28074 16600 28080 16612
rect 28132 16600 28138 16652
rect 30098 16600 30104 16652
rect 30156 16600 30162 16652
rect 31128 16649 31156 16748
rect 32217 16745 32229 16779
rect 32263 16776 32275 16779
rect 33134 16776 33140 16788
rect 32263 16748 33140 16776
rect 32263 16745 32275 16748
rect 32217 16739 32275 16745
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 34517 16779 34575 16785
rect 34517 16745 34529 16779
rect 34563 16776 34575 16779
rect 34790 16776 34796 16788
rect 34563 16748 34796 16776
rect 34563 16745 34575 16748
rect 34517 16739 34575 16745
rect 34790 16736 34796 16748
rect 34848 16736 34854 16788
rect 31294 16668 31300 16720
rect 31352 16708 31358 16720
rect 32125 16711 32183 16717
rect 32125 16708 32137 16711
rect 31352 16680 32137 16708
rect 31352 16668 31358 16680
rect 32125 16677 32137 16680
rect 32171 16677 32183 16711
rect 32125 16671 32183 16677
rect 32490 16668 32496 16720
rect 32548 16668 32554 16720
rect 31021 16643 31079 16649
rect 31021 16640 31033 16643
rect 30484 16612 31033 16640
rect 25317 16575 25375 16581
rect 25317 16541 25329 16575
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16572 30067 16575
rect 30484 16572 30512 16612
rect 31021 16609 31033 16612
rect 31067 16609 31079 16643
rect 31021 16603 31079 16609
rect 31113 16643 31171 16649
rect 31113 16609 31125 16643
rect 31159 16609 31171 16643
rect 31754 16640 31760 16652
rect 31113 16603 31171 16609
rect 31220 16612 31760 16640
rect 30055 16544 30512 16572
rect 30558 16575 30616 16581
rect 30055 16541 30067 16544
rect 30009 16535 30067 16541
rect 30558 16541 30570 16575
rect 30604 16572 30616 16575
rect 31036 16572 31064 16603
rect 31220 16572 31248 16612
rect 31754 16600 31760 16612
rect 31812 16640 31818 16652
rect 32309 16643 32367 16649
rect 31812 16612 32076 16640
rect 31812 16600 31818 16612
rect 30604 16544 30880 16572
rect 31036 16544 31248 16572
rect 31297 16575 31355 16581
rect 30604 16541 30616 16544
rect 30558 16535 30616 16541
rect 19426 16504 19432 16516
rect 19260 16476 19432 16504
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 19978 16464 19984 16516
rect 20036 16464 20042 16516
rect 22554 16464 22560 16516
rect 22612 16464 22618 16516
rect 23014 16464 23020 16516
rect 23072 16464 23078 16516
rect 23934 16464 23940 16516
rect 23992 16504 23998 16516
rect 26053 16507 26111 16513
rect 26053 16504 26065 16507
rect 23992 16476 26065 16504
rect 23992 16464 23998 16476
rect 26053 16473 26065 16476
rect 26099 16504 26111 16507
rect 27065 16507 27123 16513
rect 27065 16504 27077 16507
rect 26099 16476 27077 16504
rect 26099 16473 26111 16476
rect 26053 16467 26111 16473
rect 27065 16473 27077 16476
rect 27111 16473 27123 16507
rect 27065 16467 27123 16473
rect 11422 16436 11428 16448
rect 9968 16408 11428 16436
rect 11422 16396 11428 16408
rect 11480 16436 11486 16448
rect 11609 16439 11667 16445
rect 11609 16436 11621 16439
rect 11480 16408 11621 16436
rect 11480 16396 11486 16408
rect 11609 16405 11621 16408
rect 11655 16405 11667 16439
rect 11609 16399 11667 16405
rect 15930 16396 15936 16448
rect 15988 16396 15994 16448
rect 20993 16439 21051 16445
rect 20993 16405 21005 16439
rect 21039 16436 21051 16439
rect 21082 16436 21088 16448
rect 21039 16408 21088 16436
rect 21039 16405 21051 16408
rect 20993 16399 21051 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 21174 16396 21180 16448
rect 21232 16396 21238 16448
rect 24026 16396 24032 16448
rect 24084 16396 24090 16448
rect 27080 16436 27108 16467
rect 27982 16464 27988 16516
rect 28040 16464 28046 16516
rect 28994 16464 29000 16516
rect 29052 16504 29058 16516
rect 29273 16507 29331 16513
rect 29273 16504 29285 16507
rect 29052 16476 29285 16504
rect 29052 16464 29058 16476
rect 29273 16473 29285 16476
rect 29319 16504 29331 16507
rect 29362 16504 29368 16516
rect 29319 16476 29368 16504
rect 29319 16473 29331 16476
rect 29273 16467 29331 16473
rect 29362 16464 29368 16476
rect 29420 16464 29426 16516
rect 30852 16504 30880 16544
rect 31297 16541 31309 16575
rect 31343 16541 31355 16575
rect 31297 16535 31355 16541
rect 31113 16507 31171 16513
rect 31113 16504 31125 16507
rect 30852 16476 31125 16504
rect 31113 16473 31125 16476
rect 31159 16473 31171 16507
rect 31312 16504 31340 16535
rect 31386 16532 31392 16584
rect 31444 16532 31450 16584
rect 32048 16581 32076 16612
rect 32309 16609 32321 16643
rect 32355 16609 32367 16643
rect 32309 16603 32367 16609
rect 32033 16575 32091 16581
rect 32033 16541 32045 16575
rect 32079 16541 32091 16575
rect 32033 16535 32091 16541
rect 31113 16467 31171 16473
rect 31266 16476 31340 16504
rect 32324 16504 32352 16603
rect 32398 16600 32404 16652
rect 32456 16640 32462 16652
rect 32456 16612 32628 16640
rect 32456 16600 32462 16612
rect 32600 16581 32628 16612
rect 32674 16600 32680 16652
rect 32732 16640 32738 16652
rect 33045 16643 33103 16649
rect 33045 16640 33057 16643
rect 32732 16612 33057 16640
rect 32732 16600 32738 16612
rect 33045 16609 33057 16612
rect 33091 16609 33103 16643
rect 33045 16603 33103 16609
rect 32585 16575 32643 16581
rect 32585 16541 32597 16575
rect 32631 16541 32643 16575
rect 32585 16535 32643 16541
rect 32766 16532 32772 16584
rect 32824 16532 32830 16584
rect 33318 16504 33324 16516
rect 32324 16476 33324 16504
rect 29454 16436 29460 16448
rect 27080 16408 29460 16436
rect 29454 16396 29460 16408
rect 29512 16396 29518 16448
rect 30377 16439 30435 16445
rect 30377 16405 30389 16439
rect 30423 16436 30435 16439
rect 30466 16436 30472 16448
rect 30423 16408 30472 16436
rect 30423 16405 30435 16408
rect 30377 16399 30435 16405
rect 30466 16396 30472 16408
rect 30524 16396 30530 16448
rect 30558 16396 30564 16448
rect 30616 16396 30622 16448
rect 30650 16396 30656 16448
rect 30708 16436 30714 16448
rect 31266 16436 31294 16476
rect 33318 16464 33324 16476
rect 33376 16464 33382 16516
rect 36170 16504 36176 16516
rect 34270 16476 36176 16504
rect 30708 16408 31294 16436
rect 30708 16396 30714 16408
rect 31662 16396 31668 16448
rect 31720 16436 31726 16448
rect 34348 16436 34376 16476
rect 36170 16464 36176 16476
rect 36228 16464 36234 16516
rect 31720 16408 34376 16436
rect 31720 16396 31726 16408
rect 1104 16346 38824 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 38824 16346
rect 1104 16272 38824 16294
rect 2593 16235 2651 16241
rect 2593 16201 2605 16235
rect 2639 16232 2651 16235
rect 2866 16232 2872 16244
rect 2639 16204 2872 16232
rect 2639 16201 2651 16204
rect 2593 16195 2651 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 4154 16232 4160 16244
rect 3436 16204 4160 16232
rect 1670 16124 1676 16176
rect 1728 16164 1734 16176
rect 2225 16167 2283 16173
rect 2225 16164 2237 16167
rect 1728 16136 2237 16164
rect 1728 16124 1734 16136
rect 2225 16133 2237 16136
rect 2271 16133 2283 16167
rect 2225 16127 2283 16133
rect 2498 16124 2504 16176
rect 2556 16164 2562 16176
rect 2685 16167 2743 16173
rect 2685 16164 2697 16167
rect 2556 16136 2697 16164
rect 2556 16124 2562 16136
rect 2685 16133 2697 16136
rect 2731 16133 2743 16167
rect 2685 16127 2743 16133
rect 2406 16056 2412 16108
rect 2464 16056 2470 16108
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 3436 16105 3464 16204
rect 4154 16192 4160 16204
rect 4212 16232 4218 16244
rect 5442 16232 5448 16244
rect 4212 16204 5448 16232
rect 4212 16192 4218 16204
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 7616 16204 8309 16232
rect 7616 16192 7622 16204
rect 8297 16201 8309 16204
rect 8343 16201 8355 16235
rect 8297 16195 8355 16201
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 9456 16204 10977 16232
rect 9456 16192 9462 16204
rect 10965 16201 10977 16204
rect 11011 16232 11023 16235
rect 11330 16232 11336 16244
rect 11011 16204 11336 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11330 16192 11336 16204
rect 11388 16232 11394 16244
rect 13633 16235 13691 16241
rect 11388 16204 12434 16232
rect 11388 16192 11394 16204
rect 4062 16164 4068 16176
rect 3528 16136 4068 16164
rect 3528 16105 3556 16136
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 3329 16099 3387 16105
rect 3329 16096 3341 16099
rect 2832 16068 3341 16096
rect 2832 16056 2838 16068
rect 3329 16065 3341 16068
rect 3375 16065 3387 16099
rect 3329 16059 3387 16065
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 3513 16099 3571 16105
rect 3513 16065 3525 16099
rect 3559 16065 3571 16099
rect 5074 16096 5080 16108
rect 4922 16068 5080 16096
rect 3513 16059 3571 16065
rect 5074 16056 5080 16068
rect 5132 16096 5138 16108
rect 5132 16068 5396 16096
rect 5132 16056 5138 16068
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 16028 2375 16031
rect 2958 16028 2964 16040
rect 2363 16000 2964 16028
rect 2363 15997 2375 16000
rect 2317 15991 2375 15997
rect 2958 15988 2964 16000
rect 3016 16028 3022 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 3016 16000 3157 16028
rect 3016 15988 3022 16000
rect 3145 15997 3157 16000
rect 3191 15997 3203 16031
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3145 15991 3203 15997
rect 3436 16000 3801 16028
rect 3436 15969 3464 16000
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15929 3479 15963
rect 3421 15923 3479 15929
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 4890 15892 4896 15904
rect 3292 15864 4896 15892
rect 3292 15852 3298 15864
rect 4890 15852 4896 15864
rect 4948 15892 4954 15904
rect 5261 15895 5319 15901
rect 5261 15892 5273 15895
rect 4948 15864 5273 15892
rect 4948 15852 4954 15864
rect 5261 15861 5273 15864
rect 5307 15861 5319 15895
rect 5368 15892 5396 16068
rect 5460 16037 5488 16192
rect 6822 16164 6828 16176
rect 6564 16136 6828 16164
rect 5534 16056 5540 16108
rect 5592 16056 5598 16108
rect 6564 16105 6592 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 9122 16124 9128 16176
rect 9180 16164 9186 16176
rect 9493 16167 9551 16173
rect 9493 16164 9505 16167
rect 9180 16136 9505 16164
rect 9180 16124 9186 16136
rect 9493 16133 9505 16136
rect 9539 16133 9551 16167
rect 9493 16127 9551 16133
rect 10042 16124 10048 16176
rect 10100 16124 10106 16176
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 7926 16056 7932 16108
rect 7984 16056 7990 16108
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 8527 16068 8800 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 15997 5503 16031
rect 5445 15991 5503 15997
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 6362 16028 6368 16040
rect 5951 16000 6368 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6362 15988 6368 16000
rect 6420 15988 6426 16040
rect 6822 15988 6828 16040
rect 6880 15988 6886 16040
rect 7944 16028 7972 16056
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 7944 16000 8677 16028
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 8665 15991 8723 15997
rect 8772 15892 8800 16068
rect 9214 15988 9220 16040
rect 9272 15988 9278 16040
rect 5368 15864 8800 15892
rect 12406 15892 12434 16204
rect 13633 16201 13645 16235
rect 13679 16232 13691 16235
rect 15286 16232 15292 16244
rect 13679 16204 15292 16232
rect 13679 16201 13691 16204
rect 13633 16195 13691 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 15562 16192 15568 16244
rect 15620 16192 15626 16244
rect 17310 16192 17316 16244
rect 17368 16192 17374 16244
rect 18598 16192 18604 16244
rect 18656 16192 18662 16244
rect 19886 16192 19892 16244
rect 19944 16232 19950 16244
rect 20073 16235 20131 16241
rect 20073 16232 20085 16235
rect 19944 16204 20085 16232
rect 19944 16192 19950 16204
rect 20073 16201 20085 16204
rect 20119 16201 20131 16235
rect 20073 16195 20131 16201
rect 20162 16192 20168 16244
rect 20220 16192 20226 16244
rect 20559 16235 20617 16241
rect 20559 16201 20571 16235
rect 20605 16232 20617 16235
rect 21174 16232 21180 16244
rect 20605 16204 21180 16232
rect 20605 16201 20617 16204
rect 20559 16195 20617 16201
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22612 16204 23029 16232
rect 22612 16192 22618 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 23017 16195 23075 16201
rect 23385 16235 23443 16241
rect 23385 16201 23397 16235
rect 23431 16232 23443 16235
rect 24026 16232 24032 16244
rect 23431 16204 24032 16232
rect 23431 16201 23443 16204
rect 23385 16195 23443 16201
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 26697 16235 26755 16241
rect 26697 16232 26709 16235
rect 25188 16204 26709 16232
rect 25188 16192 25194 16204
rect 26697 16201 26709 16204
rect 26743 16201 26755 16235
rect 26697 16195 26755 16201
rect 13078 16124 13084 16176
rect 13136 16164 13142 16176
rect 13173 16167 13231 16173
rect 13173 16164 13185 16167
rect 13136 16136 13185 16164
rect 13136 16124 13142 16136
rect 13173 16133 13185 16136
rect 13219 16164 13231 16167
rect 15381 16167 15439 16173
rect 13219 16136 13952 16164
rect 13219 16133 13231 16136
rect 13173 16127 13231 16133
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13495 16068 13737 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 13725 16065 13737 16068
rect 13771 16096 13783 16099
rect 13814 16096 13820 16108
rect 13771 16068 13820 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 13357 16031 13415 16037
rect 13357 15997 13369 16031
rect 13403 16028 13415 16031
rect 13630 16028 13636 16040
rect 13403 16000 13636 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 13740 15960 13768 16059
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 13924 16105 13952 16136
rect 15381 16133 15393 16167
rect 15427 16164 15439 16167
rect 15838 16164 15844 16176
rect 15427 16136 15844 16164
rect 15427 16133 15439 16136
rect 15381 16127 15439 16133
rect 15838 16124 15844 16136
rect 15896 16124 15902 16176
rect 20349 16167 20407 16173
rect 20349 16133 20361 16167
rect 20395 16133 20407 16167
rect 20349 16127 20407 16133
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 13924 16028 13952 16059
rect 14734 16056 14740 16108
rect 14792 16056 14798 16108
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 15252 16068 15301 16096
rect 15252 16056 15258 16068
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15289 16059 15347 16065
rect 15396 16068 15485 16096
rect 15396 16040 15424 16068
rect 15473 16065 15485 16068
rect 15519 16096 15531 16099
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15519 16068 15761 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 16022 16056 16028 16108
rect 16080 16056 16086 16108
rect 16209 16099 16267 16105
rect 16209 16065 16221 16099
rect 16255 16065 16267 16099
rect 16209 16059 16267 16065
rect 14826 16028 14832 16040
rect 13924 16000 14832 16028
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 16028 15071 16031
rect 15059 16000 15240 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 15102 15960 15108 15972
rect 13740 15932 15108 15960
rect 15102 15920 15108 15932
rect 15160 15920 15166 15972
rect 15212 15960 15240 16000
rect 15378 15988 15384 16040
rect 15436 15988 15442 16040
rect 15654 15960 15660 15972
rect 15212 15932 15660 15960
rect 15654 15920 15660 15932
rect 15712 15920 15718 15972
rect 16224 15904 16252 16059
rect 16666 16056 16672 16108
rect 16724 16056 16730 16108
rect 16758 16056 16764 16108
rect 16816 16096 16822 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16816 16068 16865 16096
rect 16816 16056 16822 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 17175 16068 17724 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 17144 16028 17172 16059
rect 16448 16000 17172 16028
rect 16448 15988 16454 16000
rect 17696 15960 17724 16068
rect 17954 16056 17960 16108
rect 18012 16056 18018 16108
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 18156 16028 18184 16059
rect 18230 16056 18236 16108
rect 18288 16056 18294 16108
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16096 18383 16099
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 18371 16068 18705 16096
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 18693 16065 18705 16068
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 18782 16056 18788 16108
rect 18840 16096 18846 16108
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 18840 16068 19257 16096
rect 18840 16056 18846 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 20254 16056 20260 16108
rect 20312 16056 20318 16108
rect 19610 16028 19616 16040
rect 18156 16000 19616 16028
rect 19610 15988 19616 16000
rect 19668 16028 19674 16040
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 19668 16000 19809 16028
rect 19668 15988 19674 16000
rect 19797 15997 19809 16000
rect 19843 16028 19855 16031
rect 20162 16028 20168 16040
rect 19843 16000 20168 16028
rect 19843 15997 19855 16000
rect 19797 15991 19855 15997
rect 20162 15988 20168 16000
rect 20220 16028 20226 16040
rect 20364 16028 20392 16127
rect 21082 16124 21088 16176
rect 21140 16164 21146 16176
rect 23477 16167 23535 16173
rect 21140 16136 21588 16164
rect 21140 16124 21146 16136
rect 20806 16056 20812 16108
rect 20864 16056 20870 16108
rect 21560 16105 21588 16136
rect 23477 16133 23489 16167
rect 23523 16164 23535 16167
rect 24118 16164 24124 16176
rect 23523 16136 24124 16164
rect 23523 16133 23535 16136
rect 23477 16127 23535 16133
rect 24118 16124 24124 16136
rect 24176 16124 24182 16176
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21453 16099 21511 16105
rect 21453 16096 21465 16099
rect 21039 16068 21465 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21453 16065 21465 16068
rect 21499 16065 21511 16099
rect 21453 16059 21511 16065
rect 21545 16099 21603 16105
rect 21545 16065 21557 16099
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 20220 16000 20392 16028
rect 20220 15988 20226 16000
rect 20530 15988 20536 16040
rect 20588 16028 20594 16040
rect 21008 16028 21036 16059
rect 24946 16056 24952 16108
rect 25004 16056 25010 16108
rect 26712 16096 26740 16195
rect 28074 16192 28080 16244
rect 28132 16192 28138 16244
rect 28258 16192 28264 16244
rect 28316 16192 28322 16244
rect 31386 16232 31392 16244
rect 29380 16204 31392 16232
rect 29089 16167 29147 16173
rect 29089 16133 29101 16167
rect 29135 16133 29147 16167
rect 29089 16127 29147 16133
rect 27525 16099 27583 16105
rect 27525 16096 27537 16099
rect 20588 16000 21036 16028
rect 23569 16031 23627 16037
rect 20588 15988 20594 16000
rect 23569 15997 23581 16031
rect 23615 15997 23627 16031
rect 23569 15991 23627 15997
rect 19334 15960 19340 15972
rect 17696 15932 19340 15960
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 20548 15932 21189 15960
rect 13173 15895 13231 15901
rect 13173 15892 13185 15895
rect 12406 15864 13185 15892
rect 5261 15855 5319 15861
rect 13173 15861 13185 15864
rect 13219 15892 13231 15895
rect 13538 15892 13544 15904
rect 13219 15864 13544 15892
rect 13219 15861 13231 15864
rect 13173 15855 13231 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 13909 15895 13967 15901
rect 13909 15892 13921 15895
rect 13872 15864 13921 15892
rect 13872 15852 13878 15864
rect 13909 15861 13921 15864
rect 13955 15861 13967 15895
rect 13909 15855 13967 15861
rect 14366 15852 14372 15904
rect 14424 15852 14430 15904
rect 15194 15852 15200 15904
rect 15252 15892 15258 15904
rect 16206 15892 16212 15904
rect 15252 15864 16212 15892
rect 15252 15852 15258 15864
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 20548 15901 20576 15932
rect 21177 15929 21189 15932
rect 21223 15929 21235 15963
rect 21177 15923 21235 15929
rect 23198 15920 23204 15972
rect 23256 15960 23262 15972
rect 23584 15960 23612 15991
rect 25222 15988 25228 16040
rect 25280 15988 25286 16040
rect 26344 16028 26372 16082
rect 26712 16068 27537 16096
rect 27525 16065 27537 16068
rect 27571 16065 27583 16099
rect 27525 16059 27583 16065
rect 28258 16099 28316 16105
rect 28258 16065 28270 16099
rect 28304 16096 28316 16099
rect 29104 16096 29132 16127
rect 29380 16105 29408 16204
rect 31386 16192 31392 16204
rect 31444 16192 31450 16244
rect 31895 16235 31953 16241
rect 31895 16201 31907 16235
rect 31941 16232 31953 16235
rect 32214 16232 32220 16244
rect 31941 16204 32220 16232
rect 31941 16201 31953 16204
rect 31895 16195 31953 16201
rect 32214 16192 32220 16204
rect 32272 16192 32278 16244
rect 31202 16124 31208 16176
rect 31260 16124 31266 16176
rect 31662 16164 31668 16176
rect 31594 16136 31668 16164
rect 28304 16068 29132 16096
rect 29365 16099 29423 16105
rect 28304 16065 28316 16068
rect 28258 16059 28316 16065
rect 29365 16065 29377 16099
rect 29411 16065 29423 16099
rect 29365 16059 29423 16065
rect 29454 16056 29460 16108
rect 29512 16096 29518 16108
rect 31220 16096 31248 16124
rect 31594 16096 31622 16136
rect 31662 16124 31668 16136
rect 31720 16124 31726 16176
rect 32493 16099 32551 16105
rect 32493 16096 32505 16099
rect 29512 16068 30604 16096
rect 31220 16068 31622 16096
rect 31726 16068 32505 16096
rect 29512 16056 29518 16068
rect 27982 16028 27988 16040
rect 26344 16000 27988 16028
rect 27982 15988 27988 16000
rect 28040 15988 28046 16040
rect 28721 16031 28779 16037
rect 28721 15997 28733 16031
rect 28767 16028 28779 16031
rect 28994 16028 29000 16040
rect 28767 16000 29000 16028
rect 28767 15997 28779 16000
rect 28721 15991 28779 15997
rect 28994 15988 29000 16000
rect 29052 15988 29058 16040
rect 29086 15988 29092 16040
rect 29144 15988 29150 16040
rect 29546 15988 29552 16040
rect 29604 16028 29610 16040
rect 30101 16031 30159 16037
rect 30101 16028 30113 16031
rect 29604 16000 30113 16028
rect 29604 15988 29610 16000
rect 30101 15997 30113 16000
rect 30147 15997 30159 16031
rect 30101 15991 30159 15997
rect 30466 15988 30472 16040
rect 30524 15988 30530 16040
rect 30576 16028 30604 16068
rect 31726 16028 31754 16068
rect 32493 16065 32505 16068
rect 32539 16096 32551 16099
rect 33137 16099 33195 16105
rect 33137 16096 33149 16099
rect 32539 16068 33149 16096
rect 32539 16065 32551 16068
rect 32493 16059 32551 16065
rect 33137 16065 33149 16068
rect 33183 16096 33195 16099
rect 35342 16096 35348 16108
rect 33183 16068 35348 16096
rect 33183 16065 33195 16068
rect 33137 16059 33195 16065
rect 35342 16056 35348 16068
rect 35400 16056 35406 16108
rect 30576 16000 31754 16028
rect 32858 15988 32864 16040
rect 32916 16028 32922 16040
rect 33965 16031 34023 16037
rect 33965 16028 33977 16031
rect 32916 16000 33977 16028
rect 32916 15988 32922 16000
rect 33965 15997 33977 16000
rect 34011 16028 34023 16031
rect 34606 16028 34612 16040
rect 34011 16000 34612 16028
rect 34011 15997 34023 16000
rect 33965 15991 34023 15997
rect 34606 15988 34612 16000
rect 34664 16028 34670 16040
rect 34790 16028 34796 16040
rect 34664 16000 34796 16028
rect 34664 15988 34670 16000
rect 34790 15988 34796 16000
rect 34848 15988 34854 16040
rect 23256 15932 23612 15960
rect 23256 15920 23262 15932
rect 27798 15920 27804 15972
rect 27856 15960 27862 15972
rect 28626 15960 28632 15972
rect 27856 15932 28632 15960
rect 27856 15920 27862 15932
rect 28626 15920 28632 15932
rect 28684 15920 28690 15972
rect 32769 15963 32827 15969
rect 32769 15929 32781 15963
rect 32815 15960 32827 15963
rect 33134 15960 33140 15972
rect 32815 15932 33140 15960
rect 32815 15929 32827 15932
rect 32769 15923 32827 15929
rect 33134 15920 33140 15932
rect 33192 15920 33198 15972
rect 20533 15895 20591 15901
rect 20533 15861 20545 15895
rect 20579 15861 20591 15895
rect 20533 15855 20591 15861
rect 20714 15852 20720 15904
rect 20772 15852 20778 15904
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 26878 15852 26884 15904
rect 26936 15892 26942 15904
rect 26973 15895 27031 15901
rect 26973 15892 26985 15895
rect 26936 15864 26985 15892
rect 26936 15852 26942 15864
rect 26973 15861 26985 15864
rect 27019 15861 27031 15895
rect 26973 15855 27031 15861
rect 29273 15895 29331 15901
rect 29273 15861 29285 15895
rect 29319 15892 29331 15895
rect 30650 15892 30656 15904
rect 29319 15864 30656 15892
rect 29319 15861 29331 15864
rect 29273 15855 29331 15861
rect 30650 15852 30656 15864
rect 30708 15852 30714 15904
rect 32861 15895 32919 15901
rect 32861 15861 32873 15895
rect 32907 15892 32919 15895
rect 32950 15892 32956 15904
rect 32907 15864 32956 15892
rect 32907 15861 32919 15864
rect 32861 15855 32919 15861
rect 32950 15852 32956 15864
rect 33008 15852 33014 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 2556 15660 2881 15688
rect 2556 15648 2562 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 2869 15651 2927 15657
rect 4157 15691 4215 15697
rect 4157 15657 4169 15691
rect 4203 15688 4215 15691
rect 4614 15688 4620 15700
rect 4203 15660 4620 15688
rect 4203 15657 4215 15660
rect 4157 15651 4215 15657
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 5169 15691 5227 15697
rect 5169 15657 5181 15691
rect 5215 15688 5227 15691
rect 5258 15688 5264 15700
rect 5215 15660 5264 15688
rect 5215 15657 5227 15660
rect 5169 15651 5227 15657
rect 5258 15648 5264 15660
rect 5316 15688 5322 15700
rect 7006 15688 7012 15700
rect 5316 15660 7012 15688
rect 5316 15648 5322 15660
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 10870 15648 10876 15700
rect 10928 15688 10934 15700
rect 10928 15660 12572 15688
rect 10928 15648 10934 15660
rect 4246 15580 4252 15632
rect 4304 15620 4310 15632
rect 5074 15620 5080 15632
rect 4304 15592 5080 15620
rect 4304 15580 4310 15592
rect 5074 15580 5080 15592
rect 5132 15580 5138 15632
rect 12544 15629 12572 15660
rect 13262 15648 13268 15700
rect 13320 15648 13326 15700
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 15933 15691 15991 15697
rect 15933 15688 15945 15691
rect 15436 15660 15945 15688
rect 15436 15648 15442 15660
rect 15933 15657 15945 15660
rect 15979 15657 15991 15691
rect 15933 15651 15991 15657
rect 16022 15648 16028 15700
rect 16080 15688 16086 15700
rect 16485 15691 16543 15697
rect 16485 15688 16497 15691
rect 16080 15660 16497 15688
rect 16080 15648 16086 15660
rect 16485 15657 16497 15660
rect 16531 15657 16543 15691
rect 16485 15651 16543 15657
rect 16942 15648 16948 15700
rect 17000 15688 17006 15700
rect 17589 15691 17647 15697
rect 17589 15688 17601 15691
rect 17000 15660 17601 15688
rect 17000 15648 17006 15660
rect 17589 15657 17601 15660
rect 17635 15688 17647 15691
rect 18414 15688 18420 15700
rect 17635 15660 18420 15688
rect 17635 15657 17647 15660
rect 17589 15651 17647 15657
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 23106 15648 23112 15700
rect 23164 15688 23170 15700
rect 29549 15691 29607 15697
rect 29549 15688 29561 15691
rect 23164 15660 29561 15688
rect 23164 15648 23170 15660
rect 29549 15657 29561 15660
rect 29595 15657 29607 15691
rect 29549 15651 29607 15657
rect 12529 15623 12587 15629
rect 12529 15589 12541 15623
rect 12575 15620 12587 15623
rect 13630 15620 13636 15632
rect 12575 15592 13636 15620
rect 12575 15589 12587 15592
rect 12529 15583 12587 15589
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 4062 15552 4068 15564
rect 3283 15524 4068 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 4062 15512 4068 15524
rect 4120 15552 4126 15564
rect 4433 15555 4491 15561
rect 4433 15552 4445 15555
rect 4120 15524 4445 15552
rect 4120 15512 4126 15524
rect 4433 15521 4445 15524
rect 4479 15521 4491 15555
rect 5350 15552 5356 15564
rect 4433 15515 4491 15521
rect 4724 15524 5356 15552
rect 2498 15444 2504 15496
rect 2556 15444 2562 15496
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 2958 15484 2964 15496
rect 2731 15456 2964 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3050 15444 3056 15496
rect 3108 15444 3114 15496
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15484 4399 15487
rect 4724 15484 4752 15524
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 4387 15456 4752 15484
rect 4801 15487 4859 15493
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 4801 15453 4813 15487
rect 4847 15484 4859 15487
rect 5258 15484 5264 15496
rect 4847 15456 5264 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 12636 15493 12664 15592
rect 13630 15580 13636 15592
rect 13688 15580 13694 15632
rect 16390 15580 16396 15632
rect 16448 15580 16454 15632
rect 16666 15580 16672 15632
rect 16724 15620 16730 15632
rect 16850 15620 16856 15632
rect 16724 15592 16856 15620
rect 16724 15580 16730 15592
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 25222 15580 25228 15632
rect 25280 15580 25286 15632
rect 25608 15592 25820 15620
rect 12710 15512 12716 15564
rect 12768 15552 12774 15564
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 12768 15524 14105 15552
rect 12768 15512 12774 15524
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 14093 15515 14151 15521
rect 14366 15512 14372 15564
rect 14424 15512 14430 15564
rect 14826 15512 14832 15564
rect 14884 15552 14890 15564
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 14884 15524 15853 15552
rect 14884 15512 14890 15524
rect 15841 15521 15853 15524
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 16022 15512 16028 15564
rect 16080 15512 16086 15564
rect 18046 15552 18052 15564
rect 17788 15524 18052 15552
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 9272 15456 10057 15484
rect 9272 15444 9278 15456
rect 10045 15453 10057 15456
rect 10091 15484 10103 15487
rect 10781 15487 10839 15493
rect 10781 15484 10793 15487
rect 10091 15456 10793 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10781 15453 10793 15456
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 12805 15487 12863 15493
rect 12805 15453 12817 15487
rect 12851 15484 12863 15487
rect 12894 15484 12900 15496
rect 12851 15456 12900 15484
rect 12851 15453 12863 15456
rect 12805 15447 12863 15453
rect 3142 15376 3148 15428
rect 3200 15416 3206 15428
rect 4709 15419 4767 15425
rect 4709 15416 4721 15419
rect 3200 15388 4721 15416
rect 3200 15376 3206 15388
rect 4709 15385 4721 15388
rect 4755 15385 4767 15419
rect 4709 15379 4767 15385
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 2593 15351 2651 15357
rect 2593 15348 2605 15351
rect 2464 15320 2605 15348
rect 2464 15308 2470 15320
rect 2593 15317 2605 15320
rect 2639 15317 2651 15351
rect 2593 15311 2651 15317
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15348 4675 15351
rect 4890 15348 4896 15360
rect 4663 15320 4896 15348
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 10796 15348 10824 15447
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13078 15444 13084 15496
rect 13136 15444 13142 15496
rect 13538 15444 13544 15496
rect 13596 15444 13602 15496
rect 13722 15444 13728 15496
rect 13780 15444 13786 15496
rect 13814 15444 13820 15496
rect 13872 15444 13878 15496
rect 15470 15444 15476 15496
rect 15528 15444 15534 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15804 15456 15945 15484
rect 15804 15444 15810 15456
rect 15933 15453 15945 15456
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 16206 15444 16212 15496
rect 16264 15444 16270 15496
rect 17788 15493 17816 15524
rect 18046 15512 18052 15524
rect 18104 15552 18110 15564
rect 18104 15524 18460 15552
rect 18104 15512 18110 15524
rect 18432 15493 18460 15524
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 22005 15555 22063 15561
rect 22005 15552 22017 15555
rect 20772 15524 22017 15552
rect 20772 15512 20778 15524
rect 22005 15521 22017 15524
rect 22051 15521 22063 15555
rect 22005 15515 22063 15521
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 25608 15552 25636 15592
rect 24176 15524 25636 15552
rect 24176 15512 24182 15524
rect 25682 15512 25688 15564
rect 25740 15512 25746 15564
rect 25792 15561 25820 15592
rect 27798 15580 27804 15632
rect 27856 15580 27862 15632
rect 25777 15555 25835 15561
rect 25777 15521 25789 15555
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 17773 15487 17831 15493
rect 17773 15453 17785 15487
rect 17819 15453 17831 15487
rect 17773 15447 17831 15453
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15484 18015 15487
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 18003 15456 18245 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 18233 15453 18245 15456
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15484 18475 15487
rect 18874 15484 18880 15496
rect 18463 15456 18880 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 11054 15376 11060 15428
rect 11112 15376 11118 15428
rect 11790 15376 11796 15428
rect 11848 15376 11854 15428
rect 12710 15416 12716 15428
rect 12452 15388 12716 15416
rect 12452 15348 12480 15388
rect 12710 15376 12716 15388
rect 12768 15376 12774 15428
rect 12986 15376 12992 15428
rect 13044 15416 13050 15428
rect 13357 15419 13415 15425
rect 13357 15416 13369 15419
rect 13044 15388 13369 15416
rect 13044 15376 13050 15388
rect 13357 15385 13369 15388
rect 13403 15385 13415 15419
rect 13357 15379 13415 15385
rect 16758 15376 16764 15428
rect 16816 15416 16822 15428
rect 16945 15419 17003 15425
rect 16945 15416 16957 15419
rect 16816 15388 16957 15416
rect 16816 15376 16822 15388
rect 16945 15385 16957 15388
rect 16991 15385 17003 15419
rect 16945 15379 17003 15385
rect 17126 15376 17132 15428
rect 17184 15416 17190 15428
rect 18049 15419 18107 15425
rect 18049 15416 18061 15419
rect 17184 15388 18061 15416
rect 17184 15376 17190 15388
rect 18049 15385 18061 15388
rect 18095 15385 18107 15419
rect 18248 15416 18276 15447
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 18969 15487 19027 15493
rect 18969 15453 18981 15487
rect 19015 15484 19027 15487
rect 19058 15484 19064 15496
rect 19015 15456 19064 15484
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 19058 15444 19064 15456
rect 19116 15484 19122 15496
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19116 15456 19993 15484
rect 19116 15444 19122 15456
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15484 22339 15487
rect 22649 15487 22707 15493
rect 22649 15484 22661 15487
rect 22327 15456 22661 15484
rect 22327 15453 22339 15456
rect 22281 15447 22339 15453
rect 22649 15453 22661 15456
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 18690 15416 18696 15428
rect 18248 15388 18696 15416
rect 18049 15379 18107 15385
rect 18690 15376 18696 15388
rect 18748 15416 18754 15428
rect 18748 15388 18920 15416
rect 18748 15376 18754 15388
rect 10796 15320 12480 15348
rect 15654 15308 15660 15360
rect 15712 15348 15718 15360
rect 17144 15348 17172 15376
rect 18892 15360 18920 15388
rect 19242 15376 19248 15428
rect 19300 15376 19306 15428
rect 22002 15416 22008 15428
rect 21574 15388 22008 15416
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 22094 15376 22100 15428
rect 22152 15416 22158 15428
rect 22296 15416 22324 15447
rect 24946 15444 24952 15496
rect 25004 15444 25010 15496
rect 25593 15487 25651 15493
rect 25593 15453 25605 15487
rect 25639 15484 25651 15487
rect 26878 15484 26884 15496
rect 25639 15456 26884 15484
rect 25639 15453 25651 15456
rect 25593 15447 25651 15453
rect 26878 15444 26884 15456
rect 26936 15444 26942 15496
rect 26970 15444 26976 15496
rect 27028 15444 27034 15496
rect 29564 15484 29592 15651
rect 32585 15555 32643 15561
rect 32585 15521 32597 15555
rect 32631 15552 32643 15555
rect 32858 15552 32864 15564
rect 32631 15524 32864 15552
rect 32631 15521 32643 15524
rect 32585 15515 32643 15521
rect 32858 15512 32864 15524
rect 32916 15512 32922 15564
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29564 15456 29745 15484
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 37274 15444 37280 15496
rect 37332 15444 37338 15496
rect 22152 15388 22324 15416
rect 22152 15376 22158 15388
rect 28166 15376 28172 15428
rect 28224 15376 28230 15428
rect 32861 15419 32919 15425
rect 32861 15385 32873 15419
rect 32907 15416 32919 15419
rect 32950 15416 32956 15428
rect 32907 15388 32956 15416
rect 32907 15385 32919 15388
rect 32861 15379 32919 15385
rect 32950 15376 32956 15388
rect 33008 15376 33014 15428
rect 34422 15416 34428 15428
rect 34086 15388 34428 15416
rect 34422 15376 34428 15388
rect 34480 15376 34486 15428
rect 34514 15376 34520 15428
rect 34572 15416 34578 15428
rect 35253 15419 35311 15425
rect 35253 15416 35265 15419
rect 34572 15388 35265 15416
rect 34572 15376 34578 15388
rect 35253 15385 35265 15388
rect 35299 15385 35311 15419
rect 35253 15379 35311 15385
rect 35434 15376 35440 15428
rect 35492 15376 35498 15428
rect 15712 15320 17172 15348
rect 15712 15308 15718 15320
rect 18874 15308 18880 15360
rect 18932 15308 18938 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 20530 15348 20536 15360
rect 19484 15320 20536 15348
rect 19484 15308 19490 15320
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 23934 15348 23940 15360
rect 23716 15320 23940 15348
rect 23716 15308 23722 15320
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 24118 15308 24124 15360
rect 24176 15308 24182 15360
rect 24394 15308 24400 15360
rect 24452 15308 24458 15360
rect 27614 15308 27620 15360
rect 27672 15308 27678 15360
rect 27706 15308 27712 15360
rect 27764 15308 27770 15360
rect 30098 15308 30104 15360
rect 30156 15348 30162 15360
rect 31021 15351 31079 15357
rect 31021 15348 31033 15351
rect 30156 15320 31033 15348
rect 30156 15308 30162 15320
rect 31021 15317 31033 15320
rect 31067 15348 31079 15351
rect 31573 15351 31631 15357
rect 31573 15348 31585 15351
rect 31067 15320 31585 15348
rect 31067 15317 31079 15320
rect 31021 15311 31079 15317
rect 31573 15317 31585 15320
rect 31619 15317 31631 15351
rect 31573 15311 31631 15317
rect 34333 15351 34391 15357
rect 34333 15317 34345 15351
rect 34379 15348 34391 15351
rect 34698 15348 34704 15360
rect 34379 15320 34704 15348
rect 34379 15317 34391 15320
rect 34333 15311 34391 15317
rect 34698 15308 34704 15320
rect 34756 15308 34762 15360
rect 36630 15308 36636 15360
rect 36688 15308 36694 15360
rect 38470 15308 38476 15360
rect 38528 15308 38534 15360
rect 1104 15258 38824 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 38824 15258
rect 1104 15184 38824 15206
rect 3602 15104 3608 15156
rect 3660 15144 3666 15156
rect 5718 15144 5724 15156
rect 3660 15116 5724 15144
rect 3660 15104 3666 15116
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 8294 15144 8300 15156
rect 6656 15116 8300 15144
rect 4614 15036 4620 15088
rect 4672 15076 4678 15088
rect 4801 15079 4859 15085
rect 4801 15076 4813 15079
rect 4672 15048 4813 15076
rect 4672 15036 4678 15048
rect 4801 15045 4813 15048
rect 4847 15045 4859 15079
rect 4801 15039 4859 15045
rect 5442 15036 5448 15088
rect 5500 15076 5506 15088
rect 5500 15048 6132 15076
rect 5500 15036 5506 15048
rect 1394 14968 1400 15020
rect 1452 14968 1458 15020
rect 2774 14968 2780 15020
rect 2832 14968 2838 15020
rect 2958 14968 2964 15020
rect 3016 15008 3022 15020
rect 3016 14980 5028 15008
rect 3016 14968 3022 14980
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 2222 14940 2228 14952
rect 1719 14912 2228 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14940 3203 14943
rect 3881 14943 3939 14949
rect 3881 14940 3893 14943
rect 3191 14912 3893 14940
rect 3191 14909 3203 14912
rect 3145 14903 3203 14909
rect 3881 14909 3893 14912
rect 3927 14940 3939 14943
rect 4062 14940 4068 14952
rect 3927 14912 4068 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4522 14900 4528 14952
rect 4580 14940 4586 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4580 14912 4905 14940
rect 4580 14900 4586 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 3234 14764 3240 14816
rect 3292 14764 3298 14816
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 4246 14804 4252 14816
rect 3752 14776 4252 14804
rect 3752 14764 3758 14776
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4614 14764 4620 14816
rect 4672 14804 4678 14816
rect 4801 14807 4859 14813
rect 4801 14804 4813 14807
rect 4672 14776 4813 14804
rect 4672 14764 4678 14776
rect 4801 14773 4813 14776
rect 4847 14773 4859 14807
rect 5000 14804 5028 14980
rect 5074 14968 5080 15020
rect 5132 14968 5138 15020
rect 5626 15008 5632 15020
rect 5276 14980 5632 15008
rect 5276 14881 5304 14980
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 6104 15017 6132 15048
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 14977 5963 15011
rect 5905 14971 5963 14977
rect 6089 15011 6147 15017
rect 6089 14977 6101 15011
rect 6135 15008 6147 15011
rect 6546 15008 6552 15020
rect 6135 14980 6552 15008
rect 6135 14977 6147 14980
rect 6089 14971 6147 14977
rect 5350 14900 5356 14952
rect 5408 14940 5414 14952
rect 5920 14940 5948 14971
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 6656 15017 6684 15116
rect 8294 15104 8300 15116
rect 8352 15144 8358 15156
rect 9214 15144 9220 15156
rect 8352 15116 9220 15144
rect 8352 15104 8358 15116
rect 7466 15036 7472 15088
rect 7524 15036 7530 15088
rect 8772 15017 8800 15116
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 10870 15144 10876 15156
rect 9916 15116 10876 15144
rect 9916 15104 9922 15116
rect 10870 15104 10876 15116
rect 10928 15144 10934 15156
rect 10965 15147 11023 15153
rect 10965 15144 10977 15147
rect 10928 15116 10977 15144
rect 10928 15104 10934 15116
rect 10965 15113 10977 15116
rect 11011 15113 11023 15147
rect 10965 15107 11023 15113
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11333 15147 11391 15153
rect 11333 15144 11345 15147
rect 11112 15116 11345 15144
rect 11112 15104 11118 15116
rect 11333 15113 11345 15116
rect 11379 15113 11391 15147
rect 11333 15107 11391 15113
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 12250 15144 12256 15156
rect 11848 15116 12256 15144
rect 11848 15104 11854 15116
rect 12250 15104 12256 15116
rect 12308 15144 12314 15156
rect 13630 15144 13636 15156
rect 12308 15116 13636 15144
rect 12308 15104 12314 15116
rect 13630 15104 13636 15116
rect 13688 15104 13694 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 14274 15144 14280 15156
rect 13872 15116 14280 15144
rect 13872 15104 13878 15116
rect 14274 15104 14280 15116
rect 14332 15144 14338 15156
rect 14461 15147 14519 15153
rect 14461 15144 14473 15147
rect 14332 15116 14473 15144
rect 14332 15104 14338 15116
rect 14461 15113 14473 15116
rect 14507 15113 14519 15147
rect 14461 15107 14519 15113
rect 14553 15147 14611 15153
rect 14553 15113 14565 15147
rect 14599 15144 14611 15147
rect 14734 15144 14740 15156
rect 14599 15116 14740 15144
rect 14599 15113 14611 15116
rect 14553 15107 14611 15113
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 18509 15147 18567 15153
rect 18509 15144 18521 15147
rect 17788 15116 18521 15144
rect 10042 15036 10048 15088
rect 10100 15036 10106 15088
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11480 15048 11529 15076
rect 11480 15036 11486 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 13078 15076 13084 15088
rect 11517 15039 11575 15045
rect 11624 15048 13084 15076
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 6917 14943 6975 14949
rect 6917 14940 6929 14943
rect 5408 14912 5948 14940
rect 6012 14912 6929 14940
rect 5408 14900 5414 14912
rect 5261 14875 5319 14881
rect 5261 14841 5273 14875
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 5721 14875 5779 14881
rect 5721 14841 5733 14875
rect 5767 14872 5779 14875
rect 6012 14872 6040 14912
rect 6917 14909 6929 14912
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 8662 14900 8668 14952
rect 8720 14900 8726 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 9582 14940 9588 14952
rect 9079 14912 9588 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 10686 14900 10692 14952
rect 10744 14900 10750 14952
rect 10873 14943 10931 14949
rect 10873 14909 10885 14943
rect 10919 14940 10931 14943
rect 11624 14940 11652 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 14826 15076 14832 15088
rect 14214 15062 14832 15076
rect 14200 15048 14832 15062
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12710 15008 12716 15020
rect 12492 14980 12716 15008
rect 12492 14968 12498 14980
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 10919 14912 11652 14940
rect 10919 14909 10931 14912
rect 10873 14903 10931 14909
rect 12342 14900 12348 14952
rect 12400 14940 12406 14952
rect 12529 14943 12587 14949
rect 12529 14940 12541 14943
rect 12400 14912 12541 14940
rect 12400 14900 12406 14912
rect 12529 14909 12541 14912
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 12986 14900 12992 14952
rect 13044 14900 13050 14952
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 14200 14940 14228 15048
rect 14826 15036 14832 15048
rect 14884 15076 14890 15088
rect 15470 15076 15476 15088
rect 14884 15048 15476 15076
rect 14884 15036 14890 15048
rect 15470 15036 15476 15048
rect 15528 15036 15534 15088
rect 17788 15017 17816 15116
rect 18509 15113 18521 15116
rect 18555 15113 18567 15147
rect 18509 15107 18567 15113
rect 18782 15104 18788 15156
rect 18840 15144 18846 15156
rect 19518 15144 19524 15156
rect 18840 15116 19524 15144
rect 18840 15104 18846 15116
rect 19518 15104 19524 15116
rect 19576 15104 19582 15156
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 20254 15144 20260 15156
rect 19751 15116 20260 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 23937 15147 23995 15153
rect 22060 15116 23796 15144
rect 22060 15104 22066 15116
rect 18877 15079 18935 15085
rect 18877 15045 18889 15079
rect 18923 15076 18935 15079
rect 19889 15079 19947 15085
rect 19889 15076 19901 15079
rect 18923 15048 19901 15076
rect 18923 15045 18935 15048
rect 18877 15039 18935 15045
rect 19889 15045 19901 15048
rect 19935 15045 19947 15079
rect 19889 15039 19947 15045
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 20714 15076 20720 15088
rect 20211 15048 20720 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 20714 15036 20720 15048
rect 20772 15076 20778 15088
rect 21266 15076 21272 15088
rect 20772 15048 21272 15076
rect 20772 15036 20778 15048
rect 21266 15036 21272 15048
rect 21324 15036 21330 15088
rect 23768 15076 23796 15116
rect 23937 15113 23949 15147
rect 23983 15144 23995 15147
rect 24946 15144 24952 15156
rect 23983 15116 24952 15144
rect 23983 15113 23995 15116
rect 23937 15107 23995 15113
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 28166 15104 28172 15156
rect 28224 15144 28230 15156
rect 28721 15147 28779 15153
rect 28721 15144 28733 15147
rect 28224 15116 28733 15144
rect 28224 15104 28230 15116
rect 28721 15113 28733 15116
rect 28767 15113 28779 15147
rect 28721 15107 28779 15113
rect 29454 15104 29460 15156
rect 29512 15144 29518 15156
rect 30098 15144 30104 15156
rect 29512 15116 30104 15144
rect 29512 15104 29518 15116
rect 30098 15104 30104 15116
rect 30156 15104 30162 15156
rect 35986 15144 35992 15156
rect 35360 15116 35992 15144
rect 23842 15076 23848 15088
rect 23690 15048 23848 15076
rect 23842 15036 23848 15048
rect 23900 15076 23906 15088
rect 23900 15048 24794 15076
rect 23900 15036 23906 15048
rect 27982 15036 27988 15088
rect 28040 15036 28046 15088
rect 33134 15036 33140 15088
rect 33192 15036 33198 15088
rect 34422 15076 34428 15088
rect 34362 15048 34428 15076
rect 34422 15036 34428 15048
rect 34480 15076 34486 15088
rect 35360 15076 35388 15116
rect 35986 15104 35992 15116
rect 36044 15144 36050 15156
rect 36044 15116 36400 15144
rect 36044 15104 36050 15116
rect 36372 15076 36400 15116
rect 37458 15076 37464 15088
rect 34480 15048 35388 15076
rect 36294 15048 37464 15076
rect 34480 15036 34486 15048
rect 37458 15036 37464 15048
rect 37516 15036 37522 15088
rect 17681 15011 17739 15017
rect 17681 15008 17693 15011
rect 17512 14980 17693 15008
rect 13688 14912 14228 14940
rect 13688 14900 13694 14912
rect 15102 14900 15108 14952
rect 15160 14900 15166 14952
rect 5767 14844 6040 14872
rect 17512 14872 17540 14980
rect 17681 14977 17693 14980
rect 17727 14977 17739 15011
rect 17681 14971 17739 14977
rect 17773 15011 17831 15017
rect 17773 14977 17785 15011
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 17954 14968 17960 15020
rect 18012 14968 18018 15020
rect 18690 14968 18696 15020
rect 18748 14968 18754 15020
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 17589 14943 17647 14949
rect 17589 14909 17601 14943
rect 17635 14940 17647 14943
rect 17972 14940 18000 14968
rect 17635 14912 18000 14940
rect 18800 14940 18828 14971
rect 18966 14968 18972 15020
rect 19024 15008 19030 15020
rect 19061 15011 19119 15017
rect 19061 15008 19073 15011
rect 19024 14980 19073 15008
rect 19024 14968 19030 14980
rect 19061 14977 19073 14980
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 19150 14968 19156 15020
rect 19208 14968 19214 15020
rect 19426 14968 19432 15020
rect 19484 14968 19490 15020
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 14977 19579 15011
rect 19521 14971 19579 14977
rect 18874 14940 18880 14952
rect 18800 14912 18880 14940
rect 17635 14909 17647 14912
rect 17589 14903 17647 14909
rect 18874 14900 18880 14912
rect 18932 14900 18938 14952
rect 19168 14940 19196 14968
rect 19536 14940 19564 14971
rect 19702 14968 19708 15020
rect 19760 15008 19766 15020
rect 19797 15011 19855 15017
rect 19797 15008 19809 15011
rect 19760 14980 19809 15008
rect 19760 14968 19766 14980
rect 19797 14977 19809 14980
rect 19843 14977 19855 15011
rect 19797 14971 19855 14977
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20088 14940 20116 14971
rect 20346 14968 20352 15020
rect 20404 14968 20410 15020
rect 24029 15011 24087 15017
rect 24029 15008 24041 15011
rect 23676 14980 24041 15008
rect 20806 14940 20812 14952
rect 18984 14912 20812 14940
rect 18984 14872 19012 14912
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22189 14943 22247 14949
rect 22189 14940 22201 14943
rect 22152 14912 22201 14940
rect 22152 14900 22158 14912
rect 22189 14909 22201 14912
rect 22235 14909 22247 14943
rect 22189 14903 22247 14909
rect 22462 14900 22468 14952
rect 22520 14900 22526 14952
rect 17512 14844 19012 14872
rect 5767 14841 5779 14844
rect 5721 14835 5779 14841
rect 5736 14804 5764 14835
rect 19242 14832 19248 14884
rect 19300 14832 19306 14884
rect 19978 14832 19984 14884
rect 20036 14872 20042 14884
rect 20036 14844 22094 14872
rect 20036 14832 20042 14844
rect 5000 14776 5764 14804
rect 4801 14767 4859 14773
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 5997 14807 6055 14813
rect 5997 14804 6009 14807
rect 5868 14776 6009 14804
rect 5868 14764 5874 14776
rect 5997 14773 6009 14776
rect 6043 14773 6055 14807
rect 5997 14767 6055 14773
rect 10502 14764 10508 14816
rect 10560 14764 10566 14816
rect 18417 14807 18475 14813
rect 18417 14773 18429 14807
rect 18463 14804 18475 14807
rect 18782 14804 18788 14816
rect 18463 14776 18788 14804
rect 18463 14773 18475 14776
rect 18417 14767 18475 14773
rect 18782 14764 18788 14776
rect 18840 14764 18846 14816
rect 18874 14764 18880 14816
rect 18932 14804 18938 14816
rect 19996 14804 20024 14832
rect 18932 14776 20024 14804
rect 18932 14764 18938 14776
rect 20530 14764 20536 14816
rect 20588 14764 20594 14816
rect 22066 14804 22094 14844
rect 23198 14804 23204 14816
rect 22066 14776 23204 14804
rect 23198 14764 23204 14776
rect 23256 14804 23262 14816
rect 23676 14804 23704 14980
rect 24029 14977 24041 14980
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 24210 14968 24216 15020
rect 24268 14968 24274 15020
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 15008 26295 15011
rect 26786 15008 26792 15020
rect 26283 14980 26792 15008
rect 26283 14977 26295 14980
rect 26237 14971 26295 14977
rect 26786 14968 26792 14980
rect 26844 15008 26850 15020
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26844 14980 26985 15008
rect 26844 14968 26850 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 29822 14968 29828 15020
rect 29880 15008 29886 15020
rect 30377 15011 30435 15017
rect 30377 15008 30389 15011
rect 29880 14980 30389 15008
rect 29880 14968 29886 14980
rect 30377 14977 30389 14980
rect 30423 14977 30435 15011
rect 30377 14971 30435 14977
rect 30561 15011 30619 15017
rect 30561 14977 30573 15011
rect 30607 15008 30619 15011
rect 30742 15008 30748 15020
rect 30607 14980 30748 15008
rect 30607 14977 30619 14980
rect 30561 14971 30619 14977
rect 30742 14968 30748 14980
rect 30800 14968 30806 15020
rect 32858 14968 32864 15020
rect 32916 14968 32922 15020
rect 36630 14968 36636 15020
rect 36688 14968 36694 15020
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 24176 14912 24317 14940
rect 24176 14900 24182 14912
rect 24305 14909 24317 14912
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 25498 14900 25504 14952
rect 25556 14940 25562 14952
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25556 14912 25973 14940
rect 25556 14900 25562 14912
rect 25961 14909 25973 14912
rect 26007 14909 26019 14943
rect 25961 14903 26019 14909
rect 27249 14943 27307 14949
rect 27249 14909 27261 14943
rect 27295 14940 27307 14943
rect 27706 14940 27712 14952
rect 27295 14912 27712 14940
rect 27295 14909 27307 14912
rect 27249 14903 27307 14909
rect 27706 14900 27712 14912
rect 27764 14900 27770 14952
rect 34790 14900 34796 14952
rect 34848 14900 34854 14952
rect 35069 14943 35127 14949
rect 35069 14909 35081 14943
rect 35115 14940 35127 14943
rect 35434 14940 35440 14952
rect 35115 14912 35440 14940
rect 35115 14909 35127 14912
rect 35069 14903 35127 14909
rect 35434 14900 35440 14912
rect 35492 14900 35498 14952
rect 36078 14832 36084 14884
rect 36136 14872 36142 14884
rect 36725 14875 36783 14881
rect 36725 14872 36737 14875
rect 36136 14844 36737 14872
rect 36136 14832 36142 14844
rect 36725 14841 36737 14844
rect 36771 14841 36783 14875
rect 36725 14835 36783 14841
rect 23256 14776 23704 14804
rect 23256 14764 23262 14776
rect 24026 14764 24032 14816
rect 24084 14804 24090 14816
rect 24121 14807 24179 14813
rect 24121 14804 24133 14807
rect 24084 14776 24133 14804
rect 24084 14764 24090 14776
rect 24121 14773 24133 14776
rect 24167 14773 24179 14807
rect 24121 14767 24179 14773
rect 24489 14807 24547 14813
rect 24489 14773 24501 14807
rect 24535 14804 24547 14807
rect 24670 14804 24676 14816
rect 24535 14776 24676 14804
rect 24535 14773 24547 14776
rect 24489 14767 24547 14773
rect 24670 14764 24676 14776
rect 24728 14764 24734 14816
rect 30745 14807 30803 14813
rect 30745 14773 30757 14807
rect 30791 14804 30803 14807
rect 31018 14804 31024 14816
rect 30791 14776 31024 14804
rect 30791 14773 30803 14776
rect 30745 14767 30803 14773
rect 31018 14764 31024 14776
rect 31076 14764 31082 14816
rect 34606 14764 34612 14816
rect 34664 14764 34670 14816
rect 36538 14764 36544 14816
rect 36596 14804 36602 14816
rect 37274 14804 37280 14816
rect 36596 14776 37280 14804
rect 36596 14764 36602 14776
rect 37274 14764 37280 14776
rect 37332 14764 37338 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 2222 14560 2228 14612
rect 2280 14560 2286 14612
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 4571 14572 4752 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 4724 14544 4752 14572
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 4856 14572 5089 14600
rect 4856 14560 4862 14572
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 5169 14603 5227 14609
rect 5169 14569 5181 14603
rect 5215 14600 5227 14603
rect 5258 14600 5264 14612
rect 5215 14572 5264 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 9582 14560 9588 14612
rect 9640 14560 9646 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 11422 14600 11428 14612
rect 11204 14572 11428 14600
rect 11204 14560 11210 14572
rect 11422 14560 11428 14572
rect 11480 14600 11486 14612
rect 12342 14600 12348 14612
rect 11480 14572 12348 14600
rect 11480 14560 11486 14572
rect 12342 14560 12348 14572
rect 12400 14600 12406 14612
rect 13906 14600 13912 14612
rect 12400 14572 13912 14600
rect 12400 14560 12406 14572
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 17313 14603 17371 14609
rect 17313 14569 17325 14603
rect 17359 14600 17371 14603
rect 18046 14600 18052 14612
rect 17359 14572 18052 14600
rect 17359 14569 17371 14572
rect 17313 14563 17371 14569
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19978 14600 19984 14612
rect 19392 14572 19984 14600
rect 19392 14560 19398 14572
rect 19978 14560 19984 14572
rect 20036 14600 20042 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 20036 14572 20085 14600
rect 20036 14560 20042 14572
rect 20073 14569 20085 14572
rect 20119 14600 20131 14603
rect 20346 14600 20352 14612
rect 20119 14572 20352 14600
rect 20119 14569 20131 14572
rect 20073 14563 20131 14569
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 22462 14560 22468 14612
rect 22520 14600 22526 14612
rect 23661 14603 23719 14609
rect 23661 14600 23673 14603
rect 22520 14572 23673 14600
rect 22520 14560 22526 14572
rect 23661 14569 23673 14572
rect 23707 14569 23719 14603
rect 23661 14563 23719 14569
rect 24121 14603 24179 14609
rect 24121 14569 24133 14603
rect 24167 14600 24179 14603
rect 24394 14600 24400 14612
rect 24167 14572 24400 14600
rect 24167 14569 24179 14572
rect 24121 14563 24179 14569
rect 24394 14560 24400 14572
rect 24452 14560 24458 14612
rect 25038 14600 25044 14612
rect 24596 14572 25044 14600
rect 2133 14535 2191 14541
rect 2133 14501 2145 14535
rect 2179 14532 2191 14535
rect 4249 14535 4307 14541
rect 2179 14504 3832 14532
rect 2179 14501 2191 14504
rect 2133 14495 2191 14501
rect 2685 14467 2743 14473
rect 2685 14433 2697 14467
rect 2731 14464 2743 14467
rect 3234 14464 3240 14476
rect 2731 14436 3240 14464
rect 2731 14433 2743 14436
rect 2685 14427 2743 14433
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 3602 14424 3608 14476
rect 3660 14424 3666 14476
rect 1854 14356 1860 14408
rect 1912 14356 1918 14408
rect 2406 14356 2412 14408
rect 2464 14356 2470 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 3050 14396 3056 14408
rect 2639 14368 3056 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 3050 14356 3056 14368
rect 3108 14396 3114 14408
rect 3804 14405 3832 14504
rect 4249 14501 4261 14535
rect 4295 14532 4307 14535
rect 4614 14532 4620 14544
rect 4295 14504 4620 14532
rect 4295 14501 4307 14504
rect 4249 14495 4307 14501
rect 4614 14492 4620 14504
rect 4672 14492 4678 14544
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 4764 14504 5488 14532
rect 4764 14492 4770 14504
rect 4798 14424 4804 14476
rect 4856 14464 4862 14476
rect 5460 14473 5488 14504
rect 8662 14492 8668 14544
rect 8720 14532 8726 14544
rect 9033 14535 9091 14541
rect 9033 14532 9045 14535
rect 8720 14504 9045 14532
rect 8720 14492 8726 14504
rect 9033 14501 9045 14504
rect 9079 14532 9091 14535
rect 9079 14504 12434 14532
rect 9079 14501 9091 14504
rect 9033 14495 9091 14501
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 4856 14436 5365 14464
rect 4856 14424 4862 14436
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5718 14464 5724 14476
rect 5675 14436 5724 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 10686 14464 10692 14476
rect 10275 14436 10692 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 11330 14464 11336 14476
rect 10980 14436 11336 14464
rect 3789 14399 3847 14405
rect 3108 14368 3464 14396
rect 3108 14356 3114 14368
rect 2133 14331 2191 14337
rect 2133 14297 2145 14331
rect 2179 14328 2191 14331
rect 2961 14331 3019 14337
rect 2961 14328 2973 14331
rect 2179 14300 2973 14328
rect 2179 14297 2191 14300
rect 2133 14291 2191 14297
rect 2961 14297 2973 14300
rect 3007 14297 3019 14331
rect 3436 14328 3464 14368
rect 3789 14365 3801 14399
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3936 14368 3985 14396
rect 3936 14356 3942 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4338 14356 4344 14408
rect 4396 14356 4402 14408
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 3896 14328 3924 14356
rect 3436 14300 3924 14328
rect 2961 14291 3019 14297
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 4433 14331 4491 14337
rect 4433 14328 4445 14331
rect 4120 14300 4445 14328
rect 4120 14288 4126 14300
rect 4433 14297 4445 14300
rect 4479 14297 4491 14331
rect 4908 14328 4936 14359
rect 5350 14328 5356 14340
rect 4908 14300 5356 14328
rect 4433 14291 4491 14297
rect 5350 14288 5356 14300
rect 5408 14328 5414 14340
rect 5552 14328 5580 14359
rect 5902 14356 5908 14408
rect 5960 14356 5966 14408
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14396 10103 14399
rect 10980 14396 11008 14436
rect 11330 14424 11336 14436
rect 11388 14464 11394 14476
rect 12158 14464 12164 14476
rect 11388 14436 12164 14464
rect 11388 14424 11394 14436
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12406 14464 12434 14504
rect 12986 14492 12992 14544
rect 13044 14492 13050 14544
rect 16393 14535 16451 14541
rect 16393 14532 16405 14535
rect 13556 14504 16405 14532
rect 13556 14464 13584 14504
rect 16393 14501 16405 14504
rect 16439 14501 16451 14535
rect 24596 14532 24624 14572
rect 25038 14560 25044 14572
rect 25096 14560 25102 14612
rect 25498 14560 25504 14612
rect 25556 14560 25562 14612
rect 26789 14603 26847 14609
rect 26789 14569 26801 14603
rect 26835 14600 26847 14603
rect 26970 14600 26976 14612
rect 26835 14572 26976 14600
rect 26835 14569 26847 14572
rect 26789 14563 26847 14569
rect 26970 14560 26976 14572
rect 27028 14560 27034 14612
rect 29822 14600 29828 14612
rect 29196 14572 29828 14600
rect 16393 14495 16451 14501
rect 23860 14504 24624 14532
rect 24673 14535 24731 14541
rect 12406 14436 13584 14464
rect 13630 14424 13636 14476
rect 13688 14424 13694 14476
rect 10091 14368 11008 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 12618 14396 12624 14408
rect 11112 14368 12624 14396
rect 11112 14356 11118 14368
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14396 13415 14399
rect 13814 14396 13820 14408
rect 13403 14368 13820 14396
rect 13403 14365 13415 14368
rect 13357 14359 13415 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 13906 14356 13912 14408
rect 13964 14396 13970 14408
rect 16206 14396 16212 14408
rect 13964 14368 16212 14396
rect 13964 14356 13970 14368
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16408 14396 16436 14495
rect 18782 14424 18788 14476
rect 18840 14424 18846 14476
rect 23474 14424 23480 14476
rect 23532 14464 23538 14476
rect 23860 14464 23888 14504
rect 24673 14501 24685 14535
rect 24719 14532 24731 14535
rect 25222 14532 25228 14544
rect 24719 14504 25228 14532
rect 24719 14501 24731 14504
rect 24673 14495 24731 14501
rect 25222 14492 25228 14504
rect 25280 14492 25286 14544
rect 24762 14464 24768 14476
rect 23532 14436 23888 14464
rect 23532 14424 23538 14436
rect 16574 14396 16580 14408
rect 16408 14368 16580 14396
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 19058 14356 19064 14408
rect 19116 14356 19122 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19208 14368 19809 14396
rect 19208 14356 19214 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22094 14396 22100 14408
rect 21867 14368 22100 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 22094 14356 22100 14368
rect 22152 14396 22158 14408
rect 23860 14405 23888 14436
rect 24228 14436 24768 14464
rect 24228 14408 24256 14436
rect 24762 14424 24768 14436
rect 24820 14464 24826 14476
rect 24857 14467 24915 14473
rect 24857 14464 24869 14467
rect 24820 14436 24869 14464
rect 24820 14424 24826 14436
rect 24857 14433 24869 14436
rect 24903 14433 24915 14467
rect 24857 14427 24915 14433
rect 25038 14424 25044 14476
rect 25096 14424 25102 14476
rect 26878 14424 26884 14476
rect 26936 14424 26942 14476
rect 27157 14467 27215 14473
rect 27157 14433 27169 14467
rect 27203 14464 27215 14467
rect 27614 14464 27620 14476
rect 27203 14436 27620 14464
rect 27203 14433 27215 14436
rect 27157 14427 27215 14433
rect 27614 14424 27620 14436
rect 27672 14424 27678 14476
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22152 14368 22845 14396
rect 22152 14356 22158 14368
rect 22833 14365 22845 14368
rect 22879 14396 22891 14399
rect 23845 14399 23903 14405
rect 22879 14368 23704 14396
rect 22879 14365 22891 14368
rect 22833 14359 22891 14365
rect 5408 14300 5580 14328
rect 5408 14288 5414 14300
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2682 14260 2688 14272
rect 1995 14232 2688 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 3881 14263 3939 14269
rect 3881 14260 3893 14263
rect 3384 14232 3893 14260
rect 3384 14220 3390 14232
rect 3881 14229 3893 14232
rect 3927 14229 3939 14263
rect 5552 14260 5580 14300
rect 6178 14288 6184 14340
rect 6236 14288 6242 14340
rect 7466 14328 7472 14340
rect 7406 14300 7472 14328
rect 7466 14288 7472 14300
rect 7524 14288 7530 14340
rect 9953 14331 10011 14337
rect 9953 14297 9965 14331
rect 9999 14328 10011 14331
rect 10502 14328 10508 14340
rect 9999 14300 10508 14328
rect 9999 14297 10011 14300
rect 9953 14291 10011 14297
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 12802 14288 12808 14340
rect 12860 14328 12866 14340
rect 12897 14331 12955 14337
rect 12897 14328 12909 14331
rect 12860 14300 12909 14328
rect 12860 14288 12866 14300
rect 12897 14297 12909 14300
rect 12943 14328 12955 14331
rect 14182 14328 14188 14340
rect 12943 14300 14188 14328
rect 12943 14297 12955 14300
rect 12897 14291 12955 14297
rect 14182 14288 14188 14300
rect 14240 14288 14246 14340
rect 15289 14331 15347 14337
rect 15289 14297 15301 14331
rect 15335 14328 15347 14331
rect 16942 14328 16948 14340
rect 15335 14300 16948 14328
rect 15335 14297 15347 14300
rect 15289 14291 15347 14297
rect 16942 14288 16948 14300
rect 17000 14288 17006 14340
rect 18138 14288 18144 14340
rect 18196 14288 18202 14340
rect 21082 14288 21088 14340
rect 21140 14328 21146 14340
rect 21140 14300 21220 14328
rect 21140 14288 21146 14300
rect 7650 14260 7656 14272
rect 5552 14232 7656 14260
rect 3881 14223 3939 14229
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 10413 14263 10471 14269
rect 10413 14260 10425 14263
rect 10284 14232 10425 14260
rect 10284 14220 10290 14232
rect 10413 14229 10425 14232
rect 10459 14229 10471 14263
rect 10413 14223 10471 14229
rect 13446 14220 13452 14272
rect 13504 14220 13510 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 14734 14260 14740 14272
rect 13688 14232 14740 14260
rect 13688 14220 13694 14232
rect 14734 14220 14740 14232
rect 14792 14260 14798 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14792 14232 15025 14260
rect 14792 14220 14798 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 16761 14263 16819 14269
rect 16761 14229 16773 14263
rect 16807 14260 16819 14263
rect 17034 14260 17040 14272
rect 16807 14232 17040 14260
rect 16807 14229 16819 14232
rect 16761 14223 16819 14229
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 17770 14220 17776 14272
rect 17828 14260 17834 14272
rect 18690 14260 18696 14272
rect 17828 14232 18696 14260
rect 17828 14220 17834 14232
rect 18690 14220 18696 14232
rect 18748 14260 18754 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 18748 14232 19257 14260
rect 18748 14220 18754 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 21192 14260 21220 14300
rect 21542 14288 21548 14340
rect 21600 14288 21606 14340
rect 23566 14288 23572 14340
rect 23624 14288 23630 14340
rect 23676 14328 23704 14368
rect 23845 14365 23857 14399
rect 23891 14365 23903 14399
rect 23845 14359 23903 14365
rect 23937 14399 23995 14405
rect 23937 14365 23949 14399
rect 23983 14396 23995 14399
rect 24026 14396 24032 14408
rect 23983 14368 24032 14396
rect 23983 14365 23995 14368
rect 23937 14359 23995 14365
rect 24026 14356 24032 14368
rect 24084 14356 24090 14408
rect 24210 14356 24216 14408
rect 24268 14356 24274 14408
rect 24302 14356 24308 14408
rect 24360 14396 24366 14408
rect 24397 14399 24455 14405
rect 24397 14396 24409 14399
rect 24360 14368 24409 14396
rect 24360 14356 24366 14368
rect 24397 14365 24409 14368
rect 24443 14365 24455 14399
rect 26234 14396 26240 14408
rect 24397 14359 24455 14365
rect 24504 14368 26240 14396
rect 24504 14328 24532 14368
rect 26234 14356 26240 14368
rect 26292 14356 26298 14408
rect 26510 14356 26516 14408
rect 26568 14356 26574 14408
rect 29196 14405 29224 14572
rect 29822 14560 29828 14572
rect 29880 14560 29886 14612
rect 30834 14560 30840 14612
rect 30892 14600 30898 14612
rect 33229 14603 33287 14609
rect 33229 14600 33241 14603
rect 30892 14572 33241 14600
rect 30892 14560 30898 14572
rect 33229 14569 33241 14572
rect 33275 14569 33287 14603
rect 33229 14563 33287 14569
rect 34514 14560 34520 14612
rect 34572 14600 34578 14612
rect 34793 14603 34851 14609
rect 34793 14600 34805 14603
rect 34572 14572 34805 14600
rect 34572 14560 34578 14572
rect 34793 14569 34805 14572
rect 34839 14569 34851 14603
rect 34793 14563 34851 14569
rect 35253 14603 35311 14609
rect 35253 14569 35265 14603
rect 35299 14600 35311 14603
rect 35434 14600 35440 14612
rect 35299 14572 35440 14600
rect 35299 14569 35311 14572
rect 35253 14563 35311 14569
rect 35434 14560 35440 14572
rect 35492 14560 35498 14612
rect 30926 14492 30932 14544
rect 30984 14532 30990 14544
rect 31297 14535 31355 14541
rect 31297 14532 31309 14535
rect 30984 14504 31309 14532
rect 30984 14492 30990 14504
rect 31297 14501 31309 14504
rect 31343 14501 31355 14535
rect 31297 14495 31355 14501
rect 32858 14492 32864 14544
rect 32916 14492 32922 14544
rect 34606 14492 34612 14544
rect 34664 14532 34670 14544
rect 34885 14535 34943 14541
rect 34885 14532 34897 14535
rect 34664 14504 34897 14532
rect 34664 14492 34670 14504
rect 34885 14501 34897 14504
rect 34931 14501 34943 14535
rect 34885 14495 34943 14501
rect 36633 14535 36691 14541
rect 36633 14501 36645 14535
rect 36679 14532 36691 14535
rect 36679 14504 36860 14532
rect 36679 14501 36691 14504
rect 36633 14495 36691 14501
rect 29546 14424 29552 14476
rect 29604 14464 29610 14476
rect 30190 14464 30196 14476
rect 29604 14436 30196 14464
rect 29604 14424 29610 14436
rect 30190 14424 30196 14436
rect 30248 14464 30254 14476
rect 31481 14467 31539 14473
rect 31481 14464 31493 14467
rect 30248 14436 31493 14464
rect 30248 14424 30254 14436
rect 31481 14433 31493 14436
rect 31527 14464 31539 14467
rect 32876 14464 32904 14492
rect 31527 14436 32904 14464
rect 31527 14433 31539 14436
rect 31481 14427 31539 14433
rect 34698 14424 34704 14476
rect 34756 14424 34762 14476
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 36832 14464 36860 14504
rect 37001 14467 37059 14473
rect 37001 14464 37013 14467
rect 34848 14436 36768 14464
rect 36832 14436 37013 14464
rect 34848 14424 34854 14436
rect 36740 14408 36768 14436
rect 37001 14433 37013 14436
rect 37047 14433 37059 14467
rect 37001 14427 37059 14433
rect 29181 14399 29239 14405
rect 29181 14365 29193 14399
rect 29227 14365 29239 14399
rect 29181 14359 29239 14365
rect 29362 14356 29368 14408
rect 29420 14356 29426 14408
rect 34977 14399 35035 14405
rect 34977 14396 34989 14399
rect 34808 14368 34989 14396
rect 34808 14340 34836 14368
rect 34977 14365 34989 14368
rect 35023 14365 35035 14399
rect 34977 14359 35035 14365
rect 35066 14356 35072 14408
rect 35124 14356 35130 14408
rect 35529 14399 35587 14405
rect 35529 14365 35541 14399
rect 35575 14396 35587 14399
rect 35986 14396 35992 14408
rect 35575 14368 35992 14396
rect 35575 14365 35587 14368
rect 35529 14359 35587 14365
rect 35986 14356 35992 14368
rect 36044 14356 36050 14408
rect 36354 14356 36360 14408
rect 36412 14356 36418 14408
rect 36722 14356 36728 14408
rect 36780 14356 36786 14408
rect 23676 14300 24532 14328
rect 24670 14288 24676 14340
rect 24728 14328 24734 14340
rect 25133 14331 25191 14337
rect 25133 14328 25145 14331
rect 24728 14300 25145 14328
rect 24728 14288 24734 14300
rect 25133 14297 25145 14300
rect 25179 14297 25191 14331
rect 25133 14291 25191 14297
rect 26789 14331 26847 14337
rect 26789 14297 26801 14331
rect 26835 14328 26847 14331
rect 27062 14328 27068 14340
rect 26835 14300 27068 14328
rect 26835 14297 26847 14300
rect 26789 14291 26847 14297
rect 27062 14288 27068 14300
rect 27120 14288 27126 14340
rect 27890 14288 27896 14340
rect 27948 14288 27954 14340
rect 29273 14331 29331 14337
rect 29273 14297 29285 14331
rect 29319 14328 29331 14331
rect 29825 14331 29883 14337
rect 29825 14328 29837 14331
rect 29319 14300 29837 14328
rect 29319 14297 29331 14300
rect 29273 14291 29331 14297
rect 29825 14297 29837 14300
rect 29871 14297 29883 14331
rect 31110 14328 31116 14340
rect 31050 14300 31116 14328
rect 29825 14291 29883 14297
rect 31110 14288 31116 14300
rect 31168 14288 31174 14340
rect 31202 14288 31208 14340
rect 31260 14328 31266 14340
rect 31757 14331 31815 14337
rect 31757 14328 31769 14331
rect 31260 14300 31769 14328
rect 31260 14288 31266 14300
rect 31757 14297 31769 14300
rect 31803 14297 31815 14331
rect 31757 14291 31815 14297
rect 31956 14300 32246 14328
rect 22002 14260 22008 14272
rect 21192 14232 22008 14260
rect 19245 14223 19303 14229
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 24489 14263 24547 14269
rect 24489 14229 24501 14263
rect 24535 14260 24547 14263
rect 24946 14260 24952 14272
rect 24535 14232 24952 14260
rect 24535 14229 24547 14232
rect 24489 14223 24547 14229
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 26605 14263 26663 14269
rect 26605 14229 26617 14263
rect 26651 14260 26663 14263
rect 27522 14260 27528 14272
rect 26651 14232 27528 14260
rect 26651 14229 26663 14232
rect 26605 14223 26663 14229
rect 27522 14220 27528 14232
rect 27580 14220 27586 14272
rect 28626 14220 28632 14272
rect 28684 14220 28690 14272
rect 31128 14260 31156 14288
rect 31294 14260 31300 14272
rect 31128 14232 31300 14260
rect 31294 14220 31300 14232
rect 31352 14260 31358 14272
rect 31956 14260 31984 14300
rect 34790 14288 34796 14340
rect 34848 14288 34854 14340
rect 35437 14331 35495 14337
rect 35437 14297 35449 14331
rect 35483 14328 35495 14331
rect 36078 14328 36084 14340
rect 35483 14300 36084 14328
rect 35483 14297 35495 14300
rect 35437 14291 35495 14297
rect 36078 14288 36084 14300
rect 36136 14288 36142 14340
rect 36630 14288 36636 14340
rect 36688 14288 36694 14340
rect 37458 14288 37464 14340
rect 37516 14288 37522 14340
rect 31352 14232 31984 14260
rect 36449 14263 36507 14269
rect 31352 14220 31358 14232
rect 36449 14229 36461 14263
rect 36495 14260 36507 14263
rect 37366 14260 37372 14272
rect 36495 14232 37372 14260
rect 36495 14229 36507 14232
rect 36449 14223 36507 14229
rect 37366 14220 37372 14232
rect 37424 14220 37430 14272
rect 38473 14263 38531 14269
rect 38473 14229 38485 14263
rect 38519 14260 38531 14263
rect 38519 14232 38884 14260
rect 38519 14229 38531 14232
rect 38473 14223 38531 14229
rect 1104 14170 38824 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 38824 14170
rect 1104 14096 38824 14118
rect 3513 14059 3571 14065
rect 3513 14025 3525 14059
rect 3559 14056 3571 14059
rect 3602 14056 3608 14068
rect 3559 14028 3608 14056
rect 3559 14025 3571 14028
rect 3513 14019 3571 14025
rect 3602 14016 3608 14028
rect 3660 14056 3666 14068
rect 3970 14056 3976 14068
rect 3660 14028 3976 14056
rect 3660 14016 3666 14028
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 5350 14056 5356 14068
rect 5184 14028 5356 14056
rect 2774 13948 2780 14000
rect 2832 13948 2838 14000
rect 3694 13948 3700 14000
rect 3752 13948 3758 14000
rect 4338 13948 4344 14000
rect 4396 13988 4402 14000
rect 5184 13997 5212 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5997 14059 6055 14065
rect 5997 14025 6009 14059
rect 6043 14056 6055 14059
rect 6178 14056 6184 14068
rect 6043 14028 6184 14056
rect 6043 14025 6055 14028
rect 5997 14019 6055 14025
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 9861 14059 9919 14065
rect 9861 14025 9873 14059
rect 9907 14056 9919 14059
rect 11054 14056 11060 14068
rect 9907 14028 11060 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 12345 14059 12403 14065
rect 12345 14025 12357 14059
rect 12391 14056 12403 14059
rect 12894 14056 12900 14068
rect 12391 14028 12900 14056
rect 12391 14025 12403 14028
rect 12345 14019 12403 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 13722 14016 13728 14068
rect 13780 14016 13786 14068
rect 17678 14056 17684 14068
rect 16684 14028 17684 14056
rect 4969 13991 5027 13997
rect 4969 13988 4981 13991
rect 4396 13960 4981 13988
rect 4396 13948 4402 13960
rect 4969 13957 4981 13960
rect 5015 13988 5027 13991
rect 5169 13991 5227 13997
rect 5015 13960 5120 13988
rect 5015 13957 5027 13960
rect 4969 13951 5027 13957
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1452 13892 1777 13920
rect 1452 13880 1458 13892
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 5092 13920 5120 13960
rect 5169 13957 5181 13991
rect 5215 13957 5227 13991
rect 5169 13951 5227 13957
rect 5626 13948 5632 14000
rect 5684 13948 5690 14000
rect 5845 13991 5903 13997
rect 5845 13957 5857 13991
rect 5891 13988 5903 13991
rect 7469 13991 7527 13997
rect 7469 13988 7481 13991
rect 5891 13960 7481 13988
rect 5891 13957 5903 13960
rect 5845 13951 5903 13957
rect 7469 13957 7481 13960
rect 7515 13957 7527 13991
rect 8294 13988 8300 14000
rect 7469 13951 7527 13957
rect 8128 13960 8300 13988
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5092 13892 5273 13920
rect 1765 13883 1823 13889
rect 5261 13889 5273 13892
rect 5307 13920 5319 13923
rect 5350 13920 5356 13932
rect 5307 13892 5356 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13920 5595 13923
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 5583 13892 6377 13920
rect 5583 13889 5595 13892
rect 5537 13883 5595 13889
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 6546 13880 6552 13932
rect 6604 13920 6610 13932
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 6604 13892 7113 13920
rect 6604 13880 6610 13892
rect 7101 13889 7113 13892
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7285 13923 7343 13929
rect 7285 13889 7297 13923
rect 7331 13920 7343 13923
rect 7650 13920 7656 13932
rect 7331 13892 7656 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 8128 13929 8156 13960
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 9950 13988 9956 14000
rect 9614 13960 9956 13988
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 11241 13991 11299 13997
rect 11241 13957 11253 13991
rect 11287 13988 11299 13991
rect 11287 13960 13308 13988
rect 11287 13957 11299 13960
rect 11241 13951 11299 13957
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13889 8171 13923
rect 8113 13883 8171 13889
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 10284 13892 10333 13920
rect 10284 13880 10290 13892
rect 10321 13889 10333 13892
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 10413 13923 10471 13929
rect 10413 13889 10425 13923
rect 10459 13920 10471 13923
rect 10502 13920 10508 13932
rect 10459 13892 10508 13920
rect 10459 13889 10471 13892
rect 10413 13883 10471 13889
rect 10502 13880 10508 13892
rect 10560 13920 10566 13932
rect 10560 13892 11008 13920
rect 10560 13880 10566 13892
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 2832 13824 3985 13852
rect 2832 13812 2838 13824
rect 3973 13821 3985 13824
rect 4019 13852 4031 13855
rect 4154 13852 4160 13864
rect 4019 13824 4160 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 5000 13824 6929 13852
rect 2028 13719 2086 13725
rect 2028 13685 2040 13719
rect 2074 13716 2086 13719
rect 3326 13716 3332 13728
rect 2074 13688 3332 13716
rect 2074 13685 2086 13688
rect 2028 13679 2086 13685
rect 3326 13676 3332 13688
rect 3384 13676 3390 13728
rect 4798 13676 4804 13728
rect 4856 13676 4862 13728
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 5000 13725 5028 13824
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13821 10655 13855
rect 10980 13852 11008 13892
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 11112 13892 11161 13920
rect 11112 13880 11118 13892
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 11333 13923 11391 13929
rect 11333 13889 11345 13923
rect 11379 13920 11391 13923
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11379 13892 11713 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 11701 13889 11713 13892
rect 11747 13920 11759 13923
rect 11790 13920 11796 13932
rect 11747 13892 11796 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 11348 13852 11376 13883
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 10980 13824 11376 13852
rect 11900 13852 11928 13883
rect 12158 13880 12164 13932
rect 12216 13880 12222 13932
rect 12618 13880 12624 13932
rect 12676 13880 12682 13932
rect 12894 13880 12900 13932
rect 12952 13880 12958 13932
rect 13280 13929 13308 13960
rect 14826 13948 14832 14000
rect 14884 13948 14890 14000
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 11900 13824 12449 13852
rect 10597 13815 10655 13821
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 9953 13787 10011 13793
rect 9953 13784 9965 13787
rect 9416 13756 9965 13784
rect 4985 13719 5043 13725
rect 4985 13716 4997 13719
rect 4948 13688 4997 13716
rect 4948 13676 4954 13688
rect 4985 13685 4997 13688
rect 5031 13685 5043 13719
rect 4985 13679 5043 13685
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 5537 13719 5595 13725
rect 5537 13716 5549 13719
rect 5316 13688 5549 13716
rect 5316 13676 5322 13688
rect 5537 13685 5549 13688
rect 5583 13685 5595 13719
rect 5537 13679 5595 13685
rect 5810 13676 5816 13728
rect 5868 13676 5874 13728
rect 8376 13719 8434 13725
rect 8376 13685 8388 13719
rect 8422 13716 8434 13719
rect 9416 13716 9444 13756
rect 9953 13753 9965 13756
rect 9999 13753 10011 13787
rect 9953 13747 10011 13753
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10612 13784 10640 13815
rect 12986 13812 12992 13864
rect 13044 13852 13050 13864
rect 13096 13852 13124 13883
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 13412 13892 13553 13920
rect 13412 13880 13418 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13449 13855 13507 13861
rect 13449 13852 13461 13855
rect 13044 13824 13461 13852
rect 13044 13812 13050 13824
rect 13449 13821 13461 13824
rect 13495 13821 13507 13855
rect 13449 13815 13507 13821
rect 15470 13812 15476 13864
rect 15528 13812 15534 13864
rect 15746 13812 15752 13864
rect 15804 13812 15810 13864
rect 16684 13861 16712 14028
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 17770 14016 17776 14068
rect 17828 14016 17834 14068
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18874 14056 18880 14068
rect 18012 14028 18880 14056
rect 18012 14016 18018 14028
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 19702 14016 19708 14068
rect 19760 14016 19766 14068
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 20717 14059 20775 14065
rect 20220 14028 20392 14056
rect 20220 14016 20226 14028
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 17236 13960 18245 13988
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13920 17003 13923
rect 17034 13920 17040 13932
rect 16991 13892 17040 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 17034 13880 17040 13892
rect 17092 13920 17098 13932
rect 17236 13929 17264 13960
rect 18233 13957 18245 13960
rect 18279 13957 18291 13991
rect 18233 13951 18291 13957
rect 19245 13991 19303 13997
rect 19245 13957 19257 13991
rect 19291 13988 19303 13991
rect 19334 13988 19340 14000
rect 19291 13960 19340 13988
rect 19291 13957 19303 13960
rect 19245 13951 19303 13957
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 19426 13948 19432 14000
rect 19484 13997 19490 14000
rect 19484 13991 19503 13997
rect 19491 13957 19503 13991
rect 19484 13951 19503 13957
rect 19484 13948 19490 13951
rect 17221 13923 17279 13929
rect 17092 13892 17172 13920
rect 17092 13880 17098 13892
rect 16669 13855 16727 13861
rect 16669 13821 16681 13855
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 10100 13756 12434 13784
rect 10100 13744 10106 13756
rect 8422 13688 9444 13716
rect 12406 13728 12434 13756
rect 13354 13744 13360 13796
rect 13412 13744 13418 13796
rect 17144 13784 17172 13892
rect 17221 13889 17233 13923
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 17911 13892 18092 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 17880 13852 17908 13883
rect 17644 13824 17908 13852
rect 17644 13812 17650 13824
rect 17954 13812 17960 13864
rect 18012 13812 18018 13864
rect 18064 13852 18092 13892
rect 18690 13880 18696 13932
rect 18748 13920 18754 13932
rect 18969 13923 19027 13929
rect 18969 13920 18981 13923
rect 18748 13892 18981 13920
rect 18748 13880 18754 13892
rect 18969 13889 18981 13892
rect 19015 13889 19027 13923
rect 18969 13883 19027 13889
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13920 19211 13923
rect 19720 13920 19748 14016
rect 20254 13988 20260 14000
rect 19904 13960 20260 13988
rect 19904 13929 19932 13960
rect 20254 13948 20260 13960
rect 20312 13948 20318 14000
rect 20364 13997 20392 14028
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 21542 14056 21548 14068
rect 20763 14028 21548 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 24302 14016 24308 14068
rect 24360 14056 24366 14068
rect 24489 14059 24547 14065
rect 24489 14056 24501 14059
rect 24360 14028 24501 14056
rect 24360 14016 24366 14028
rect 24489 14025 24501 14028
rect 24535 14025 24547 14059
rect 24489 14019 24547 14025
rect 24762 14016 24768 14068
rect 24820 14056 24826 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 24820 14028 25053 14056
rect 24820 14016 24826 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 27062 14016 27068 14068
rect 27120 14016 27126 14068
rect 27522 14016 27528 14068
rect 27580 14056 27586 14068
rect 27709 14059 27767 14065
rect 27709 14056 27721 14059
rect 27580 14028 27721 14056
rect 27580 14016 27586 14028
rect 27709 14025 27721 14028
rect 27755 14025 27767 14059
rect 27709 14019 27767 14025
rect 29362 14016 29368 14068
rect 29420 14056 29426 14068
rect 30285 14059 30343 14065
rect 30285 14056 30297 14059
rect 29420 14028 30297 14056
rect 29420 14016 29426 14028
rect 30285 14025 30297 14028
rect 30331 14025 30343 14059
rect 30285 14019 30343 14025
rect 31018 14016 31024 14068
rect 31076 14016 31082 14068
rect 31202 14016 31208 14068
rect 31260 14016 31266 14068
rect 32953 14059 33011 14065
rect 32953 14025 32965 14059
rect 32999 14056 33011 14059
rect 33689 14059 33747 14065
rect 33689 14056 33701 14059
rect 32999 14028 33701 14056
rect 32999 14025 33011 14028
rect 32953 14019 33011 14025
rect 33689 14025 33701 14028
rect 33735 14025 33747 14059
rect 33689 14019 33747 14025
rect 35329 14059 35387 14065
rect 35329 14025 35341 14059
rect 35375 14056 35387 14059
rect 35986 14056 35992 14068
rect 35375 14028 35992 14056
rect 35375 14025 35387 14028
rect 35329 14019 35387 14025
rect 35986 14016 35992 14028
rect 36044 14016 36050 14068
rect 36630 14016 36636 14068
rect 36688 14056 36694 14068
rect 36817 14059 36875 14065
rect 36817 14056 36829 14059
rect 36688 14028 36829 14056
rect 36688 14016 36694 14028
rect 36817 14025 36829 14028
rect 36863 14025 36875 14059
rect 36817 14019 36875 14025
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 37553 14059 37611 14065
rect 37553 14056 37565 14059
rect 37424 14028 37565 14056
rect 37424 14016 37430 14028
rect 37553 14025 37565 14028
rect 37599 14025 37611 14059
rect 37553 14019 37611 14025
rect 20349 13991 20407 13997
rect 20349 13957 20361 13991
rect 20395 13957 20407 13991
rect 20349 13951 20407 13957
rect 20565 13991 20623 13997
rect 20565 13957 20577 13991
rect 20611 13988 20623 13991
rect 20901 13991 20959 13997
rect 20901 13988 20913 13991
rect 20611 13960 20913 13988
rect 20611 13957 20623 13960
rect 20565 13951 20623 13957
rect 20901 13957 20913 13960
rect 20947 13957 20959 13991
rect 22094 13988 22100 14000
rect 20901 13951 20959 13957
rect 21836 13960 22100 13988
rect 19199 13892 19748 13920
rect 19889 13923 19947 13929
rect 19199 13889 19211 13892
rect 19153 13883 19211 13889
rect 19889 13889 19901 13923
rect 19935 13889 19947 13923
rect 19889 13883 19947 13889
rect 19978 13880 19984 13932
rect 20036 13880 20042 13932
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13920 20223 13923
rect 20438 13920 20444 13932
rect 20211 13892 20444 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 21836 13929 21864 13960
rect 22094 13948 22100 13960
rect 22152 13948 22158 14000
rect 23842 13988 23848 14000
rect 23322 13960 23848 13988
rect 23842 13948 23848 13960
rect 23900 13948 23906 14000
rect 24320 13988 24348 14016
rect 24044 13960 24348 13988
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13889 21051 13923
rect 20993 13883 21051 13889
rect 21821 13923 21879 13929
rect 21821 13889 21833 13923
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 18064 13824 18797 13852
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19518 13852 19524 13864
rect 19107 13824 19524 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19518 13812 19524 13824
rect 19576 13812 19582 13864
rect 19610 13812 19616 13864
rect 19668 13852 19674 13864
rect 21008 13852 21036 13883
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24044 13929 24072 13960
rect 24670 13948 24676 14000
rect 24728 13988 24734 14000
rect 24728 13960 24992 13988
rect 24728 13948 24734 13960
rect 24964 13929 24992 13960
rect 29822 13948 29828 14000
rect 29880 13948 29886 14000
rect 33137 13991 33195 13997
rect 29932 13960 30144 13988
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 23532 13892 23765 13920
rect 23532 13880 23538 13892
rect 23753 13889 23765 13892
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 24029 13923 24087 13929
rect 24029 13889 24041 13923
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 24121 13883 24179 13889
rect 24213 13923 24271 13929
rect 24213 13889 24225 13923
rect 24259 13920 24271 13923
rect 24397 13923 24455 13929
rect 24397 13920 24409 13923
rect 24259 13892 24409 13920
rect 24259 13889 24271 13892
rect 24213 13883 24271 13889
rect 24397 13889 24409 13892
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13889 25007 13923
rect 24949 13883 25007 13889
rect 19668 13824 21036 13852
rect 19668 13812 19674 13824
rect 22094 13812 22100 13864
rect 22152 13812 22158 13864
rect 23768 13852 23796 13883
rect 24136 13852 24164 13883
rect 26694 13880 26700 13932
rect 26752 13920 26758 13932
rect 27341 13923 27399 13929
rect 27341 13920 27353 13923
rect 26752 13892 27353 13920
rect 26752 13880 26758 13892
rect 27341 13889 27353 13892
rect 27387 13920 27399 13923
rect 28353 13923 28411 13929
rect 28353 13920 28365 13923
rect 27387 13892 28365 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 28353 13889 28365 13892
rect 28399 13920 28411 13923
rect 28626 13920 28632 13932
rect 28399 13892 28632 13920
rect 28399 13889 28411 13892
rect 28353 13883 28411 13889
rect 28626 13880 28632 13892
rect 28684 13880 28690 13932
rect 24854 13852 24860 13864
rect 23768 13824 24164 13852
rect 24688 13824 24860 13852
rect 17972 13784 18000 13812
rect 20073 13787 20131 13793
rect 20073 13784 20085 13787
rect 17144 13756 18000 13784
rect 19444 13756 20085 13784
rect 12406 13688 12440 13728
rect 8422 13685 8434 13688
rect 8376 13679 8434 13685
rect 12434 13676 12440 13688
rect 12492 13716 12498 13728
rect 13170 13716 13176 13728
rect 12492 13688 13176 13716
rect 12492 13676 12498 13688
rect 13170 13676 13176 13688
rect 13228 13716 13234 13728
rect 13630 13716 13636 13728
rect 13228 13688 13636 13716
rect 13228 13676 13234 13688
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 13998 13676 14004 13728
rect 14056 13676 14062 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 16761 13719 16819 13725
rect 16761 13716 16773 13719
rect 16632 13688 16773 13716
rect 16632 13676 16638 13688
rect 16761 13685 16773 13688
rect 16807 13685 16819 13719
rect 16761 13679 16819 13685
rect 16853 13719 16911 13725
rect 16853 13685 16865 13719
rect 16899 13716 16911 13719
rect 17129 13719 17187 13725
rect 17129 13716 17141 13719
rect 16899 13688 17141 13716
rect 16899 13685 16911 13688
rect 16853 13679 16911 13685
rect 17129 13685 17141 13688
rect 17175 13685 17187 13719
rect 17129 13679 17187 13685
rect 17402 13676 17408 13728
rect 17460 13676 17466 13728
rect 19444 13725 19472 13756
rect 20073 13753 20085 13756
rect 20119 13784 20131 13787
rect 20714 13784 20720 13796
rect 20119 13756 20720 13784
rect 20119 13753 20131 13756
rect 20073 13747 20131 13753
rect 20714 13744 20720 13756
rect 20772 13744 20778 13796
rect 23753 13787 23811 13793
rect 23753 13753 23765 13787
rect 23799 13784 23811 13787
rect 23934 13784 23940 13796
rect 23799 13756 23940 13784
rect 23799 13753 23811 13756
rect 23753 13747 23811 13753
rect 23934 13744 23940 13756
rect 23992 13744 23998 13796
rect 24688 13793 24716 13824
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 27065 13855 27123 13861
rect 27065 13821 27077 13855
rect 27111 13852 27123 13855
rect 27798 13852 27804 13864
rect 27111 13824 27804 13852
rect 27111 13821 27123 13824
rect 27065 13815 27123 13821
rect 27798 13812 27804 13824
rect 27856 13852 27862 13864
rect 28534 13852 28540 13864
rect 27856 13824 28540 13852
rect 27856 13812 27862 13824
rect 28534 13812 28540 13824
rect 28592 13852 28598 13864
rect 29932 13852 29960 13960
rect 30009 13923 30067 13929
rect 30009 13889 30021 13923
rect 30055 13889 30067 13923
rect 30009 13883 30067 13889
rect 28592 13824 29960 13852
rect 28592 13812 28598 13824
rect 24673 13787 24731 13793
rect 24673 13753 24685 13787
rect 24719 13753 24731 13787
rect 24673 13747 24731 13753
rect 26510 13744 26516 13796
rect 26568 13784 26574 13796
rect 27249 13787 27307 13793
rect 27249 13784 27261 13787
rect 26568 13756 27261 13784
rect 26568 13744 26574 13756
rect 27249 13753 27261 13756
rect 27295 13784 27307 13787
rect 28166 13784 28172 13796
rect 27295 13756 28172 13784
rect 27295 13753 27307 13756
rect 27249 13747 27307 13753
rect 28166 13744 28172 13756
rect 28224 13744 28230 13796
rect 30024 13784 30052 13883
rect 30116 13852 30144 13960
rect 33137 13957 33149 13991
rect 33183 13988 33195 13991
rect 33229 13991 33287 13997
rect 33229 13988 33241 13991
rect 33183 13960 33241 13988
rect 33183 13957 33195 13960
rect 33137 13951 33195 13957
rect 33229 13957 33241 13960
rect 33275 13957 33287 13991
rect 33229 13951 33287 13957
rect 34606 13948 34612 14000
rect 34664 13988 34670 14000
rect 35529 13991 35587 13997
rect 35529 13988 35541 13991
rect 34664 13960 35541 13988
rect 34664 13948 34670 13960
rect 35529 13957 35541 13960
rect 35575 13988 35587 13991
rect 35897 13991 35955 13997
rect 35897 13988 35909 13991
rect 35575 13960 35909 13988
rect 35575 13957 35587 13960
rect 35529 13951 35587 13957
rect 35897 13957 35909 13960
rect 35943 13957 35955 13991
rect 35897 13951 35955 13957
rect 36265 13991 36323 13997
rect 36265 13957 36277 13991
rect 36311 13988 36323 13991
rect 36354 13988 36360 14000
rect 36311 13960 36360 13988
rect 36311 13957 36323 13960
rect 36265 13951 36323 13957
rect 30193 13923 30251 13929
rect 30193 13889 30205 13923
rect 30239 13920 30251 13923
rect 30561 13923 30619 13929
rect 30561 13920 30573 13923
rect 30239 13892 30573 13920
rect 30239 13889 30251 13892
rect 30193 13883 30251 13889
rect 30561 13889 30573 13892
rect 30607 13920 30619 13923
rect 30926 13920 30932 13932
rect 30607 13892 30932 13920
rect 30607 13889 30619 13892
rect 30561 13883 30619 13889
rect 30926 13880 30932 13892
rect 30984 13880 30990 13932
rect 31573 13923 31631 13929
rect 31573 13889 31585 13923
rect 31619 13920 31631 13923
rect 31662 13920 31668 13932
rect 31619 13892 31668 13920
rect 31619 13889 31631 13892
rect 31573 13883 31631 13889
rect 31662 13880 31668 13892
rect 31720 13920 31726 13932
rect 32861 13923 32919 13929
rect 32861 13920 32873 13923
rect 31720 13892 32873 13920
rect 31720 13880 31726 13892
rect 32861 13889 32873 13892
rect 32907 13920 32919 13923
rect 33413 13923 33471 13929
rect 33413 13920 33425 13923
rect 32907 13892 33425 13920
rect 32907 13889 32919 13892
rect 32861 13883 32919 13889
rect 33413 13889 33425 13892
rect 33459 13889 33471 13923
rect 33413 13883 33471 13889
rect 33502 13880 33508 13932
rect 33560 13920 33566 13932
rect 34241 13923 34299 13929
rect 34241 13920 34253 13923
rect 33560 13892 34253 13920
rect 33560 13880 33566 13892
rect 34241 13889 34253 13892
rect 34287 13889 34299 13923
rect 35434 13920 35440 13932
rect 34241 13883 34299 13889
rect 35084 13892 35440 13920
rect 35084 13864 35112 13892
rect 35434 13880 35440 13892
rect 35492 13920 35498 13932
rect 35713 13923 35771 13929
rect 35713 13920 35725 13923
rect 35492 13892 35725 13920
rect 35492 13880 35498 13892
rect 35713 13889 35725 13892
rect 35759 13889 35771 13923
rect 35713 13883 35771 13889
rect 30285 13855 30343 13861
rect 30285 13852 30297 13855
rect 30116 13824 30297 13852
rect 30285 13821 30297 13824
rect 30331 13821 30343 13855
rect 33229 13855 33287 13861
rect 33229 13852 33241 13855
rect 30285 13815 30343 13821
rect 32784 13824 33241 13852
rect 30300 13784 30328 13815
rect 30024 13756 30236 13784
rect 30300 13756 30604 13784
rect 30208 13728 30236 13756
rect 19429 13719 19487 13725
rect 19429 13685 19441 13719
rect 19475 13685 19487 13719
rect 19429 13679 19487 13685
rect 19610 13676 19616 13728
rect 19668 13676 19674 13728
rect 20530 13676 20536 13728
rect 20588 13676 20594 13728
rect 23569 13719 23627 13725
rect 23569 13685 23581 13719
rect 23615 13716 23627 13719
rect 23658 13716 23664 13728
rect 23615 13688 23664 13716
rect 23615 13685 23627 13688
rect 23569 13679 23627 13685
rect 23658 13676 23664 13688
rect 23716 13676 23722 13728
rect 24857 13719 24915 13725
rect 24857 13685 24869 13719
rect 24903 13716 24915 13719
rect 24946 13716 24952 13728
rect 24903 13688 24952 13716
rect 24903 13685 24915 13688
rect 24857 13679 24915 13685
rect 24946 13676 24952 13688
rect 25004 13676 25010 13728
rect 30190 13676 30196 13728
rect 30248 13716 30254 13728
rect 30469 13719 30527 13725
rect 30469 13716 30481 13719
rect 30248 13688 30481 13716
rect 30248 13676 30254 13688
rect 30469 13685 30481 13688
rect 30515 13685 30527 13719
rect 30576 13716 30604 13756
rect 30650 13744 30656 13796
rect 30708 13744 30714 13796
rect 31754 13784 31760 13796
rect 31036 13756 31760 13784
rect 31036 13725 31064 13756
rect 31754 13744 31760 13756
rect 31812 13784 31818 13796
rect 32784 13784 32812 13824
rect 33229 13821 33241 13824
rect 33275 13852 33287 13855
rect 35066 13852 35072 13864
rect 33275 13824 35072 13852
rect 33275 13821 33287 13824
rect 33229 13815 33287 13821
rect 35066 13812 35072 13824
rect 35124 13812 35130 13864
rect 35912 13852 35940 13951
rect 36354 13948 36360 13960
rect 36412 13988 36418 14000
rect 36412 13960 37044 13988
rect 36412 13948 36418 13960
rect 35986 13880 35992 13932
rect 36044 13880 36050 13932
rect 36078 13880 36084 13932
rect 36136 13920 36142 13932
rect 37016 13929 37044 13960
rect 37001 13923 37059 13929
rect 36136 13892 36952 13920
rect 36136 13880 36142 13892
rect 36817 13855 36875 13861
rect 36817 13852 36829 13855
rect 35912 13824 36829 13852
rect 36817 13821 36829 13824
rect 36863 13821 36875 13855
rect 36924 13852 36952 13892
rect 37001 13889 37013 13923
rect 37047 13889 37059 13923
rect 37001 13883 37059 13889
rect 37093 13923 37151 13929
rect 37093 13889 37105 13923
rect 37139 13920 37151 13923
rect 38197 13923 38255 13929
rect 38197 13920 38209 13923
rect 37139 13892 38209 13920
rect 37139 13889 37151 13892
rect 37093 13883 37151 13889
rect 38197 13889 38209 13892
rect 38243 13920 38255 13923
rect 38856 13920 38884 14232
rect 38243 13892 38884 13920
rect 38243 13889 38255 13892
rect 38197 13883 38255 13889
rect 37108 13852 37136 13883
rect 36924 13824 37136 13852
rect 36817 13815 36875 13821
rect 31812 13756 32812 13784
rect 36832 13784 36860 13815
rect 37274 13784 37280 13796
rect 36832 13756 37280 13784
rect 31812 13744 31818 13756
rect 37274 13744 37280 13756
rect 37332 13744 37338 13796
rect 31021 13719 31079 13725
rect 31021 13716 31033 13719
rect 30576 13688 31033 13716
rect 30469 13679 30527 13685
rect 31021 13685 31033 13688
rect 31067 13685 31079 13719
rect 31021 13679 31079 13685
rect 31481 13719 31539 13725
rect 31481 13685 31493 13719
rect 31527 13716 31539 13719
rect 31570 13716 31576 13728
rect 31527 13688 31576 13716
rect 31527 13685 31539 13688
rect 31481 13679 31539 13685
rect 31570 13676 31576 13688
rect 31628 13676 31634 13728
rect 32858 13676 32864 13728
rect 32916 13716 32922 13728
rect 33137 13719 33195 13725
rect 33137 13716 33149 13719
rect 32916 13688 33149 13716
rect 32916 13676 32922 13688
rect 33137 13685 33149 13688
rect 33183 13685 33195 13719
rect 33137 13679 33195 13685
rect 34698 13676 34704 13728
rect 34756 13716 34762 13728
rect 35161 13719 35219 13725
rect 35161 13716 35173 13719
rect 34756 13688 35173 13716
rect 34756 13676 34762 13688
rect 35161 13685 35173 13688
rect 35207 13685 35219 13719
rect 35161 13679 35219 13685
rect 35345 13719 35403 13725
rect 35345 13685 35357 13719
rect 35391 13716 35403 13719
rect 35434 13716 35440 13728
rect 35391 13688 35440 13716
rect 35391 13685 35403 13688
rect 35345 13679 35403 13685
rect 35434 13676 35440 13688
rect 35492 13676 35498 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3789 13515 3847 13521
rect 2832 13484 3648 13512
rect 2832 13472 2838 13484
rect 1854 13336 1860 13388
rect 1912 13376 1918 13388
rect 2317 13379 2375 13385
rect 2317 13376 2329 13379
rect 1912 13348 2329 13376
rect 1912 13336 1918 13348
rect 2317 13345 2329 13348
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 2332 13172 2360 13339
rect 2774 13336 2780 13388
rect 2832 13336 2838 13388
rect 3620 13385 3648 13484
rect 3789 13481 3801 13515
rect 3835 13512 3847 13515
rect 3878 13512 3884 13524
rect 3835 13484 3884 13512
rect 3835 13481 3847 13484
rect 3789 13475 3847 13481
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 3970 13472 3976 13524
rect 4028 13472 4034 13524
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 5040 13484 6101 13512
rect 5040 13472 5046 13484
rect 6089 13481 6101 13484
rect 6135 13481 6147 13515
rect 6089 13475 6147 13481
rect 12986 13472 12992 13524
rect 13044 13472 13050 13524
rect 13354 13472 13360 13524
rect 13412 13472 13418 13524
rect 15289 13515 15347 13521
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 15470 13512 15476 13524
rect 15335 13484 15476 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 17586 13521 17592 13524
rect 17543 13515 17592 13521
rect 17543 13481 17555 13515
rect 17589 13481 17592 13515
rect 17543 13475 17592 13481
rect 17586 13472 17592 13475
rect 17644 13472 17650 13524
rect 17678 13472 17684 13524
rect 17736 13512 17742 13524
rect 19337 13515 19395 13521
rect 19337 13512 19349 13515
rect 17736 13484 19349 13512
rect 17736 13472 17742 13484
rect 19337 13481 19349 13484
rect 19383 13512 19395 13515
rect 19426 13512 19432 13524
rect 19383 13484 19432 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19426 13472 19432 13484
rect 19484 13512 19490 13524
rect 20162 13512 20168 13524
rect 19484 13484 20168 13512
rect 19484 13472 19490 13484
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 20625 13515 20683 13521
rect 20625 13481 20637 13515
rect 20671 13512 20683 13515
rect 20714 13512 20720 13524
rect 20671 13484 20720 13512
rect 20671 13481 20683 13484
rect 20625 13475 20683 13481
rect 20714 13472 20720 13484
rect 20772 13512 20778 13524
rect 21082 13512 21088 13524
rect 20772 13484 21088 13512
rect 20772 13472 20778 13484
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 21910 13472 21916 13524
rect 21968 13472 21974 13524
rect 22094 13472 22100 13524
rect 22152 13472 22158 13524
rect 23477 13515 23535 13521
rect 23477 13481 23489 13515
rect 23523 13512 23535 13515
rect 24946 13512 24952 13524
rect 23523 13484 24952 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 24946 13472 24952 13484
rect 25004 13472 25010 13524
rect 25222 13472 25228 13524
rect 25280 13472 25286 13524
rect 29822 13472 29828 13524
rect 29880 13512 29886 13524
rect 31294 13512 31300 13524
rect 29880 13484 31300 13512
rect 29880 13472 29886 13484
rect 31294 13472 31300 13484
rect 31352 13472 31358 13524
rect 35986 13472 35992 13524
rect 36044 13512 36050 13524
rect 36170 13512 36176 13524
rect 36044 13484 36176 13512
rect 36044 13472 36050 13484
rect 36170 13472 36176 13484
rect 36228 13512 36234 13524
rect 36449 13515 36507 13521
rect 36449 13512 36461 13515
rect 36228 13484 36461 13512
rect 36228 13472 36234 13484
rect 36449 13481 36461 13484
rect 36495 13481 36507 13515
rect 36449 13475 36507 13481
rect 7837 13447 7895 13453
rect 7837 13413 7849 13447
rect 7883 13444 7895 13447
rect 9214 13444 9220 13456
rect 7883 13416 9220 13444
rect 7883 13413 7895 13416
rect 7837 13407 7895 13413
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 13633 13447 13691 13453
rect 13633 13413 13645 13447
rect 13679 13444 13691 13447
rect 13722 13444 13728 13456
rect 13679 13416 13728 13444
rect 13679 13413 13691 13416
rect 13633 13407 13691 13413
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 21269 13447 21327 13453
rect 21269 13444 21281 13447
rect 20088 13416 21281 13444
rect 3605 13379 3663 13385
rect 3605 13345 3617 13379
rect 3651 13376 3663 13379
rect 4614 13376 4620 13388
rect 3651 13348 4620 13376
rect 3651 13345 3663 13348
rect 3605 13339 3663 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 7392 13348 7941 13376
rect 7392 13320 7420 13348
rect 7929 13345 7941 13348
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13376 9459 13379
rect 10042 13376 10048 13388
rect 9447 13348 10048 13376
rect 9447 13345 9459 13348
rect 9401 13339 9459 13345
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 11793 13379 11851 13385
rect 11793 13345 11805 13379
rect 11839 13376 11851 13379
rect 12342 13376 12348 13388
rect 11839 13348 12348 13376
rect 11839 13345 11851 13348
rect 11793 13339 11851 13345
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 12434 13336 12440 13388
rect 12492 13336 12498 13388
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12676 13348 12817 13376
rect 12676 13336 12682 13348
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 13446 13376 13452 13388
rect 12805 13339 12863 13345
rect 12912 13348 13452 13376
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2455 13280 2973 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 2961 13271 3019 13277
rect 3620 13280 4353 13308
rect 2498 13200 2504 13252
rect 2556 13240 2562 13252
rect 3620 13240 3648 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 8478 13308 8484 13320
rect 7607 13280 8484 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 10226 13308 10232 13320
rect 9539 13280 10232 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13308 12311 13311
rect 12526 13308 12532 13320
rect 12299 13280 12532 13308
rect 12299 13277 12311 13280
rect 12253 13271 12311 13277
rect 12526 13268 12532 13280
rect 12584 13308 12590 13320
rect 12912 13308 12940 13348
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 14734 13336 14740 13388
rect 14792 13336 14798 13388
rect 15746 13336 15752 13388
rect 15804 13336 15810 13388
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13376 16175 13379
rect 16574 13376 16580 13388
rect 16163 13348 16580 13376
rect 16163 13345 16175 13348
rect 16117 13339 16175 13345
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 12584 13280 12940 13308
rect 12989 13311 13047 13317
rect 12584 13268 12590 13280
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13262 13308 13268 13320
rect 13035 13280 13268 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 4157 13243 4215 13249
rect 2556 13212 3648 13240
rect 3712 13212 3924 13240
rect 2556 13200 2562 13212
rect 3712 13172 3740 13212
rect 2332 13144 3740 13172
rect 3896 13172 3924 13212
rect 4157 13209 4169 13243
rect 4203 13240 4215 13243
rect 4522 13240 4528 13252
rect 4203 13212 4528 13240
rect 4203 13209 4215 13212
rect 4157 13203 4215 13209
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 4614 13200 4620 13252
rect 4672 13200 4678 13252
rect 7837 13243 7895 13249
rect 3957 13175 4015 13181
rect 3957 13172 3969 13175
rect 3896 13144 3969 13172
rect 3957 13141 3969 13144
rect 4003 13172 4015 13175
rect 4798 13172 4804 13184
rect 4003 13144 4804 13172
rect 4003 13141 4015 13144
rect 3957 13135 4015 13141
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 5832 13172 5860 13240
rect 7837 13209 7849 13243
rect 7883 13240 7895 13243
rect 9122 13240 9128 13252
rect 7883 13212 9128 13240
rect 7883 13209 7895 13212
rect 7837 13203 7895 13209
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 10134 13200 10140 13252
rect 10192 13240 10198 13252
rect 11517 13243 11575 13249
rect 10192 13212 10350 13240
rect 10192 13200 10198 13212
rect 11517 13209 11529 13243
rect 11563 13209 11575 13243
rect 11517 13203 11575 13209
rect 5500 13144 5860 13172
rect 5500 13132 5506 13144
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 6972 13144 7297 13172
rect 6972 13132 6978 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 7285 13135 7343 13141
rect 7650 13132 7656 13184
rect 7708 13132 7714 13184
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9732 13144 9965 13172
rect 9732 13132 9738 13144
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 9953 13135 10011 13141
rect 10045 13175 10103 13181
rect 10045 13141 10057 13175
rect 10091 13172 10103 13175
rect 11422 13172 11428 13184
rect 10091 13144 11428 13172
rect 10091 13141 10103 13144
rect 10045 13135 10103 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11532 13172 11560 13203
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 12713 13243 12771 13249
rect 12713 13240 12725 13243
rect 11848 13212 12725 13240
rect 11848 13200 11854 13212
rect 12713 13209 12725 13212
rect 12759 13209 12771 13243
rect 12713 13203 12771 13209
rect 12802 13200 12808 13252
rect 12860 13240 12866 13252
rect 13004 13240 13032 13271
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 13541 13311 13599 13317
rect 13541 13308 13553 13311
rect 13412 13280 13553 13308
rect 13412 13268 13418 13280
rect 13541 13277 13553 13280
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 12860 13212 13032 13240
rect 13740 13240 13768 13271
rect 13814 13268 13820 13320
rect 13872 13268 13878 13320
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14056 13280 14933 13308
rect 14056 13268 14062 13280
rect 14921 13277 14933 13280
rect 14967 13308 14979 13311
rect 15102 13308 15108 13320
rect 14967 13280 15108 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 16022 13308 16028 13320
rect 15856 13280 16028 13308
rect 14458 13240 14464 13252
rect 13740 13212 14464 13240
rect 12860 13200 12866 13212
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 15856 13240 15884 13280
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 18509 13311 18567 13317
rect 18509 13308 18521 13311
rect 18472 13280 18521 13308
rect 18472 13268 18478 13280
rect 18509 13277 18521 13280
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 19518 13268 19524 13320
rect 19576 13268 19582 13320
rect 19610 13268 19616 13320
rect 19668 13308 19674 13320
rect 20088 13317 20116 13416
rect 21269 13413 21281 13416
rect 21315 13413 21327 13447
rect 21269 13407 21327 13413
rect 20254 13336 20260 13388
rect 20312 13336 20318 13388
rect 21085 13379 21143 13385
rect 21085 13345 21097 13379
rect 21131 13345 21143 13379
rect 21928 13376 21956 13472
rect 24210 13444 24216 13456
rect 22664 13416 24216 13444
rect 22664 13385 22692 13416
rect 24210 13404 24216 13416
rect 24268 13404 24274 13456
rect 27801 13447 27859 13453
rect 27801 13413 27813 13447
rect 27847 13444 27859 13447
rect 27890 13444 27896 13456
rect 27847 13416 27896 13444
rect 27847 13413 27859 13416
rect 27801 13407 27859 13413
rect 27890 13404 27896 13416
rect 27948 13404 27954 13456
rect 28626 13404 28632 13456
rect 28684 13404 28690 13456
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 21928 13348 22661 13376
rect 21085 13339 21143 13345
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 23934 13376 23940 13388
rect 22649 13339 22707 13345
rect 23216 13348 23940 13376
rect 20073 13311 20131 13317
rect 20073 13308 20085 13311
rect 19668 13280 20085 13308
rect 19668 13268 19674 13280
rect 20073 13277 20085 13280
rect 20119 13277 20131 13311
rect 20073 13271 20131 13277
rect 20162 13268 20168 13320
rect 20220 13308 20226 13320
rect 21100 13308 21128 13339
rect 20220 13280 21128 13308
rect 21361 13311 21419 13317
rect 20220 13268 20226 13280
rect 21361 13277 21373 13311
rect 21407 13308 21419 13311
rect 21542 13308 21548 13320
rect 21407 13280 21548 13308
rect 21407 13277 21419 13280
rect 21361 13271 21419 13277
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13308 22615 13311
rect 23216 13308 23244 13348
rect 23934 13336 23940 13348
rect 23992 13336 23998 13388
rect 24946 13376 24952 13388
rect 24596 13348 24952 13376
rect 22603 13280 23244 13308
rect 23293 13311 23351 13317
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 23293 13277 23305 13311
rect 23339 13308 23351 13311
rect 23382 13308 23388 13320
rect 23339 13280 23388 13308
rect 23339 13277 23351 13280
rect 23293 13271 23351 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13308 23627 13311
rect 23658 13308 23664 13320
rect 23615 13280 23664 13308
rect 23615 13277 23627 13280
rect 23569 13271 23627 13277
rect 17678 13240 17684 13252
rect 14752 13212 15884 13240
rect 17158 13212 17684 13240
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11532 13144 11897 13172
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 12434 13172 12440 13184
rect 12391 13144 12440 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 12434 13132 12440 13144
rect 12492 13172 12498 13184
rect 12986 13172 12992 13184
rect 12492 13144 12992 13172
rect 12492 13132 12498 13144
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 14752 13172 14780 13212
rect 17678 13200 17684 13212
rect 17736 13240 17742 13252
rect 18138 13240 18144 13252
rect 17736 13212 18144 13240
rect 17736 13200 17742 13212
rect 18138 13200 18144 13212
rect 18196 13200 18202 13252
rect 20901 13243 20959 13249
rect 20901 13209 20913 13243
rect 20947 13240 20959 13243
rect 21174 13240 21180 13252
rect 20947 13212 21180 13240
rect 20947 13209 20959 13212
rect 20901 13203 20959 13209
rect 21174 13200 21180 13212
rect 21232 13240 21238 13252
rect 21634 13240 21640 13252
rect 21232 13212 21640 13240
rect 21232 13200 21238 13212
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 22465 13243 22523 13249
rect 22465 13209 22477 13243
rect 22511 13240 22523 13243
rect 23584 13240 23612 13271
rect 23658 13268 23664 13280
rect 23716 13308 23722 13320
rect 23845 13311 23903 13317
rect 23845 13308 23857 13311
rect 23716 13280 23857 13308
rect 23716 13268 23722 13280
rect 23845 13277 23857 13280
rect 23891 13308 23903 13311
rect 24210 13308 24216 13320
rect 23891 13280 24216 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 24596 13317 24624 13348
rect 24946 13336 24952 13348
rect 25004 13376 25010 13388
rect 25593 13379 25651 13385
rect 25593 13376 25605 13379
rect 25004 13348 25605 13376
rect 25004 13336 25010 13348
rect 25593 13345 25605 13348
rect 25639 13345 25651 13379
rect 25593 13339 25651 13345
rect 28166 13336 28172 13388
rect 28224 13376 28230 13388
rect 28353 13379 28411 13385
rect 28353 13376 28365 13379
rect 28224 13348 28365 13376
rect 28224 13336 28230 13348
rect 28353 13345 28365 13348
rect 28399 13345 28411 13379
rect 28353 13339 28411 13345
rect 28445 13379 28503 13385
rect 28445 13345 28457 13379
rect 28491 13376 28503 13379
rect 28644 13376 28672 13404
rect 28491 13348 28672 13376
rect 28491 13345 28503 13348
rect 28445 13339 28503 13345
rect 30374 13336 30380 13388
rect 30432 13376 30438 13388
rect 30561 13379 30619 13385
rect 30561 13376 30573 13379
rect 30432 13348 30573 13376
rect 30432 13336 30438 13348
rect 30561 13345 30573 13348
rect 30607 13345 30619 13379
rect 30561 13339 30619 13345
rect 32493 13379 32551 13385
rect 32493 13345 32505 13379
rect 32539 13376 32551 13379
rect 32766 13376 32772 13388
rect 32539 13348 32772 13376
rect 32539 13345 32551 13348
rect 32493 13339 32551 13345
rect 32766 13336 32772 13348
rect 32824 13376 32830 13388
rect 34701 13379 34759 13385
rect 34701 13376 34713 13379
rect 32824 13348 34713 13376
rect 32824 13336 32830 13348
rect 34701 13345 34713 13348
rect 34747 13376 34759 13379
rect 35986 13376 35992 13388
rect 34747 13348 35992 13376
rect 34747 13345 34759 13348
rect 34701 13339 34759 13345
rect 35986 13336 35992 13348
rect 36044 13336 36050 13388
rect 36722 13336 36728 13388
rect 36780 13336 36786 13388
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 24854 13268 24860 13320
rect 24912 13268 24918 13320
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 22511 13212 23612 13240
rect 22511 13209 22523 13212
rect 22465 13203 22523 13209
rect 23750 13200 23756 13252
rect 23808 13240 23814 13252
rect 24397 13243 24455 13249
rect 24397 13240 24409 13243
rect 23808 13212 24409 13240
rect 23808 13200 23814 13212
rect 24397 13209 24409 13212
rect 24443 13209 24455 13243
rect 24397 13203 24455 13209
rect 25056 13240 25084 13271
rect 25130 13268 25136 13320
rect 25188 13268 25194 13320
rect 25409 13311 25467 13317
rect 25409 13277 25421 13311
rect 25455 13277 25467 13311
rect 25409 13271 25467 13277
rect 25424 13240 25452 13271
rect 26510 13268 26516 13320
rect 26568 13268 26574 13320
rect 26602 13268 26608 13320
rect 26660 13308 26666 13320
rect 26789 13311 26847 13317
rect 26789 13308 26801 13311
rect 26660 13280 26801 13308
rect 26660 13268 26666 13280
rect 26789 13277 26801 13280
rect 26835 13308 26847 13311
rect 28537 13311 28595 13317
rect 26835 13280 27752 13308
rect 26835 13277 26847 13280
rect 26789 13271 26847 13277
rect 25056 13212 25452 13240
rect 13219 13144 14780 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 14826 13132 14832 13184
rect 14884 13132 14890 13184
rect 18690 13132 18696 13184
rect 18748 13132 18754 13184
rect 19886 13132 19892 13184
rect 19944 13132 19950 13184
rect 21082 13132 21088 13184
rect 21140 13132 21146 13184
rect 23106 13132 23112 13184
rect 23164 13132 23170 13184
rect 24213 13175 24271 13181
rect 24213 13141 24225 13175
rect 24259 13172 24271 13175
rect 25056 13172 25084 13212
rect 26694 13200 26700 13252
rect 26752 13200 26758 13252
rect 27614 13200 27620 13252
rect 27672 13200 27678 13252
rect 27724 13240 27752 13280
rect 28537 13277 28549 13311
rect 28583 13277 28595 13311
rect 28537 13271 28595 13277
rect 28552 13240 28580 13271
rect 28626 13268 28632 13320
rect 28684 13268 28690 13320
rect 34330 13308 34336 13320
rect 33902 13280 34336 13308
rect 34330 13268 34336 13280
rect 34388 13268 34394 13320
rect 28718 13240 28724 13252
rect 27724 13212 28724 13240
rect 28718 13200 28724 13212
rect 28776 13200 28782 13252
rect 29086 13200 29092 13252
rect 29144 13240 29150 13252
rect 29641 13243 29699 13249
rect 29641 13240 29653 13243
rect 29144 13212 29653 13240
rect 29144 13200 29150 13212
rect 29641 13209 29653 13212
rect 29687 13240 29699 13243
rect 29917 13243 29975 13249
rect 29917 13240 29929 13243
rect 29687 13212 29929 13240
rect 29687 13209 29699 13212
rect 29641 13203 29699 13209
rect 29917 13209 29929 13212
rect 29963 13209 29975 13243
rect 29917 13203 29975 13209
rect 30837 13243 30895 13249
rect 30837 13209 30849 13243
rect 30883 13240 30895 13243
rect 31110 13240 31116 13252
rect 30883 13212 31116 13240
rect 30883 13209 30895 13212
rect 30837 13203 30895 13209
rect 31110 13200 31116 13212
rect 31168 13200 31174 13252
rect 31294 13200 31300 13252
rect 31352 13200 31358 13252
rect 32769 13243 32827 13249
rect 32769 13209 32781 13243
rect 32815 13240 32827 13243
rect 32858 13240 32864 13252
rect 32815 13212 32864 13240
rect 32815 13209 32827 13212
rect 32769 13203 32827 13209
rect 32858 13200 32864 13212
rect 32916 13200 32922 13252
rect 34517 13243 34575 13249
rect 34517 13240 34529 13243
rect 34072 13212 34529 13240
rect 24259 13144 25084 13172
rect 26789 13175 26847 13181
rect 24259 13141 24271 13144
rect 24213 13135 24271 13141
rect 26789 13141 26801 13175
rect 26835 13172 26847 13175
rect 26878 13172 26884 13184
rect 26835 13144 26884 13172
rect 26835 13141 26847 13144
rect 26789 13135 26847 13141
rect 26878 13132 26884 13144
rect 26936 13132 26942 13184
rect 28169 13175 28227 13181
rect 28169 13141 28181 13175
rect 28215 13172 28227 13175
rect 28258 13172 28264 13184
rect 28215 13144 28264 13172
rect 28215 13141 28227 13144
rect 28169 13135 28227 13141
rect 28258 13132 28264 13144
rect 28316 13132 28322 13184
rect 29730 13132 29736 13184
rect 29788 13132 29794 13184
rect 31202 13132 31208 13184
rect 31260 13172 31266 13184
rect 32309 13175 32367 13181
rect 32309 13172 32321 13175
rect 31260 13144 32321 13172
rect 31260 13132 31266 13144
rect 32309 13141 32321 13144
rect 32355 13141 32367 13175
rect 32309 13135 32367 13141
rect 33502 13132 33508 13184
rect 33560 13172 33566 13184
rect 34072 13172 34100 13212
rect 34517 13209 34529 13212
rect 34563 13209 34575 13243
rect 34517 13203 34575 13209
rect 34698 13200 34704 13252
rect 34756 13240 34762 13252
rect 34977 13243 35035 13249
rect 34977 13240 34989 13243
rect 34756 13212 34989 13240
rect 34756 13200 34762 13212
rect 34977 13209 34989 13212
rect 35023 13209 35035 13243
rect 36202 13212 36308 13240
rect 34977 13203 35035 13209
rect 33560 13144 34100 13172
rect 36280 13172 36308 13212
rect 36998 13200 37004 13252
rect 37056 13200 37062 13252
rect 37458 13240 37464 13252
rect 37108 13212 37464 13240
rect 37108 13172 37136 13212
rect 37458 13200 37464 13212
rect 37516 13200 37522 13252
rect 36280 13144 37136 13172
rect 38473 13175 38531 13181
rect 33560 13132 33566 13144
rect 38473 13141 38485 13175
rect 38519 13172 38531 13175
rect 38519 13144 38884 13172
rect 38519 13141 38531 13144
rect 38473 13135 38531 13141
rect 1104 13082 38824 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 38824 13082
rect 1104 13008 38824 13030
rect 4249 12971 4307 12977
rect 4249 12937 4261 12971
rect 4295 12968 4307 12971
rect 4522 12968 4528 12980
rect 4295 12940 4528 12968
rect 4295 12937 4307 12940
rect 4249 12931 4307 12937
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4672 12940 4813 12968
rect 4672 12928 4678 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 4801 12931 4859 12937
rect 4982 12928 4988 12980
rect 5040 12968 5046 12980
rect 5534 12968 5540 12980
rect 5040 12940 5540 12968
rect 5040 12928 5046 12940
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 11149 12971 11207 12977
rect 11149 12968 11161 12971
rect 9640 12940 11161 12968
rect 9640 12928 9646 12940
rect 11149 12937 11161 12940
rect 11195 12937 11207 12971
rect 11149 12931 11207 12937
rect 12161 12971 12219 12977
rect 12161 12937 12173 12971
rect 12207 12968 12219 12971
rect 12526 12968 12532 12980
rect 12207 12940 12532 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 2774 12860 2780 12912
rect 2832 12860 2838 12912
rect 4154 12900 4160 12912
rect 4002 12872 4160 12900
rect 4154 12860 4160 12872
rect 4212 12900 4218 12912
rect 5442 12900 5448 12912
rect 4212 12872 5448 12900
rect 4212 12860 4218 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 6914 12860 6920 12912
rect 6972 12860 6978 12912
rect 7466 12860 7472 12912
rect 7524 12860 7530 12912
rect 9674 12860 9680 12912
rect 9732 12860 9738 12912
rect 10134 12860 10140 12912
rect 10192 12860 10198 12912
rect 11164 12900 11192 12931
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 12621 12971 12679 12977
rect 12621 12937 12633 12971
rect 12667 12968 12679 12971
rect 12894 12968 12900 12980
rect 12667 12940 12900 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 18785 12971 18843 12977
rect 18785 12937 18797 12971
rect 18831 12968 18843 12971
rect 19150 12968 19156 12980
rect 18831 12940 19156 12968
rect 18831 12937 18843 12940
rect 18785 12931 18843 12937
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 21542 12928 21548 12980
rect 21600 12928 21606 12980
rect 21634 12928 21640 12980
rect 21692 12968 21698 12980
rect 27614 12968 27620 12980
rect 21692 12940 27620 12968
rect 21692 12928 21698 12940
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 28626 12928 28632 12980
rect 28684 12968 28690 12980
rect 28810 12968 28816 12980
rect 28684 12940 28816 12968
rect 28684 12928 28690 12940
rect 28810 12928 28816 12940
rect 28868 12928 28874 12980
rect 30650 12928 30656 12980
rect 30708 12928 30714 12980
rect 31110 12928 31116 12980
rect 31168 12928 31174 12980
rect 31294 12928 31300 12980
rect 31352 12968 31358 12980
rect 33410 12968 33416 12980
rect 31352 12940 33416 12968
rect 31352 12928 31358 12940
rect 33410 12928 33416 12940
rect 33468 12928 33474 12980
rect 35434 12928 35440 12980
rect 35492 12968 35498 12980
rect 35713 12971 35771 12977
rect 35713 12968 35725 12971
rect 35492 12940 35725 12968
rect 35492 12928 35498 12940
rect 35713 12937 35725 12940
rect 35759 12937 35771 12971
rect 35713 12931 35771 12937
rect 36354 12928 36360 12980
rect 36412 12968 36418 12980
rect 36449 12971 36507 12977
rect 36449 12968 36461 12971
rect 36412 12940 36461 12968
rect 36412 12928 36418 12940
rect 36449 12937 36461 12940
rect 36495 12937 36507 12971
rect 36449 12931 36507 12937
rect 12434 12900 12440 12912
rect 11164 12872 12440 12900
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 14918 12860 14924 12912
rect 14976 12860 14982 12912
rect 15746 12860 15752 12912
rect 15804 12900 15810 12912
rect 17313 12903 17371 12909
rect 15804 12872 15976 12900
rect 15804 12860 15810 12872
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12832 4583 12835
rect 4614 12832 4620 12844
rect 4571 12804 4620 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12832 4767 12835
rect 4798 12832 4804 12844
rect 4755 12804 4804 12832
rect 4755 12801 4767 12804
rect 4709 12795 4767 12801
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12832 4951 12835
rect 5258 12832 5264 12844
rect 4939 12804 5264 12832
rect 4939 12801 4951 12804
rect 4893 12795 4951 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 6178 12832 6184 12844
rect 5960 12804 6184 12832
rect 5960 12792 5966 12804
rect 6178 12792 6184 12804
rect 6236 12832 6242 12844
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 6236 12804 6653 12832
rect 6236 12792 6242 12804
rect 6641 12801 6653 12804
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8352 12804 9413 12832
rect 8352 12792 8358 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 11422 12792 11428 12844
rect 11480 12832 11486 12844
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11480 12804 11529 12832
rect 11480 12792 11486 12804
rect 11517 12801 11529 12804
rect 11563 12832 11575 12835
rect 12802 12832 12808 12844
rect 11563 12804 12808 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 13078 12792 13084 12844
rect 13136 12792 13142 12844
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 13538 12832 13544 12844
rect 13311 12804 13544 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 15948 12841 15976 12872
rect 17313 12869 17325 12903
rect 17359 12900 17371 12903
rect 17402 12900 17408 12912
rect 17359 12872 17408 12900
rect 17359 12869 17371 12872
rect 17313 12863 17371 12869
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 18046 12860 18052 12912
rect 18104 12860 18110 12912
rect 24946 12900 24952 12912
rect 24044 12872 24952 12900
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16574 12832 16580 12844
rect 15979 12804 16580 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16574 12792 16580 12804
rect 16632 12832 16638 12844
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16632 12804 17049 12832
rect 16632 12792 16638 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 19484 12804 19533 12832
rect 19484 12792 19490 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12832 19763 12835
rect 19886 12832 19892 12844
rect 19751 12804 19892 12832
rect 19751 12801 19763 12804
rect 19705 12795 19763 12801
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12832 20131 12835
rect 21082 12832 21088 12844
rect 20119 12804 21088 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 23753 12835 23811 12841
rect 23753 12801 23765 12835
rect 23799 12832 23811 12835
rect 23842 12832 23848 12844
rect 23799 12804 23848 12832
rect 23799 12801 23811 12804
rect 23753 12795 23811 12801
rect 23842 12792 23848 12804
rect 23900 12792 23906 12844
rect 24044 12841 24072 12872
rect 24946 12860 24952 12872
rect 25004 12860 25010 12912
rect 26418 12860 26424 12912
rect 26476 12900 26482 12912
rect 26694 12900 26700 12912
rect 26476 12872 26700 12900
rect 26476 12860 26482 12872
rect 26694 12860 26700 12872
rect 26752 12900 26758 12912
rect 27522 12900 27528 12912
rect 26752 12872 27528 12900
rect 26752 12860 26758 12872
rect 27522 12860 27528 12872
rect 27580 12860 27586 12912
rect 27890 12860 27896 12912
rect 27948 12860 27954 12912
rect 29822 12860 29828 12912
rect 29880 12860 29886 12912
rect 30374 12860 30380 12912
rect 30432 12900 30438 12912
rect 30668 12900 30696 12928
rect 33045 12903 33103 12909
rect 30432 12872 30604 12900
rect 30668 12872 31524 12900
rect 30432 12860 30438 12872
rect 24029 12835 24087 12841
rect 24029 12801 24041 12835
rect 24075 12801 24087 12835
rect 24029 12795 24087 12801
rect 24210 12792 24216 12844
rect 24268 12792 24274 12844
rect 24670 12792 24676 12844
rect 24728 12832 24734 12844
rect 25130 12832 25136 12844
rect 24728 12804 25136 12832
rect 24728 12792 24734 12804
rect 25130 12792 25136 12804
rect 25188 12792 25194 12844
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12832 26387 12835
rect 26510 12832 26516 12844
rect 26375 12804 26516 12832
rect 26375 12801 26387 12804
rect 26329 12795 26387 12801
rect 26510 12792 26516 12804
rect 26568 12792 26574 12844
rect 26602 12792 26608 12844
rect 26660 12792 26666 12844
rect 30576 12841 30604 12872
rect 31496 12844 31524 12872
rect 33045 12869 33057 12903
rect 33091 12900 33103 12903
rect 33226 12900 33232 12912
rect 33091 12872 33232 12900
rect 33091 12869 33103 12872
rect 33045 12863 33103 12869
rect 33226 12860 33232 12872
rect 33284 12860 33290 12912
rect 36464 12900 36492 12931
rect 36998 12928 37004 12980
rect 37056 12928 37062 12980
rect 37277 12903 37335 12909
rect 37277 12900 37289 12903
rect 36004 12872 36308 12900
rect 36464 12872 36952 12900
rect 30561 12835 30619 12841
rect 30561 12801 30573 12835
rect 30607 12801 30619 12835
rect 30561 12795 30619 12801
rect 30837 12835 30895 12841
rect 30837 12801 30849 12835
rect 30883 12801 30895 12835
rect 30837 12795 30895 12801
rect 2498 12724 2504 12776
rect 2556 12724 2562 12776
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4982 12764 4988 12776
rect 4387 12736 4988 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4816 12708 4844 12736
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 9214 12724 9220 12776
rect 9272 12724 9278 12776
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 14148 12736 14197 12764
rect 14148 12724 14154 12736
rect 14185 12733 14197 12736
rect 14231 12733 14243 12767
rect 14185 12727 14243 12733
rect 15654 12724 15660 12776
rect 15712 12724 15718 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20165 12767 20223 12773
rect 20165 12764 20177 12767
rect 19843 12736 20177 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 20165 12733 20177 12736
rect 20211 12733 20223 12767
rect 20165 12727 20223 12733
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20496 12736 20729 12764
rect 20496 12724 20502 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 20901 12767 20959 12773
rect 20901 12733 20913 12767
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 4798 12656 4804 12708
rect 4856 12656 4862 12708
rect 8389 12699 8447 12705
rect 8389 12665 8401 12699
rect 8435 12696 8447 12699
rect 8478 12696 8484 12708
rect 8435 12668 8484 12696
rect 8435 12665 8447 12668
rect 8389 12659 8447 12665
rect 8478 12656 8484 12668
rect 8536 12696 8542 12708
rect 8536 12668 8800 12696
rect 8536 12656 8542 12668
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 8018 12628 8024 12640
rect 7524 12600 8024 12628
rect 7524 12588 7530 12600
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 8628 12600 8677 12628
rect 8628 12588 8634 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 8772 12628 8800 12668
rect 19610 12656 19616 12708
rect 19668 12696 19674 12708
rect 20073 12699 20131 12705
rect 20073 12696 20085 12699
rect 19668 12668 20085 12696
rect 19668 12656 19674 12668
rect 20073 12665 20085 12668
rect 20119 12665 20131 12699
rect 20073 12659 20131 12665
rect 20254 12656 20260 12708
rect 20312 12696 20318 12708
rect 20806 12696 20812 12708
rect 20312 12668 20812 12696
rect 20312 12656 20318 12668
rect 20806 12656 20812 12668
rect 20864 12696 20870 12708
rect 20916 12696 20944 12727
rect 26234 12724 26240 12776
rect 26292 12764 26298 12776
rect 26973 12767 27031 12773
rect 26973 12764 26985 12767
rect 26292 12736 26985 12764
rect 26292 12724 26298 12736
rect 26973 12733 26985 12736
rect 27019 12733 27031 12767
rect 26973 12727 27031 12733
rect 27246 12724 27252 12776
rect 27304 12724 27310 12776
rect 28534 12724 28540 12776
rect 28592 12764 28598 12776
rect 30285 12767 30343 12773
rect 30285 12764 30297 12767
rect 28592 12736 30297 12764
rect 28592 12724 28598 12736
rect 30285 12733 30297 12736
rect 30331 12733 30343 12767
rect 30285 12727 30343 12733
rect 20864 12668 20944 12696
rect 20864 12656 20870 12668
rect 10134 12628 10140 12640
rect 8772 12600 10140 12628
rect 8665 12591 8723 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 13446 12588 13452 12640
rect 13504 12588 13510 12640
rect 19334 12588 19340 12640
rect 19392 12588 19398 12640
rect 23474 12588 23480 12640
rect 23532 12628 23538 12640
rect 23569 12631 23627 12637
rect 23569 12628 23581 12631
rect 23532 12600 23581 12628
rect 23532 12588 23538 12600
rect 23569 12597 23581 12600
rect 23615 12597 23627 12631
rect 23569 12591 23627 12597
rect 26786 12588 26792 12640
rect 26844 12588 26850 12640
rect 28718 12588 28724 12640
rect 28776 12588 28782 12640
rect 30190 12588 30196 12640
rect 30248 12628 30254 12640
rect 30852 12628 30880 12795
rect 31110 12792 31116 12844
rect 31168 12832 31174 12844
rect 31389 12835 31447 12841
rect 31389 12832 31401 12835
rect 31168 12804 31401 12832
rect 31168 12792 31174 12804
rect 31389 12801 31401 12804
rect 31435 12801 31447 12835
rect 31389 12795 31447 12801
rect 31478 12792 31484 12844
rect 31536 12792 31542 12844
rect 31570 12792 31576 12844
rect 31628 12792 31634 12844
rect 31754 12792 31760 12844
rect 31812 12792 31818 12844
rect 36004 12841 36032 12872
rect 35989 12835 36047 12841
rect 35989 12801 36001 12835
rect 36035 12801 36047 12835
rect 35989 12795 36047 12801
rect 36078 12792 36084 12844
rect 36136 12792 36142 12844
rect 36170 12792 36176 12844
rect 36228 12792 36234 12844
rect 36280 12832 36308 12872
rect 36280 12804 36584 12832
rect 31021 12767 31079 12773
rect 31021 12733 31033 12767
rect 31067 12764 31079 12767
rect 31202 12764 31208 12776
rect 31067 12736 31208 12764
rect 31067 12733 31079 12736
rect 31021 12727 31079 12733
rect 31202 12724 31208 12736
rect 31260 12724 31266 12776
rect 35897 12767 35955 12773
rect 35897 12733 35909 12767
rect 35943 12733 35955 12767
rect 36096 12764 36124 12792
rect 36262 12764 36268 12776
rect 36096 12736 36268 12764
rect 35897 12727 35955 12733
rect 32674 12656 32680 12708
rect 32732 12656 32738 12708
rect 34606 12696 34612 12708
rect 33060 12668 34612 12696
rect 31294 12628 31300 12640
rect 30248 12600 31300 12628
rect 30248 12588 30254 12600
rect 31294 12588 31300 12600
rect 31352 12588 31358 12640
rect 33060 12637 33088 12668
rect 34606 12656 34612 12668
rect 34664 12656 34670 12708
rect 35912 12696 35940 12727
rect 36262 12724 36268 12736
rect 36320 12724 36326 12776
rect 36556 12756 36584 12804
rect 36630 12792 36636 12844
rect 36688 12792 36694 12844
rect 36924 12841 36952 12872
rect 37108 12872 37289 12900
rect 37108 12841 37136 12872
rect 37277 12869 37289 12872
rect 37323 12869 37335 12903
rect 37277 12863 37335 12869
rect 36909 12835 36967 12841
rect 36909 12801 36921 12835
rect 36955 12801 36967 12835
rect 36909 12795 36967 12801
rect 37093 12835 37151 12841
rect 37093 12801 37105 12835
rect 37139 12801 37151 12835
rect 37553 12835 37611 12841
rect 37553 12832 37565 12835
rect 37093 12795 37151 12801
rect 37200 12804 37565 12832
rect 36817 12767 36875 12773
rect 36817 12764 36829 12767
rect 36740 12756 36829 12764
rect 36556 12736 36829 12756
rect 36556 12728 36768 12736
rect 36817 12733 36829 12736
rect 36863 12764 36875 12767
rect 36998 12764 37004 12776
rect 36863 12736 37004 12764
rect 36863 12733 36875 12736
rect 36817 12727 36875 12733
rect 36998 12724 37004 12736
rect 37056 12764 37062 12776
rect 37200 12764 37228 12804
rect 37553 12801 37565 12804
rect 37599 12832 37611 12835
rect 38856 12832 38884 13144
rect 37599 12804 38884 12832
rect 37599 12801 37611 12804
rect 37553 12795 37611 12801
rect 37056 12736 37228 12764
rect 37056 12724 37062 12736
rect 37274 12724 37280 12776
rect 37332 12724 37338 12776
rect 35912 12668 36676 12696
rect 36648 12640 36676 12668
rect 33045 12631 33103 12637
rect 33045 12597 33057 12631
rect 33091 12597 33103 12631
rect 33045 12591 33103 12597
rect 33134 12588 33140 12640
rect 33192 12628 33198 12640
rect 33229 12631 33287 12637
rect 33229 12628 33241 12631
rect 33192 12600 33241 12628
rect 33192 12588 33198 12600
rect 33229 12597 33241 12600
rect 33275 12597 33287 12631
rect 33229 12591 33287 12597
rect 36630 12588 36636 12640
rect 36688 12628 36694 12640
rect 37461 12631 37519 12637
rect 37461 12628 37473 12631
rect 36688 12600 37473 12628
rect 36688 12588 36694 12600
rect 37461 12597 37473 12600
rect 37507 12628 37519 12631
rect 37826 12628 37832 12640
rect 37507 12600 37832 12628
rect 37507 12597 37519 12600
rect 37461 12591 37519 12597
rect 37826 12588 37832 12600
rect 37884 12588 37890 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 4801 12427 4859 12433
rect 4801 12393 4813 12427
rect 4847 12424 4859 12427
rect 5166 12424 5172 12436
rect 4847 12396 5172 12424
rect 4847 12393 4859 12396
rect 4801 12387 4859 12393
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 4816 12356 4844 12387
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 9180 12396 9229 12424
rect 9180 12384 9186 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 10134 12384 10140 12436
rect 10192 12384 10198 12436
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 13173 12427 13231 12433
rect 13173 12424 13185 12427
rect 13136 12396 13185 12424
rect 13136 12384 13142 12396
rect 13173 12393 13185 12396
rect 13219 12393 13231 12427
rect 13173 12387 13231 12393
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13412 12396 14105 12424
rect 13412 12384 13418 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 15286 12424 15292 12436
rect 14599 12396 15292 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15381 12427 15439 12433
rect 15381 12393 15393 12427
rect 15427 12424 15439 12427
rect 15654 12424 15660 12436
rect 15427 12396 15660 12424
rect 15427 12393 15439 12396
rect 15381 12387 15439 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 17126 12424 17132 12436
rect 16224 12396 17132 12424
rect 4764 12328 4844 12356
rect 4764 12316 4770 12328
rect 5810 12316 5816 12368
rect 5868 12316 5874 12368
rect 10870 12356 10876 12368
rect 7576 12328 10876 12356
rect 4798 12288 4804 12300
rect 4356 12260 4804 12288
rect 4356 12232 4384 12260
rect 4798 12248 4804 12260
rect 4856 12288 4862 12300
rect 7576 12288 7604 12328
rect 10870 12316 10876 12328
rect 10928 12356 10934 12368
rect 11238 12356 11244 12368
rect 10928 12328 11244 12356
rect 10928 12316 10934 12328
rect 11238 12316 11244 12328
rect 11296 12316 11302 12368
rect 13446 12356 13452 12368
rect 12636 12328 13452 12356
rect 4856 12260 7604 12288
rect 4856 12248 4862 12260
rect 7650 12248 7656 12300
rect 7708 12288 7714 12300
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7708 12260 7941 12288
rect 7708 12248 7714 12260
rect 7929 12257 7941 12260
rect 7975 12288 7987 12291
rect 8110 12288 8116 12300
rect 7975 12260 8116 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8110 12248 8116 12260
rect 8168 12288 8174 12300
rect 12636 12297 12664 12328
rect 13446 12316 13452 12328
rect 13504 12356 13510 12368
rect 16224 12356 16252 12396
rect 17126 12384 17132 12396
rect 17184 12384 17190 12436
rect 20806 12384 20812 12436
rect 20864 12424 20870 12436
rect 21085 12427 21143 12433
rect 21085 12424 21097 12427
rect 20864 12396 21097 12424
rect 20864 12384 20870 12396
rect 21085 12393 21097 12396
rect 21131 12393 21143 12427
rect 21085 12387 21143 12393
rect 24857 12427 24915 12433
rect 24857 12393 24869 12427
rect 24903 12424 24915 12427
rect 25130 12424 25136 12436
rect 24903 12396 25136 12424
rect 24903 12393 24915 12396
rect 24857 12387 24915 12393
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 26789 12427 26847 12433
rect 26789 12393 26801 12427
rect 26835 12424 26847 12427
rect 26878 12424 26884 12436
rect 26835 12396 26884 12424
rect 26835 12393 26847 12396
rect 26789 12387 26847 12393
rect 26878 12384 26884 12396
rect 26936 12384 26942 12436
rect 26973 12427 27031 12433
rect 26973 12393 26985 12427
rect 27019 12424 27031 12427
rect 27246 12424 27252 12436
rect 27019 12396 27252 12424
rect 27019 12393 27031 12396
rect 26973 12387 27031 12393
rect 27246 12384 27252 12396
rect 27304 12384 27310 12436
rect 28258 12384 28264 12436
rect 28316 12424 28322 12436
rect 28353 12427 28411 12433
rect 28353 12424 28365 12427
rect 28316 12396 28365 12424
rect 28316 12384 28322 12396
rect 28353 12393 28365 12396
rect 28399 12393 28411 12427
rect 29365 12427 29423 12433
rect 29365 12424 29377 12427
rect 28353 12387 28411 12393
rect 28644 12396 29377 12424
rect 23017 12359 23075 12365
rect 23017 12356 23029 12359
rect 13504 12328 14964 12356
rect 13504 12316 13510 12328
rect 12529 12291 12587 12297
rect 8168 12260 10364 12288
rect 8168 12248 8174 12260
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 4338 12220 4344 12232
rect 3651 12192 4344 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 5077 12223 5135 12229
rect 5077 12220 5089 12223
rect 4816 12192 5089 12220
rect 3418 12112 3424 12164
rect 3476 12152 3482 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 3476 12124 4169 12152
rect 3476 12112 3482 12124
rect 4157 12121 4169 12124
rect 4203 12121 4215 12155
rect 4157 12115 4215 12121
rect 4430 12112 4436 12164
rect 4488 12152 4494 12164
rect 4816 12161 4844 12192
rect 5077 12189 5089 12192
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 5224 12192 6101 12220
rect 5224 12180 5230 12192
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 6178 12180 6184 12232
rect 6236 12180 6242 12232
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 7800 12192 8156 12220
rect 7800 12180 7806 12192
rect 4785 12155 4844 12161
rect 4785 12152 4797 12155
rect 4488 12124 4797 12152
rect 4488 12112 4494 12124
rect 4785 12121 4797 12124
rect 4831 12124 4844 12155
rect 4985 12155 5043 12161
rect 4831 12121 4843 12124
rect 4785 12115 4843 12121
rect 4985 12121 4997 12155
rect 5031 12121 5043 12155
rect 4985 12115 5043 12121
rect 5721 12155 5779 12161
rect 5721 12121 5733 12155
rect 5767 12152 5779 12155
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 5767 12124 5825 12152
rect 5767 12121 5779 12124
rect 5721 12115 5779 12121
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4522 12084 4528 12096
rect 4387 12056 4528 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 5000 12084 5028 12115
rect 6454 12112 6460 12164
rect 6512 12112 6518 12164
rect 8128 12161 8156 12192
rect 8570 12180 8576 12232
rect 8628 12180 8634 12232
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 8113 12155 8171 12161
rect 7682 12124 8064 12152
rect 5350 12084 5356 12096
rect 5000 12056 5356 12084
rect 5350 12044 5356 12056
rect 5408 12084 5414 12096
rect 5997 12087 6055 12093
rect 5997 12084 6009 12087
rect 5408 12056 6009 12084
rect 5408 12044 5414 12056
rect 5997 12053 6009 12056
rect 6043 12053 6055 12087
rect 8036 12084 8064 12124
rect 8113 12121 8125 12155
rect 8159 12121 8171 12155
rect 8113 12115 8171 12121
rect 8202 12084 8208 12096
rect 8036 12056 8208 12084
rect 5997 12047 6055 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8386 12044 8392 12096
rect 8444 12084 8450 12096
rect 8665 12087 8723 12093
rect 8665 12084 8677 12087
rect 8444 12056 8677 12084
rect 8444 12044 8450 12056
rect 8665 12053 8677 12056
rect 8711 12053 8723 12087
rect 8772 12084 8800 12183
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 9784 12152 9812 12180
rect 10336 12161 10364 12260
rect 12529 12257 12541 12291
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12257 12679 12291
rect 12621 12251 12679 12257
rect 12544 12220 12572 12251
rect 12802 12248 12808 12300
rect 12860 12288 12866 12300
rect 13722 12288 13728 12300
rect 12860 12260 13728 12288
rect 12860 12248 12866 12260
rect 13722 12248 13728 12260
rect 13780 12288 13786 12300
rect 14936 12297 14964 12328
rect 15304 12328 16252 12356
rect 22296 12328 23029 12356
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 13780 12260 14197 12288
rect 13780 12248 13786 12260
rect 13170 12220 13176 12232
rect 12544 12192 13176 12220
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 10105 12155 10163 12161
rect 10105 12152 10117 12155
rect 9784 12124 10117 12152
rect 10105 12121 10117 12124
rect 10151 12121 10163 12155
rect 10105 12115 10163 12121
rect 10321 12155 10379 12161
rect 10321 12121 10333 12155
rect 10367 12121 10379 12155
rect 10321 12115 10379 12121
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12121 11851 12155
rect 13372 12152 13400 12183
rect 13630 12180 13636 12232
rect 13688 12180 13694 12232
rect 13832 12229 13860 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 14829 12291 14887 12297
rect 14829 12257 14841 12291
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 13817 12223 13875 12229
rect 13817 12189 13829 12223
rect 13863 12189 13875 12223
rect 13817 12183 13875 12189
rect 14090 12180 14096 12232
rect 14148 12180 14154 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12189 14427 12223
rect 14844 12222 14872 12251
rect 15304 12232 15332 12328
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 18233 12291 18291 12297
rect 15795 12260 18000 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 14844 12220 15148 12222
rect 15286 12220 15292 12232
rect 14844 12194 15292 12220
rect 15120 12192 15292 12194
rect 14369 12183 14427 12189
rect 13906 12152 13912 12164
rect 13372 12124 13912 12152
rect 11793 12115 11851 12121
rect 8846 12084 8852 12096
rect 8772 12056 8852 12084
rect 8665 12047 8723 12053
rect 8846 12044 8852 12056
rect 8904 12084 8910 12096
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 8904 12056 9965 12084
rect 8904 12044 8910 12056
rect 9953 12053 9965 12056
rect 9999 12053 10011 12087
rect 9953 12047 10011 12053
rect 11606 12044 11612 12096
rect 11664 12084 11670 12096
rect 11808 12084 11836 12115
rect 13906 12112 13912 12124
rect 13964 12152 13970 12164
rect 14108 12152 14136 12180
rect 13964 12124 14136 12152
rect 13964 12112 13970 12124
rect 11664 12056 11836 12084
rect 11664 12044 11670 12056
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 12250 12084 12256 12096
rect 11940 12056 12256 12084
rect 11940 12044 11946 12056
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12713 12087 12771 12093
rect 12713 12053 12725 12087
rect 12759 12084 12771 12087
rect 12802 12084 12808 12096
rect 12759 12056 12808 12084
rect 12759 12053 12771 12056
rect 12713 12047 12771 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13078 12044 13084 12096
rect 13136 12044 13142 12096
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 13722 12084 13728 12096
rect 13596 12056 13728 12084
rect 13596 12044 13602 12056
rect 13722 12044 13728 12056
rect 13780 12084 13786 12096
rect 14384 12084 14412 12183
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15764 12152 15792 12251
rect 17494 12180 17500 12232
rect 17552 12180 17558 12232
rect 17972 12229 18000 12260
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 18690 12288 18696 12300
rect 18279 12260 18696 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 19610 12248 19616 12300
rect 19668 12248 19674 12300
rect 22296 12297 22324 12328
rect 23017 12325 23029 12328
rect 23063 12356 23075 12359
rect 23063 12328 23704 12356
rect 23063 12325 23075 12328
rect 23017 12319 23075 12325
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 23106 12248 23112 12300
rect 23164 12248 23170 12300
rect 23201 12291 23259 12297
rect 23201 12257 23213 12291
rect 23247 12288 23259 12291
rect 23474 12288 23480 12300
rect 23247 12260 23480 12288
rect 23247 12257 23259 12260
rect 23201 12251 23259 12257
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12220 18935 12223
rect 19150 12220 19156 12232
rect 18923 12192 19156 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 16942 12152 16948 12164
rect 15120 12124 15792 12152
rect 16790 12124 16948 12152
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 13780 12056 15025 12084
rect 13780 12044 13786 12056
rect 15013 12053 15025 12056
rect 15059 12084 15071 12087
rect 15120 12084 15148 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17221 12155 17279 12161
rect 17221 12121 17233 12155
rect 17267 12121 17279 12155
rect 17221 12115 17279 12121
rect 15059 12056 15148 12084
rect 17236 12084 17264 12115
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 19058 12152 19064 12164
rect 18656 12124 19064 12152
rect 18656 12112 18662 12124
rect 19058 12112 19064 12124
rect 19116 12152 19122 12164
rect 19352 12152 19380 12183
rect 20714 12180 20720 12232
rect 20772 12180 20778 12232
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12220 22247 12223
rect 22925 12223 22983 12229
rect 22925 12220 22937 12223
rect 22235 12192 22937 12220
rect 22235 12189 22247 12192
rect 22189 12183 22247 12189
rect 22925 12189 22937 12192
rect 22971 12189 22983 12223
rect 22925 12183 22983 12189
rect 19116 12124 19380 12152
rect 22940 12152 22968 12183
rect 23382 12180 23388 12232
rect 23440 12180 23446 12232
rect 23676 12229 23704 12328
rect 24486 12316 24492 12368
rect 24544 12356 24550 12368
rect 25041 12359 25099 12365
rect 25041 12356 25053 12359
rect 24544 12328 25053 12356
rect 24544 12316 24550 12328
rect 25041 12325 25053 12328
rect 25087 12325 25099 12359
rect 25041 12319 25099 12325
rect 28169 12359 28227 12365
rect 28169 12325 28181 12359
rect 28215 12356 28227 12359
rect 28534 12356 28540 12368
rect 28215 12328 28540 12356
rect 28215 12325 28227 12328
rect 28169 12319 28227 12325
rect 28534 12316 28540 12328
rect 28592 12316 28598 12368
rect 24946 12288 24952 12300
rect 24412 12260 24952 12288
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12220 23719 12223
rect 23750 12220 23756 12232
rect 23707 12192 23756 12220
rect 23707 12189 23719 12192
rect 23661 12183 23719 12189
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 23934 12180 23940 12232
rect 23992 12180 23998 12232
rect 24412 12229 24440 12260
rect 24946 12248 24952 12260
rect 25004 12288 25010 12300
rect 25409 12291 25467 12297
rect 25409 12288 25421 12291
rect 25004 12260 25421 12288
rect 25004 12248 25010 12260
rect 25409 12257 25421 12260
rect 25455 12257 25467 12291
rect 25409 12251 25467 12257
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12220 24087 12223
rect 24397 12223 24455 12229
rect 24075 12192 24256 12220
rect 24075 12189 24087 12192
rect 24029 12183 24087 12189
rect 23842 12152 23848 12164
rect 22940 12124 23848 12152
rect 19116 12112 19122 12124
rect 17589 12087 17647 12093
rect 17589 12084 17601 12087
rect 17236 12056 17601 12084
rect 15059 12053 15071 12056
rect 15013 12047 15071 12053
rect 17589 12053 17601 12056
rect 17635 12053 17647 12087
rect 17589 12047 17647 12053
rect 18049 12087 18107 12093
rect 18049 12053 18061 12087
rect 18095 12084 18107 12087
rect 18414 12084 18420 12096
rect 18095 12056 18420 12084
rect 18095 12053 18107 12056
rect 18049 12047 18107 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18969 12087 19027 12093
rect 18969 12053 18981 12087
rect 19015 12084 19027 12087
rect 20346 12084 20352 12096
rect 19015 12056 20352 12084
rect 19015 12053 19027 12056
rect 18969 12047 19027 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 21821 12087 21879 12093
rect 21821 12053 21833 12087
rect 21867 12084 21879 12087
rect 22002 12084 22008 12096
rect 21867 12056 22008 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 22741 12087 22799 12093
rect 22741 12053 22753 12087
rect 22787 12084 22799 12087
rect 23198 12084 23204 12096
rect 22787 12056 23204 12084
rect 22787 12053 22799 12056
rect 22741 12047 22799 12053
rect 23198 12044 23204 12056
rect 23256 12044 23262 12096
rect 23768 12093 23796 12124
rect 23842 12112 23848 12124
rect 23900 12112 23906 12164
rect 24118 12112 24124 12164
rect 24176 12112 24182 12164
rect 24228 12152 24256 12192
rect 24397 12189 24409 12223
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24670 12180 24676 12232
rect 24728 12180 24734 12232
rect 25501 12223 25559 12229
rect 25501 12220 25513 12223
rect 24964 12192 25513 12220
rect 24578 12152 24584 12164
rect 24228 12124 24584 12152
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 24964 12096 24992 12192
rect 25501 12189 25513 12192
rect 25547 12189 25559 12223
rect 25501 12183 25559 12189
rect 26510 12180 26516 12232
rect 26568 12220 26574 12232
rect 28644 12220 28672 12396
rect 29365 12393 29377 12396
rect 29411 12424 29423 12427
rect 30190 12424 30196 12436
rect 29411 12396 30196 12424
rect 29411 12393 29423 12396
rect 29365 12387 29423 12393
rect 30190 12384 30196 12396
rect 30248 12384 30254 12436
rect 31021 12427 31079 12433
rect 31021 12424 31033 12427
rect 30576 12396 31033 12424
rect 28718 12316 28724 12368
rect 28776 12316 28782 12368
rect 28810 12316 28816 12368
rect 28868 12316 28874 12368
rect 29822 12316 29828 12368
rect 29880 12316 29886 12368
rect 28736 12288 28764 12316
rect 28736 12260 29040 12288
rect 29012 12229 29040 12260
rect 28721 12223 28779 12229
rect 28721 12220 28733 12223
rect 26568 12192 28580 12220
rect 28644 12192 28733 12220
rect 26568 12180 26574 12192
rect 26605 12155 26663 12161
rect 26605 12121 26617 12155
rect 26651 12121 26663 12155
rect 26605 12115 26663 12121
rect 23753 12087 23811 12093
rect 23753 12053 23765 12087
rect 23799 12084 23811 12087
rect 24486 12084 24492 12096
rect 23799 12056 24492 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 24486 12044 24492 12056
rect 24544 12044 24550 12096
rect 24946 12044 24952 12096
rect 25004 12044 25010 12096
rect 25682 12044 25688 12096
rect 25740 12044 25746 12096
rect 26620 12084 26648 12115
rect 26786 12112 26792 12164
rect 26844 12161 26850 12164
rect 26844 12155 26863 12161
rect 26851 12121 26863 12155
rect 26844 12115 26863 12121
rect 26844 12112 26850 12115
rect 27522 12112 27528 12164
rect 27580 12152 27586 12164
rect 28552 12152 28580 12192
rect 28721 12189 28733 12192
rect 28767 12189 28779 12223
rect 28721 12183 28779 12189
rect 28997 12223 29055 12229
rect 28997 12189 29009 12223
rect 29043 12189 29055 12223
rect 28997 12183 29055 12189
rect 29641 12223 29699 12229
rect 29641 12189 29653 12223
rect 29687 12220 29699 12223
rect 29730 12220 29736 12232
rect 29687 12192 29736 12220
rect 29687 12189 29699 12192
rect 29641 12183 29699 12189
rect 29730 12180 29736 12192
rect 29788 12180 29794 12232
rect 30576 12229 30604 12396
rect 31021 12393 31033 12396
rect 31067 12424 31079 12427
rect 31202 12424 31208 12436
rect 31067 12396 31208 12424
rect 31067 12393 31079 12396
rect 31021 12387 31079 12393
rect 31202 12384 31208 12396
rect 31260 12424 31266 12436
rect 31297 12427 31355 12433
rect 31297 12424 31309 12427
rect 31260 12396 31309 12424
rect 31260 12384 31266 12396
rect 31297 12393 31309 12396
rect 31343 12393 31355 12427
rect 31297 12387 31355 12393
rect 32493 12427 32551 12433
rect 32493 12393 32505 12427
rect 32539 12424 32551 12427
rect 33502 12424 33508 12436
rect 32539 12396 33508 12424
rect 32539 12393 32551 12396
rect 32493 12387 32551 12393
rect 33502 12384 33508 12396
rect 33560 12384 33566 12436
rect 36262 12384 36268 12436
rect 36320 12424 36326 12436
rect 36633 12427 36691 12433
rect 36633 12424 36645 12427
rect 36320 12396 36645 12424
rect 36320 12384 36326 12396
rect 36633 12393 36645 12396
rect 36679 12393 36691 12427
rect 36633 12387 36691 12393
rect 31386 12316 31392 12368
rect 31444 12356 31450 12368
rect 31573 12359 31631 12365
rect 31573 12356 31585 12359
rect 31444 12328 31585 12356
rect 31444 12316 31450 12328
rect 31573 12325 31585 12328
rect 31619 12325 31631 12359
rect 31573 12319 31631 12325
rect 32674 12316 32680 12368
rect 32732 12316 32738 12368
rect 34885 12359 34943 12365
rect 34885 12325 34897 12359
rect 34931 12356 34943 12359
rect 34931 12328 35204 12356
rect 34931 12325 34943 12328
rect 34885 12319 34943 12325
rect 30760 12260 31800 12288
rect 30760 12232 30788 12260
rect 31772 12232 31800 12260
rect 32766 12248 32772 12300
rect 32824 12248 32830 12300
rect 33045 12291 33103 12297
rect 33045 12257 33057 12291
rect 33091 12288 33103 12291
rect 33134 12288 33140 12300
rect 33091 12260 33140 12288
rect 33091 12257 33103 12260
rect 33045 12251 33103 12257
rect 33134 12248 33140 12260
rect 33192 12248 33198 12300
rect 33410 12248 33416 12300
rect 33468 12288 33474 12300
rect 35176 12288 35204 12328
rect 36078 12316 36084 12368
rect 36136 12356 36142 12368
rect 36538 12356 36544 12368
rect 36136 12328 36544 12356
rect 36136 12316 36142 12328
rect 36538 12316 36544 12328
rect 36596 12316 36602 12368
rect 37458 12288 37464 12300
rect 33468 12260 35112 12288
rect 33468 12248 33474 12260
rect 30377 12223 30435 12229
rect 30377 12189 30389 12223
rect 30423 12189 30435 12223
rect 30377 12183 30435 12189
rect 30561 12223 30619 12229
rect 30561 12189 30573 12223
rect 30607 12189 30619 12223
rect 30561 12183 30619 12189
rect 29181 12155 29239 12161
rect 29181 12152 29193 12155
rect 27580 12124 28488 12152
rect 28552 12124 29193 12152
rect 27580 12112 27586 12124
rect 28350 12084 28356 12096
rect 26620 12056 28356 12084
rect 28350 12044 28356 12056
rect 28408 12044 28414 12096
rect 28460 12084 28488 12124
rect 29181 12121 29193 12124
rect 29227 12121 29239 12155
rect 30392 12152 30420 12183
rect 30742 12180 30748 12232
rect 30800 12180 30806 12232
rect 30837 12223 30895 12229
rect 30837 12189 30849 12223
rect 30883 12220 30895 12223
rect 30926 12220 30932 12232
rect 30883 12192 30932 12220
rect 30883 12189 30895 12192
rect 30837 12183 30895 12189
rect 30926 12180 30932 12192
rect 30984 12220 30990 12232
rect 31573 12223 31631 12229
rect 30984 12214 31524 12220
rect 31573 12214 31585 12223
rect 30984 12192 31585 12214
rect 30984 12180 30990 12192
rect 31496 12189 31585 12192
rect 31619 12189 31631 12223
rect 31496 12186 31631 12189
rect 31573 12183 31631 12186
rect 31754 12180 31760 12232
rect 31812 12180 31818 12232
rect 35084 12229 35112 12260
rect 35176 12260 37464 12288
rect 35069 12223 35127 12229
rect 35069 12189 35081 12223
rect 35115 12189 35127 12223
rect 35069 12183 35127 12189
rect 30392 12124 30972 12152
rect 29181 12115 29239 12121
rect 29089 12087 29147 12093
rect 29089 12084 29101 12087
rect 28460 12056 29101 12084
rect 29089 12053 29101 12056
rect 29135 12053 29147 12087
rect 29089 12047 29147 12053
rect 30469 12087 30527 12093
rect 30469 12053 30481 12087
rect 30515 12084 30527 12087
rect 30834 12084 30840 12096
rect 30515 12056 30840 12084
rect 30515 12053 30527 12056
rect 30469 12047 30527 12053
rect 30834 12044 30840 12056
rect 30892 12044 30898 12096
rect 30944 12084 30972 12124
rect 31018 12112 31024 12164
rect 31076 12152 31082 12164
rect 31113 12155 31171 12161
rect 31113 12152 31125 12155
rect 31076 12124 31125 12152
rect 31076 12112 31082 12124
rect 31113 12121 31125 12124
rect 31159 12121 31171 12155
rect 31113 12115 31171 12121
rect 31294 12112 31300 12164
rect 31352 12161 31358 12164
rect 31352 12155 31371 12161
rect 31359 12121 31371 12155
rect 31352 12115 31371 12121
rect 32309 12155 32367 12161
rect 32309 12121 32321 12155
rect 32355 12152 32367 12155
rect 32766 12152 32772 12164
rect 32355 12124 32772 12152
rect 32355 12121 32367 12124
rect 32309 12115 32367 12121
rect 31352 12112 31358 12115
rect 32766 12112 32772 12124
rect 32824 12112 32830 12164
rect 34330 12152 34336 12164
rect 34270 12124 34336 12152
rect 34330 12112 34336 12124
rect 34388 12152 34394 12164
rect 35176 12152 35204 12260
rect 37458 12248 37464 12260
rect 37516 12248 37522 12300
rect 35986 12180 35992 12232
rect 36044 12220 36050 12232
rect 36265 12223 36323 12229
rect 36265 12220 36277 12223
rect 36044 12192 36277 12220
rect 36044 12180 36050 12192
rect 36265 12189 36277 12192
rect 36311 12220 36323 12223
rect 36538 12220 36544 12232
rect 36311 12192 36544 12220
rect 36311 12189 36323 12192
rect 36265 12183 36323 12189
rect 36538 12180 36544 12192
rect 36596 12180 36602 12232
rect 36633 12223 36691 12229
rect 36633 12189 36645 12223
rect 36679 12189 36691 12223
rect 36633 12183 36691 12189
rect 36725 12223 36783 12229
rect 36725 12189 36737 12223
rect 36771 12220 36783 12223
rect 37090 12220 37096 12232
rect 36771 12192 37096 12220
rect 36771 12189 36783 12192
rect 36725 12183 36783 12189
rect 34388 12124 35204 12152
rect 34388 12112 34394 12124
rect 31202 12084 31208 12096
rect 30944 12056 31208 12084
rect 31202 12044 31208 12056
rect 31260 12044 31266 12096
rect 31481 12087 31539 12093
rect 31481 12053 31493 12087
rect 31527 12084 31539 12087
rect 31662 12084 31668 12096
rect 31527 12056 31668 12084
rect 31527 12053 31539 12056
rect 31481 12047 31539 12053
rect 31662 12044 31668 12056
rect 31720 12084 31726 12096
rect 32509 12087 32567 12093
rect 32509 12084 32521 12087
rect 31720 12056 32521 12084
rect 31720 12044 31726 12056
rect 32509 12053 32521 12056
rect 32555 12053 32567 12087
rect 32784 12084 32812 12112
rect 34517 12087 34575 12093
rect 34517 12084 34529 12087
rect 32784 12056 34529 12084
rect 32509 12047 32567 12053
rect 34517 12053 34529 12056
rect 34563 12053 34575 12087
rect 34517 12047 34575 12053
rect 35342 12044 35348 12096
rect 35400 12084 35406 12096
rect 35713 12087 35771 12093
rect 35713 12084 35725 12087
rect 35400 12056 35725 12084
rect 35400 12044 35406 12056
rect 35713 12053 35725 12056
rect 35759 12084 35771 12087
rect 36354 12084 36360 12096
rect 35759 12056 36360 12084
rect 35759 12053 35771 12056
rect 35713 12047 35771 12053
rect 36354 12044 36360 12056
rect 36412 12044 36418 12096
rect 36446 12044 36452 12096
rect 36504 12044 36510 12096
rect 36648 12084 36676 12183
rect 37090 12180 37096 12192
rect 37148 12180 37154 12232
rect 36814 12112 36820 12164
rect 36872 12152 36878 12164
rect 36909 12155 36967 12161
rect 36909 12152 36921 12155
rect 36872 12124 36921 12152
rect 36872 12112 36878 12124
rect 36909 12121 36921 12124
rect 36955 12121 36967 12155
rect 36909 12115 36967 12121
rect 36998 12084 37004 12096
rect 36648 12056 37004 12084
rect 36998 12044 37004 12056
rect 37056 12044 37062 12096
rect 1104 11994 38824 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 38824 11994
rect 1104 11920 38824 11942
rect 4430 11840 4436 11892
rect 4488 11840 4494 11892
rect 7742 11880 7748 11892
rect 4632 11852 7748 11880
rect 2958 11704 2964 11756
rect 3016 11704 3022 11756
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3694 11744 3700 11756
rect 3283 11716 3700 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3694 11704 3700 11716
rect 3752 11744 3758 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 3752 11716 4077 11744
rect 3752 11704 3758 11716
rect 4065 11713 4077 11716
rect 4111 11744 4123 11747
rect 4632 11744 4660 11852
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 9585 11883 9643 11889
rect 8260 11852 9444 11880
rect 8260 11840 8266 11852
rect 5442 11772 5448 11824
rect 5500 11772 5506 11824
rect 6365 11815 6423 11821
rect 6365 11781 6377 11815
rect 6411 11812 6423 11815
rect 7006 11812 7012 11824
rect 6411 11784 7012 11812
rect 6411 11781 6423 11784
rect 6365 11775 6423 11781
rect 7006 11772 7012 11784
rect 7064 11812 7070 11824
rect 7377 11815 7435 11821
rect 7377 11812 7389 11815
rect 7064 11784 7389 11812
rect 7064 11772 7070 11784
rect 7377 11781 7389 11784
rect 7423 11781 7435 11815
rect 7377 11775 7435 11781
rect 8113 11815 8171 11821
rect 8113 11781 8125 11815
rect 8159 11812 8171 11815
rect 8386 11812 8392 11824
rect 8159 11784 8392 11812
rect 8159 11781 8171 11784
rect 8113 11775 8171 11781
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 9416 11812 9444 11852
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 9766 11880 9772 11892
rect 9631 11852 9772 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10870 11840 10876 11892
rect 10928 11840 10934 11892
rect 12894 11880 12900 11892
rect 11256 11852 12900 11880
rect 10042 11812 10048 11824
rect 9338 11784 10048 11812
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10888 11812 10916 11840
rect 11149 11815 11207 11821
rect 11149 11812 11161 11815
rect 10888 11784 11161 11812
rect 11149 11781 11161 11784
rect 11195 11781 11207 11815
rect 11149 11775 11207 11781
rect 4111 11716 4660 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4338 11636 4344 11688
rect 4396 11636 4402 11688
rect 5902 11636 5908 11688
rect 5960 11636 5966 11688
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 6546 11676 6552 11688
rect 6236 11648 6552 11676
rect 6236 11636 6242 11648
rect 6546 11636 6552 11648
rect 6604 11676 6610 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 6604 11648 7205 11676
rect 6604 11636 6610 11648
rect 7193 11645 7205 11648
rect 7239 11676 7251 11679
rect 7834 11676 7840 11688
rect 7239 11648 7840 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 11256 11676 11284 11852
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 17678 11880 17684 11892
rect 17328 11852 17684 11880
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 13096 11812 13124 11840
rect 13265 11815 13323 11821
rect 13265 11812 13277 11815
rect 11940 11784 12098 11812
rect 13096 11784 13277 11812
rect 11940 11772 11946 11784
rect 13265 11781 13277 11784
rect 13311 11781 13323 11815
rect 13265 11775 13323 11781
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 17328 11812 17356 11852
rect 17678 11840 17684 11852
rect 17736 11880 17742 11892
rect 17736 11852 18276 11880
rect 17736 11840 17742 11852
rect 18248 11812 18276 11852
rect 18414 11840 18420 11892
rect 18472 11840 18478 11892
rect 20349 11883 20407 11889
rect 20349 11849 20361 11883
rect 20395 11880 20407 11883
rect 20438 11880 20444 11892
rect 20395 11852 20444 11880
rect 20395 11849 20407 11852
rect 20349 11843 20407 11849
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 23017 11883 23075 11889
rect 23017 11849 23029 11883
rect 23063 11880 23075 11883
rect 23934 11880 23940 11892
rect 23063 11852 23940 11880
rect 23063 11849 23075 11852
rect 23017 11843 23075 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 33226 11840 33232 11892
rect 33284 11840 33290 11892
rect 34790 11840 34796 11892
rect 34848 11880 34854 11892
rect 35069 11883 35127 11889
rect 35069 11880 35081 11883
rect 34848 11852 35081 11880
rect 34848 11840 34854 11852
rect 35069 11849 35081 11852
rect 35115 11849 35127 11883
rect 35069 11843 35127 11849
rect 17000 11784 17434 11812
rect 18248 11784 19366 11812
rect 17000 11772 17006 11784
rect 23382 11772 23388 11824
rect 23440 11812 23446 11824
rect 27065 11815 27123 11821
rect 27065 11812 27077 11815
rect 23440 11784 23796 11812
rect 23440 11772 23446 11784
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11744 13691 11747
rect 13722 11744 13728 11756
rect 13679 11716 13728 11744
rect 13679 11713 13691 11716
rect 13633 11707 13691 11713
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11744 13875 11747
rect 13906 11744 13912 11756
rect 13863 11716 13912 11744
rect 13863 11713 13875 11716
rect 13817 11707 13875 11713
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 7944 11648 11284 11676
rect 11793 11679 11851 11685
rect 3418 11568 3424 11620
rect 3476 11568 3482 11620
rect 4522 11568 4528 11620
rect 4580 11608 4586 11620
rect 4580 11580 4844 11608
rect 4580 11568 4586 11580
rect 4816 11552 4844 11580
rect 2866 11500 2872 11552
rect 2924 11500 2930 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 4706 11540 4712 11552
rect 3660 11512 4712 11540
rect 3660 11500 3666 11512
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 7944 11540 7972 11648
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 12802 11676 12808 11688
rect 11839 11648 12808 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11676 13599 11679
rect 14090 11676 14096 11688
rect 13587 11648 14096 11676
rect 13587 11645 13599 11648
rect 13541 11639 13599 11645
rect 14090 11636 14096 11648
rect 14148 11676 14154 11688
rect 16224 11676 16252 11707
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 20441 11747 20499 11753
rect 20441 11744 20453 11747
rect 20404 11716 20453 11744
rect 20404 11704 20410 11716
rect 20441 11713 20453 11716
rect 20487 11713 20499 11747
rect 20441 11707 20499 11713
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22557 11747 22615 11753
rect 22557 11744 22569 11747
rect 22060 11716 22569 11744
rect 22060 11704 22066 11716
rect 22557 11713 22569 11716
rect 22603 11713 22615 11747
rect 22557 11707 22615 11713
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 23768 11753 23796 11784
rect 26620 11784 27077 11812
rect 26620 11756 26648 11784
rect 27065 11781 27077 11784
rect 27111 11781 27123 11815
rect 27065 11775 27123 11781
rect 29730 11772 29736 11824
rect 29788 11812 29794 11824
rect 35342 11812 35348 11824
rect 29788 11784 35348 11812
rect 29788 11772 29794 11784
rect 35342 11772 35348 11784
rect 35400 11772 35406 11824
rect 36446 11812 36452 11824
rect 35452 11784 36452 11812
rect 23569 11747 23627 11753
rect 23569 11744 23581 11747
rect 23532 11716 23581 11744
rect 23532 11704 23538 11716
rect 23569 11713 23581 11716
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11713 23811 11747
rect 23753 11707 23811 11713
rect 16666 11676 16672 11688
rect 14148 11648 16672 11676
rect 14148 11636 14154 11648
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 16945 11679 17003 11685
rect 16945 11645 16957 11679
rect 16991 11676 17003 11679
rect 17402 11676 17408 11688
rect 16991 11648 17408 11676
rect 16991 11645 17003 11648
rect 16945 11639 17003 11645
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 17494 11636 17500 11688
rect 17552 11676 17558 11688
rect 18598 11676 18604 11688
rect 17552 11648 18604 11676
rect 17552 11636 17558 11648
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 19334 11676 19340 11688
rect 18923 11648 19340 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 19334 11636 19340 11648
rect 19392 11636 19398 11688
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11645 22155 11679
rect 23768 11676 23796 11707
rect 24670 11704 24676 11756
rect 24728 11704 24734 11756
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11744 24915 11747
rect 25682 11744 25688 11756
rect 24903 11716 25688 11744
rect 24903 11713 24915 11716
rect 24857 11707 24915 11713
rect 24302 11676 24308 11688
rect 23768 11648 24308 11676
rect 22097 11639 22155 11645
rect 13814 11568 13820 11620
rect 13872 11568 13878 11620
rect 21450 11608 21456 11620
rect 20456 11580 21456 11608
rect 4856 11512 7972 11540
rect 11241 11543 11299 11549
rect 4856 11500 4862 11512
rect 11241 11509 11253 11543
rect 11287 11540 11299 11543
rect 11606 11540 11612 11552
rect 11287 11512 11612 11540
rect 11287 11509 11299 11512
rect 11241 11503 11299 11509
rect 11606 11500 11612 11512
rect 11664 11540 11670 11552
rect 12618 11540 12624 11552
rect 11664 11512 12624 11540
rect 11664 11500 11670 11512
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 20456 11540 20484 11580
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 22112 11608 22140 11639
rect 24302 11636 24308 11648
rect 24360 11676 24366 11688
rect 24872 11676 24900 11707
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 25958 11704 25964 11756
rect 26016 11704 26022 11756
rect 26142 11704 26148 11756
rect 26200 11704 26206 11756
rect 26234 11704 26240 11756
rect 26292 11744 26298 11756
rect 26418 11744 26424 11756
rect 26292 11716 26424 11744
rect 26292 11704 26298 11716
rect 26418 11704 26424 11716
rect 26476 11704 26482 11756
rect 26513 11747 26571 11753
rect 26513 11713 26525 11747
rect 26559 11744 26571 11747
rect 26602 11744 26608 11756
rect 26559 11716 26608 11744
rect 26559 11713 26571 11716
rect 26513 11707 26571 11713
rect 26602 11704 26608 11716
rect 26660 11704 26666 11756
rect 26970 11704 26976 11756
rect 27028 11704 27034 11756
rect 27249 11747 27307 11753
rect 27249 11713 27261 11747
rect 27295 11713 27307 11747
rect 27249 11707 27307 11713
rect 30837 11747 30895 11753
rect 30837 11713 30849 11747
rect 30883 11744 30895 11747
rect 31018 11744 31024 11756
rect 30883 11716 31024 11744
rect 30883 11713 30895 11716
rect 30837 11707 30895 11713
rect 24360 11648 24900 11676
rect 26329 11679 26387 11685
rect 24360 11636 24366 11648
rect 26329 11645 26341 11679
rect 26375 11676 26387 11679
rect 26697 11679 26755 11685
rect 26375 11648 26648 11676
rect 26375 11645 26387 11648
rect 26329 11639 26387 11645
rect 26620 11620 26648 11648
rect 26697 11645 26709 11679
rect 26743 11676 26755 11679
rect 27264 11676 27292 11707
rect 31018 11704 31024 11716
rect 31076 11704 31082 11756
rect 31478 11704 31484 11756
rect 31536 11744 31542 11756
rect 33045 11747 33103 11753
rect 33045 11744 33057 11747
rect 31536 11716 33057 11744
rect 31536 11704 31542 11716
rect 33045 11713 33057 11716
rect 33091 11713 33103 11747
rect 33045 11707 33103 11713
rect 34790 11704 34796 11756
rect 34848 11744 34854 11756
rect 35452 11753 35480 11784
rect 36446 11772 36452 11784
rect 36504 11772 36510 11824
rect 36722 11772 36728 11824
rect 36780 11812 36786 11824
rect 37461 11815 37519 11821
rect 37461 11812 37473 11815
rect 36780 11784 37473 11812
rect 36780 11772 36786 11784
rect 37461 11781 37473 11784
rect 37507 11781 37519 11815
rect 37461 11775 37519 11781
rect 35253 11747 35311 11753
rect 35253 11744 35265 11747
rect 34848 11716 35265 11744
rect 34848 11704 34854 11716
rect 35253 11713 35265 11716
rect 35299 11713 35311 11747
rect 35253 11707 35311 11713
rect 35437 11747 35495 11753
rect 35437 11713 35449 11747
rect 35483 11713 35495 11747
rect 35437 11707 35495 11713
rect 35529 11747 35587 11753
rect 35529 11713 35541 11747
rect 35575 11713 35587 11747
rect 35529 11707 35587 11713
rect 26743 11648 27292 11676
rect 30929 11679 30987 11685
rect 26743 11645 26755 11648
rect 26697 11639 26755 11645
rect 30929 11645 30941 11679
rect 30975 11676 30987 11679
rect 31386 11676 31392 11688
rect 30975 11648 31392 11676
rect 30975 11645 30987 11648
rect 30929 11639 30987 11645
rect 31386 11636 31392 11648
rect 31444 11636 31450 11688
rect 32766 11636 32772 11688
rect 32824 11636 32830 11688
rect 32861 11679 32919 11685
rect 32861 11645 32873 11679
rect 32907 11645 32919 11679
rect 32861 11639 32919 11645
rect 32953 11679 33011 11685
rect 32953 11645 32965 11679
rect 32999 11676 33011 11679
rect 33226 11676 33232 11688
rect 32999 11648 33232 11676
rect 32999 11645 33011 11648
rect 32953 11639 33011 11645
rect 22925 11611 22983 11617
rect 22925 11608 22937 11611
rect 22112 11580 22937 11608
rect 22925 11577 22937 11580
rect 22971 11608 22983 11611
rect 23106 11608 23112 11620
rect 22971 11580 23112 11608
rect 22971 11577 22983 11580
rect 22925 11571 22983 11577
rect 23106 11568 23112 11580
rect 23164 11568 23170 11620
rect 26602 11568 26608 11620
rect 26660 11608 26666 11620
rect 26970 11608 26976 11620
rect 26660 11580 26976 11608
rect 26660 11568 26666 11580
rect 26970 11568 26976 11580
rect 27028 11568 27034 11620
rect 31205 11611 31263 11617
rect 31205 11577 31217 11611
rect 31251 11608 31263 11611
rect 31570 11608 31576 11620
rect 31251 11580 31576 11608
rect 31251 11577 31263 11580
rect 31205 11571 31263 11577
rect 31570 11568 31576 11580
rect 31628 11568 31634 11620
rect 32876 11608 32904 11639
rect 33226 11636 33232 11648
rect 33284 11636 33290 11688
rect 35544 11676 35572 11707
rect 35710 11704 35716 11756
rect 35768 11704 35774 11756
rect 35805 11747 35863 11753
rect 35805 11713 35817 11747
rect 35851 11744 35863 11747
rect 36354 11744 36360 11756
rect 35851 11716 36360 11744
rect 35851 11713 35863 11716
rect 35805 11707 35863 11713
rect 36354 11704 36360 11716
rect 36412 11704 36418 11756
rect 36170 11676 36176 11688
rect 35544 11648 36176 11676
rect 36170 11636 36176 11648
rect 36228 11636 36234 11688
rect 36630 11636 36636 11688
rect 36688 11636 36694 11688
rect 33594 11608 33600 11620
rect 32876 11580 33600 11608
rect 33594 11568 33600 11580
rect 33652 11568 33658 11620
rect 35342 11568 35348 11620
rect 35400 11568 35406 11620
rect 37826 11568 37832 11620
rect 37884 11568 37890 11620
rect 12952 11512 20484 11540
rect 20625 11543 20683 11549
rect 12952 11500 12958 11512
rect 20625 11509 20637 11543
rect 20671 11540 20683 11543
rect 21266 11540 21272 11552
rect 20671 11512 21272 11540
rect 20671 11509 20683 11512
rect 20625 11503 20683 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 22278 11500 22284 11552
rect 22336 11500 22342 11552
rect 23569 11543 23627 11549
rect 23569 11509 23581 11543
rect 23615 11540 23627 11543
rect 24578 11540 24584 11552
rect 23615 11512 24584 11540
rect 23615 11509 23627 11512
rect 23569 11503 23627 11509
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 24857 11543 24915 11549
rect 24857 11509 24869 11543
rect 24903 11540 24915 11543
rect 25038 11540 25044 11552
rect 24903 11512 25044 11540
rect 24903 11509 24915 11512
rect 24857 11503 24915 11509
rect 25038 11500 25044 11512
rect 25096 11500 25102 11552
rect 27433 11543 27491 11549
rect 27433 11509 27445 11543
rect 27479 11540 27491 11543
rect 28258 11540 28264 11552
rect 27479 11512 28264 11540
rect 27479 11509 27491 11512
rect 27433 11503 27491 11509
rect 28258 11500 28264 11512
rect 28316 11500 28322 11552
rect 32674 11500 32680 11552
rect 32732 11540 32738 11552
rect 34422 11540 34428 11552
rect 32732 11512 34428 11540
rect 32732 11500 32738 11512
rect 34422 11500 34428 11512
rect 34480 11540 34486 11552
rect 36538 11540 36544 11552
rect 34480 11512 36544 11540
rect 34480 11500 34486 11512
rect 36538 11500 36544 11512
rect 36596 11500 36602 11552
rect 36906 11500 36912 11552
rect 36964 11540 36970 11552
rect 37277 11543 37335 11549
rect 37277 11540 37289 11543
rect 36964 11512 37289 11540
rect 36964 11500 36970 11512
rect 37277 11509 37289 11512
rect 37323 11509 37335 11543
rect 37277 11503 37335 11509
rect 37366 11500 37372 11552
rect 37424 11540 37430 11552
rect 37461 11543 37519 11549
rect 37461 11540 37473 11543
rect 37424 11512 37473 11540
rect 37424 11500 37430 11512
rect 37461 11509 37473 11512
rect 37507 11509 37519 11543
rect 37461 11503 37519 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 2915 11308 3924 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 2498 11228 2504 11280
rect 2556 11268 2562 11280
rect 2556 11240 3832 11268
rect 2556 11228 2562 11240
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11200 2651 11203
rect 2958 11200 2964 11212
rect 2639 11172 2964 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3602 11160 3608 11212
rect 3660 11160 3666 11212
rect 1302 11092 1308 11144
rect 1360 11132 1366 11144
rect 3804 11141 3832 11240
rect 3896 11200 3924 11308
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 4672 11308 5120 11336
rect 4672 11296 4678 11308
rect 5092 11268 5120 11308
rect 5350 11296 5356 11348
rect 5408 11336 5414 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 5408 11308 5549 11336
rect 5408 11296 5414 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 5537 11299 5595 11305
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6512 11308 6929 11336
rect 6512 11296 6518 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 17034 11336 17040 11348
rect 12299 11308 12572 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 5258 11268 5264 11280
rect 5092 11240 5264 11268
rect 5258 11228 5264 11240
rect 5316 11268 5322 11280
rect 5316 11240 6684 11268
rect 5316 11228 5322 11240
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3896 11172 4077 11200
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4798 11200 4804 11212
rect 4212 11172 4804 11200
rect 4212 11160 4218 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 5902 11160 5908 11212
rect 5960 11200 5966 11212
rect 6549 11203 6607 11209
rect 6549 11200 6561 11203
rect 5960 11172 6561 11200
rect 5960 11160 5966 11172
rect 6549 11169 6561 11172
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 6656 11141 6684 11240
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 12345 11271 12403 11277
rect 7892 11240 9076 11268
rect 7892 11228 7898 11240
rect 7374 11160 7380 11212
rect 7432 11160 7438 11212
rect 8110 11160 8116 11212
rect 8168 11200 8174 11212
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 8168 11172 8217 11200
rect 8168 11160 8174 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 9048 11144 9076 11240
rect 12345 11237 12357 11271
rect 12391 11237 12403 11271
rect 12345 11231 12403 11237
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11200 10839 11203
rect 12360 11200 12388 11231
rect 10827 11172 12388 11200
rect 12544 11200 12572 11308
rect 14200 11308 17040 11336
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 14200 11268 14228 11308
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17126 11296 17132 11348
rect 17184 11296 17190 11348
rect 17402 11296 17408 11348
rect 17460 11296 17466 11348
rect 17678 11296 17684 11348
rect 17736 11336 17742 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 17736 11308 18337 11336
rect 17736 11296 17742 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18325 11299 18383 11305
rect 21637 11339 21695 11345
rect 21637 11305 21649 11339
rect 21683 11336 21695 11339
rect 21818 11336 21824 11348
rect 21683 11308 21824 11336
rect 21683 11305 21695 11308
rect 21637 11299 21695 11305
rect 12676 11240 14228 11268
rect 17144 11268 17172 11296
rect 17144 11240 17724 11268
rect 12676 11228 12682 11240
rect 12544 11172 12756 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 1397 11135 1455 11141
rect 1397 11132 1409 11135
rect 1360 11104 1409 11132
rect 1360 11092 1366 11104
rect 1397 11101 1409 11104
rect 1443 11132 1455 11135
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1443 11104 1685 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11132 6423 11135
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 6411 11104 6469 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 7331 11104 7665 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7653 11101 7665 11104
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 2516 11064 2544 11095
rect 3694 11064 3700 11076
rect 2516 11036 3700 11064
rect 3694 11024 3700 11036
rect 3752 11024 3758 11076
rect 3804 11064 3832 11095
rect 8386 11092 8392 11144
rect 8444 11092 8450 11144
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 8662 11132 8668 11144
rect 8619 11104 8668 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 9088 11104 10517 11132
rect 9088 11092 9094 11104
rect 10505 11101 10517 11104
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 11882 11092 11888 11144
rect 11940 11092 11946 11144
rect 12728 11141 12756 11172
rect 12802 11160 12808 11212
rect 12860 11160 12866 11212
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 13170 11200 13176 11212
rect 13035 11172 13176 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 14918 11160 14924 11212
rect 14976 11200 14982 11212
rect 15841 11203 15899 11209
rect 15841 11200 15853 11203
rect 14976 11172 15853 11200
rect 14976 11160 14982 11172
rect 15841 11169 15853 11172
rect 15887 11169 15899 11203
rect 15841 11163 15899 11169
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 17129 11203 17187 11209
rect 17129 11200 17141 11203
rect 16724 11172 17141 11200
rect 16724 11160 16730 11172
rect 17129 11169 17141 11172
rect 17175 11200 17187 11203
rect 17586 11200 17592 11212
rect 17175 11172 17592 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 17696 11200 17724 11240
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 17696 11172 17969 11200
rect 17957 11169 17969 11172
rect 18003 11169 18015 11203
rect 21652 11200 21680 11299
rect 21818 11296 21824 11308
rect 21876 11336 21882 11348
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 21876 11308 22017 11336
rect 21876 11296 21882 11308
rect 22005 11305 22017 11308
rect 22051 11336 22063 11339
rect 22281 11339 22339 11345
rect 22281 11336 22293 11339
rect 22051 11308 22293 11336
rect 22051 11305 22063 11308
rect 22005 11299 22063 11305
rect 22281 11305 22293 11308
rect 22327 11336 22339 11339
rect 22327 11308 24992 11336
rect 22327 11305 22339 11308
rect 22281 11299 22339 11305
rect 17957 11163 18015 11169
rect 21284 11172 21680 11200
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11132 12771 11135
rect 13354 11132 13360 11144
rect 12759 11104 13360 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 14090 11092 14096 11144
rect 14148 11092 14154 11144
rect 15470 11092 15476 11144
rect 15528 11092 15534 11144
rect 17770 11132 17776 11144
rect 16592 11104 17776 11132
rect 16592 11076 16620 11104
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 17880 11104 18613 11132
rect 3804 11036 4016 11064
rect 1578 10956 1584 11008
rect 1636 10956 1642 11008
rect 3988 10996 4016 11036
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4120 11036 4554 11064
rect 4120 11024 4126 11036
rect 14366 11024 14372 11076
rect 14424 11024 14430 11076
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 16301 11067 16359 11073
rect 16301 11064 16313 11067
rect 16264 11036 16313 11064
rect 16264 11024 16270 11036
rect 16301 11033 16313 11036
rect 16347 11064 16359 11067
rect 16393 11067 16451 11073
rect 16393 11064 16405 11067
rect 16347 11036 16405 11064
rect 16347 11033 16359 11036
rect 16301 11027 16359 11033
rect 16393 11033 16405 11036
rect 16439 11064 16451 11067
rect 16574 11064 16580 11076
rect 16439 11036 16580 11064
rect 16439 11033 16451 11036
rect 16393 11027 16451 11033
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 17880 11064 17908 11104
rect 18601 11101 18613 11104
rect 18647 11132 18659 11135
rect 18782 11132 18788 11144
rect 18647 11104 18788 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 21284 11141 21312 11172
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 21450 11092 21456 11144
rect 21508 11132 21514 11144
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 21508 11104 21833 11132
rect 21508 11092 21514 11104
rect 21821 11101 21833 11104
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 24210 11092 24216 11144
rect 24268 11132 24274 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 24268 11104 24409 11132
rect 24268 11092 24274 11104
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24578 11092 24584 11144
rect 24636 11092 24642 11144
rect 24854 11092 24860 11144
rect 24912 11092 24918 11144
rect 17092 11036 17908 11064
rect 20901 11067 20959 11073
rect 17092 11024 17098 11036
rect 20901 11033 20913 11067
rect 20947 11064 20959 11067
rect 20990 11064 20996 11076
rect 20947 11036 20996 11064
rect 20947 11033 20959 11036
rect 20901 11027 20959 11033
rect 20990 11024 20996 11036
rect 21048 11024 21054 11076
rect 24118 11024 24124 11076
rect 24176 11064 24182 11076
rect 24765 11067 24823 11073
rect 24765 11064 24777 11067
rect 24176 11036 24777 11064
rect 24176 11024 24182 11036
rect 24765 11033 24777 11036
rect 24811 11033 24823 11067
rect 24964 11064 24992 11308
rect 25958 11296 25964 11348
rect 26016 11296 26022 11348
rect 28537 11339 28595 11345
rect 28537 11305 28549 11339
rect 28583 11336 28595 11339
rect 30190 11336 30196 11348
rect 28583 11308 30196 11336
rect 28583 11305 28595 11308
rect 28537 11299 28595 11305
rect 30190 11296 30196 11308
rect 30248 11296 30254 11348
rect 31754 11296 31760 11348
rect 31812 11336 31818 11348
rect 32769 11339 32827 11345
rect 32769 11336 32781 11339
rect 31812 11308 32781 11336
rect 31812 11296 31818 11308
rect 32769 11305 32781 11308
rect 32815 11305 32827 11339
rect 32769 11299 32827 11305
rect 27617 11271 27675 11277
rect 27617 11237 27629 11271
rect 27663 11268 27675 11271
rect 28353 11271 28411 11277
rect 28353 11268 28365 11271
rect 27663 11240 28365 11268
rect 27663 11237 27675 11240
rect 27617 11231 27675 11237
rect 28353 11237 28365 11240
rect 28399 11237 28411 11271
rect 28629 11271 28687 11277
rect 28629 11268 28641 11271
rect 28353 11231 28411 11237
rect 28460 11240 28641 11268
rect 28258 11160 28264 11212
rect 28316 11200 28322 11212
rect 28460 11200 28488 11240
rect 28629 11237 28641 11240
rect 28675 11237 28687 11271
rect 30926 11268 30932 11280
rect 28629 11231 28687 11237
rect 29932 11240 30932 11268
rect 28316 11172 28488 11200
rect 28316 11160 28322 11172
rect 28534 11160 28540 11212
rect 28592 11200 28598 11212
rect 29932 11209 29960 11240
rect 30926 11228 30932 11240
rect 30984 11228 30990 11280
rect 29917 11203 29975 11209
rect 28592 11172 29040 11200
rect 28592 11160 28598 11172
rect 25958 11092 25964 11144
rect 26016 11132 26022 11144
rect 26145 11135 26203 11141
rect 26145 11132 26157 11135
rect 26016 11104 26157 11132
rect 26016 11092 26022 11104
rect 26145 11101 26157 11104
rect 26191 11101 26203 11135
rect 26145 11095 26203 11101
rect 26234 11092 26240 11144
rect 26292 11092 26298 11144
rect 26326 11092 26332 11144
rect 26384 11132 26390 11144
rect 26421 11135 26479 11141
rect 26421 11132 26433 11135
rect 26384 11104 26433 11132
rect 26384 11092 26390 11104
rect 26421 11101 26433 11104
rect 26467 11101 26479 11135
rect 26421 11095 26479 11101
rect 26510 11092 26516 11144
rect 26568 11092 26574 11144
rect 27798 11092 27804 11144
rect 27856 11092 27862 11144
rect 27890 11092 27896 11144
rect 27948 11092 27954 11144
rect 28169 11135 28227 11141
rect 28169 11101 28181 11135
rect 28215 11132 28227 11135
rect 28721 11135 28779 11141
rect 28721 11132 28733 11135
rect 28215 11104 28733 11132
rect 28215 11101 28227 11104
rect 28169 11095 28227 11101
rect 28721 11101 28733 11104
rect 28767 11132 28779 11135
rect 28810 11132 28816 11144
rect 28767 11104 28816 11132
rect 28767 11101 28779 11104
rect 28721 11095 28779 11101
rect 28810 11092 28816 11104
rect 28868 11092 28874 11144
rect 29012 11141 29040 11172
rect 29917 11169 29929 11203
rect 29963 11169 29975 11203
rect 32784 11200 32812 11299
rect 32858 11296 32864 11348
rect 32916 11296 32922 11348
rect 33321 11339 33379 11345
rect 33321 11305 33333 11339
rect 33367 11336 33379 11339
rect 33594 11336 33600 11348
rect 33367 11308 33600 11336
rect 33367 11305 33379 11308
rect 33321 11299 33379 11305
rect 33594 11296 33600 11308
rect 33652 11296 33658 11348
rect 36078 11296 36084 11348
rect 36136 11296 36142 11348
rect 36170 11296 36176 11348
rect 36228 11296 36234 11348
rect 36262 11296 36268 11348
rect 36320 11296 36326 11348
rect 37090 11336 37096 11348
rect 36648 11308 37096 11336
rect 32876 11268 32904 11296
rect 36648 11268 36676 11308
rect 37090 11296 37096 11308
rect 37148 11296 37154 11348
rect 32876 11240 33364 11268
rect 29917 11163 29975 11169
rect 30116 11172 30696 11200
rect 32784 11172 33088 11200
rect 30116 11144 30144 11172
rect 28997 11135 29055 11141
rect 28997 11101 29009 11135
rect 29043 11101 29055 11135
rect 28997 11095 29055 11101
rect 30006 11092 30012 11144
rect 30064 11092 30070 11144
rect 30098 11092 30104 11144
rect 30156 11092 30162 11144
rect 30190 11092 30196 11144
rect 30248 11092 30254 11144
rect 30668 11141 30696 11172
rect 30469 11135 30527 11141
rect 30469 11101 30481 11135
rect 30515 11101 30527 11135
rect 30469 11095 30527 11101
rect 30653 11135 30711 11141
rect 30653 11101 30665 11135
rect 30699 11101 30711 11135
rect 30653 11095 30711 11101
rect 29086 11064 29092 11076
rect 24964 11036 29092 11064
rect 24765 11027 24823 11033
rect 29086 11024 29092 11036
rect 29144 11024 29150 11076
rect 29178 11024 29184 11076
rect 29236 11024 29242 11076
rect 30024 11064 30052 11092
rect 30484 11064 30512 11095
rect 31018 11092 31024 11144
rect 31076 11132 31082 11144
rect 32858 11132 32864 11144
rect 31076 11104 32864 11132
rect 31076 11092 31082 11104
rect 32858 11092 32864 11104
rect 32916 11092 32922 11144
rect 32950 11092 32956 11144
rect 33008 11092 33014 11144
rect 33060 11141 33088 11172
rect 33045 11135 33103 11141
rect 33045 11101 33057 11135
rect 33091 11101 33103 11135
rect 33045 11095 33103 11101
rect 33226 11092 33232 11144
rect 33284 11092 33290 11144
rect 33336 11141 33364 11240
rect 36280 11240 36676 11268
rect 35161 11203 35219 11209
rect 35161 11169 35173 11203
rect 35207 11200 35219 11203
rect 35207 11172 35848 11200
rect 35207 11169 35219 11172
rect 35161 11163 35219 11169
rect 33321 11135 33379 11141
rect 33321 11101 33333 11135
rect 33367 11132 33379 11135
rect 33870 11132 33876 11144
rect 33367 11104 33876 11132
rect 33367 11101 33379 11104
rect 33321 11095 33379 11101
rect 33870 11092 33876 11104
rect 33928 11092 33934 11144
rect 35820 11141 35848 11172
rect 36280 11144 36308 11240
rect 36906 11160 36912 11212
rect 36964 11160 36970 11212
rect 36998 11160 37004 11212
rect 37056 11200 37062 11212
rect 38381 11203 38439 11209
rect 38381 11200 38393 11203
rect 37056 11172 38393 11200
rect 37056 11160 37062 11172
rect 38381 11169 38393 11172
rect 38427 11169 38439 11203
rect 38381 11163 38439 11169
rect 35345 11135 35403 11141
rect 35345 11101 35357 11135
rect 35391 11101 35403 11135
rect 35345 11095 35403 11101
rect 35437 11135 35495 11141
rect 35437 11101 35449 11135
rect 35483 11101 35495 11135
rect 35437 11095 35495 11101
rect 35621 11135 35679 11141
rect 35621 11101 35633 11135
rect 35667 11101 35679 11135
rect 35621 11095 35679 11101
rect 35713 11135 35771 11141
rect 35713 11101 35725 11135
rect 35759 11101 35771 11135
rect 35713 11095 35771 11101
rect 35805 11135 35863 11141
rect 35805 11101 35817 11135
rect 35851 11101 35863 11135
rect 35805 11095 35863 11101
rect 35989 11135 36047 11141
rect 35989 11101 36001 11135
rect 36035 11132 36047 11135
rect 36262 11132 36268 11144
rect 36035 11104 36268 11132
rect 36035 11101 36047 11104
rect 35989 11095 36047 11101
rect 30024 11036 30512 11064
rect 30926 11024 30932 11076
rect 30984 11064 30990 11076
rect 32968 11064 32996 11092
rect 35360 11064 35388 11095
rect 30984 11036 32996 11064
rect 33520 11036 35388 11064
rect 30984 11024 30990 11036
rect 4798 10996 4804 11008
rect 3988 10968 4804 10996
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 8478 10956 8484 11008
rect 8536 10956 8542 11008
rect 17770 10956 17776 11008
rect 17828 10956 17834 11008
rect 17865 10999 17923 11005
rect 17865 10965 17877 10999
rect 17911 10996 17923 10999
rect 17954 10996 17960 11008
rect 17911 10968 17960 10996
rect 17911 10965 17923 10968
rect 17865 10959 17923 10965
rect 17954 10956 17960 10968
rect 18012 10996 18018 11008
rect 18414 10996 18420 11008
rect 18012 10968 18420 10996
rect 18012 10956 18018 10968
rect 18414 10956 18420 10968
rect 18472 10956 18478 11008
rect 22738 10956 22744 11008
rect 22796 10996 22802 11008
rect 26326 10996 26332 11008
rect 22796 10968 26332 10996
rect 22796 10956 22802 10968
rect 26326 10956 26332 10968
rect 26384 10996 26390 11008
rect 28074 10996 28080 11008
rect 26384 10968 28080 10996
rect 26384 10956 26390 10968
rect 28074 10956 28080 10968
rect 28132 10956 28138 11008
rect 29365 10999 29423 11005
rect 29365 10965 29377 10999
rect 29411 10996 29423 10999
rect 30098 10996 30104 11008
rect 29411 10968 30104 10996
rect 29411 10965 29423 10968
rect 29365 10959 29423 10965
rect 30098 10956 30104 10968
rect 30156 10956 30162 11008
rect 30377 10999 30435 11005
rect 30377 10965 30389 10999
rect 30423 10996 30435 10999
rect 30466 10996 30472 11008
rect 30423 10968 30472 10996
rect 30423 10965 30435 10968
rect 30377 10959 30435 10965
rect 30466 10956 30472 10968
rect 30524 10956 30530 11008
rect 30650 10956 30656 11008
rect 30708 10996 30714 11008
rect 30837 10999 30895 11005
rect 30837 10996 30849 10999
rect 30708 10968 30849 10996
rect 30708 10956 30714 10968
rect 30837 10965 30849 10968
rect 30883 10965 30895 10999
rect 30837 10959 30895 10965
rect 32582 10956 32588 11008
rect 32640 10956 32646 11008
rect 33318 10956 33324 11008
rect 33376 10996 33382 11008
rect 33520 11005 33548 11036
rect 33505 10999 33563 11005
rect 33505 10996 33517 10999
rect 33376 10968 33517 10996
rect 33376 10956 33382 10968
rect 33505 10965 33517 10968
rect 33551 10965 33563 10999
rect 33505 10959 33563 10965
rect 34790 10956 34796 11008
rect 34848 10996 34854 11008
rect 35452 10996 35480 11095
rect 34848 10968 35480 10996
rect 35636 10996 35664 11095
rect 35728 11064 35756 11095
rect 36262 11092 36268 11104
rect 36320 11092 36326 11144
rect 36630 11092 36636 11144
rect 36688 11092 36694 11144
rect 36078 11064 36084 11076
rect 35728 11036 36084 11064
rect 36078 11024 36084 11036
rect 36136 11024 36142 11076
rect 37458 11024 37464 11076
rect 37516 11024 37522 11076
rect 36170 10996 36176 11008
rect 35636 10968 36176 10996
rect 34848 10956 34854 10968
rect 36170 10956 36176 10968
rect 36228 10956 36234 11008
rect 36265 10999 36323 11005
rect 36265 10965 36277 10999
rect 36311 10996 36323 10999
rect 36446 10996 36452 11008
rect 36311 10968 36452 10996
rect 36311 10965 36323 10968
rect 36265 10959 36323 10965
rect 36446 10956 36452 10968
rect 36504 10956 36510 11008
rect 1104 10906 38824 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 38824 10906
rect 1104 10832 38824 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 1596 10724 1624 10755
rect 3694 10752 3700 10804
rect 3752 10792 3758 10804
rect 4433 10795 4491 10801
rect 4433 10792 4445 10795
rect 3752 10764 4445 10792
rect 3752 10752 3758 10764
rect 4433 10761 4445 10764
rect 4479 10761 4491 10795
rect 8478 10792 8484 10804
rect 4433 10755 4491 10761
rect 6840 10764 8484 10792
rect 2777 10727 2835 10733
rect 1596 10696 1900 10724
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 1360 10628 1409 10656
rect 1360 10616 1366 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1872 10665 1900 10696
rect 2777 10693 2789 10727
rect 2823 10724 2835 10727
rect 2866 10724 2872 10736
rect 2823 10696 2872 10724
rect 2823 10693 2835 10696
rect 2777 10687 2835 10693
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 6840 10733 6868 10764
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 10870 10752 10876 10804
rect 10928 10752 10934 10804
rect 13357 10795 13415 10801
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13630 10792 13636 10804
rect 13403 10764 13636 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 14366 10752 14372 10804
rect 14424 10752 14430 10804
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 14918 10792 14924 10804
rect 14875 10764 14924 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 22278 10752 22284 10804
rect 22336 10792 22342 10804
rect 22922 10792 22928 10804
rect 22336 10764 22928 10792
rect 22336 10752 22342 10764
rect 22922 10752 22928 10764
rect 22980 10752 22986 10804
rect 23017 10795 23075 10801
rect 23017 10761 23029 10795
rect 23063 10792 23075 10795
rect 23290 10792 23296 10804
rect 23063 10764 23296 10792
rect 23063 10761 23075 10764
rect 23017 10755 23075 10761
rect 23290 10752 23296 10764
rect 23348 10792 23354 10804
rect 23348 10764 24624 10792
rect 23348 10752 23354 10764
rect 6825 10727 6883 10733
rect 6825 10693 6837 10727
rect 6871 10693 6883 10727
rect 8202 10724 8208 10736
rect 8050 10696 8208 10724
rect 6825 10687 6883 10693
rect 8202 10684 8208 10696
rect 8260 10724 8266 10736
rect 8260 10696 9798 10724
rect 8260 10684 8266 10696
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1636 10628 1685 10656
rect 1636 10616 1642 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 2498 10616 2504 10668
rect 2556 10616 2562 10668
rect 3878 10616 3884 10668
rect 3936 10616 3942 10668
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5350 10656 5356 10668
rect 5123 10628 5356 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8352 10628 8585 10656
rect 8352 10616 8358 10628
rect 8573 10625 8585 10628
rect 8619 10656 8631 10659
rect 8846 10656 8852 10668
rect 8619 10628 8852 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 10888 10656 10916 10752
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 12621 10727 12679 10733
rect 12621 10724 12633 10727
rect 11388 10696 12633 10724
rect 11388 10684 11394 10696
rect 12621 10693 12633 10696
rect 12667 10724 12679 10727
rect 18322 10724 18328 10736
rect 12667 10696 18328 10724
rect 12667 10693 12679 10696
rect 12621 10687 12679 10693
rect 18322 10684 18328 10696
rect 18380 10724 18386 10736
rect 18380 10696 18538 10724
rect 18380 10684 18386 10696
rect 20990 10684 20996 10736
rect 21048 10684 21054 10736
rect 23845 10727 23903 10733
rect 22066 10696 23152 10724
rect 11057 10659 11115 10665
rect 11057 10656 11069 10659
rect 10888 10628 11069 10656
rect 11057 10625 11069 10628
rect 11103 10625 11115 10659
rect 11057 10619 11115 10625
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 13412 10628 13553 10656
rect 13412 10616 13418 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 13814 10616 13820 10668
rect 13872 10616 13878 10668
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14700 10628 14749 10656
rect 14700 10616 14706 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10656 17187 10659
rect 17218 10656 17224 10668
rect 17175 10628 17224 10656
rect 17175 10625 17187 10628
rect 17129 10619 17187 10625
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17773 10659 17831 10665
rect 17773 10656 17785 10659
rect 17644 10628 17785 10656
rect 17644 10616 17650 10628
rect 17773 10625 17785 10628
rect 17819 10625 17831 10659
rect 22066 10656 22094 10696
rect 22664 10665 22692 10696
rect 17773 10619 17831 10625
rect 21468 10628 22094 10656
rect 22189 10659 22247 10665
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 2087 10560 2237 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2225 10557 2237 10560
rect 2271 10588 2283 10591
rect 4154 10588 4160 10600
rect 2271 10560 4160 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4706 10588 4712 10600
rect 4295 10560 4712 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 8404 10452 8432 10551
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8812 10560 9321 10588
rect 8812 10548 8818 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 10962 10588 10968 10600
rect 10827 10560 10968 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 10962 10548 10968 10560
rect 11020 10588 11026 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11020 10560 12081 10588
rect 11020 10548 11026 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15286 10588 15292 10600
rect 15059 10560 15292 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 20714 10588 20720 10600
rect 20027 10560 20720 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 20714 10548 20720 10560
rect 20772 10548 20778 10600
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 11517 10523 11575 10529
rect 11517 10520 11529 10523
rect 10376 10492 11529 10520
rect 10376 10480 10382 10492
rect 11517 10489 11529 10492
rect 11563 10489 11575 10523
rect 11517 10483 11575 10489
rect 21468 10464 21496 10628
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 22204 10520 22232 10619
rect 22922 10616 22928 10668
rect 22980 10616 22986 10668
rect 23124 10665 23152 10696
rect 23845 10693 23857 10727
rect 23891 10724 23903 10727
rect 24118 10724 24124 10736
rect 23891 10696 24124 10724
rect 23891 10693 23903 10696
rect 23845 10687 23903 10693
rect 24118 10684 24124 10696
rect 24176 10684 24182 10736
rect 24596 10733 24624 10764
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 24949 10795 25007 10801
rect 24949 10792 24961 10795
rect 24912 10764 24961 10792
rect 24912 10752 24918 10764
rect 24949 10761 24961 10764
rect 24995 10761 25007 10795
rect 24949 10755 25007 10761
rect 29178 10752 29184 10804
rect 29236 10752 29242 10804
rect 30190 10752 30196 10804
rect 30248 10752 30254 10804
rect 33134 10752 33140 10804
rect 33192 10792 33198 10804
rect 33962 10792 33968 10804
rect 33192 10764 33968 10792
rect 33192 10752 33198 10764
rect 33962 10752 33968 10764
rect 34020 10792 34026 10804
rect 34057 10795 34115 10801
rect 34057 10792 34069 10795
rect 34020 10764 34069 10792
rect 34020 10752 34026 10764
rect 34057 10761 34069 10764
rect 34103 10761 34115 10795
rect 34057 10755 34115 10761
rect 34425 10795 34483 10801
rect 34425 10761 34437 10795
rect 34471 10792 34483 10795
rect 34698 10792 34704 10804
rect 34471 10764 34704 10792
rect 34471 10761 34483 10764
rect 34425 10755 34483 10761
rect 34698 10752 34704 10764
rect 34756 10752 34762 10804
rect 34885 10795 34943 10801
rect 34885 10761 34897 10795
rect 34931 10792 34943 10795
rect 35342 10792 35348 10804
rect 34931 10764 35348 10792
rect 34931 10761 34943 10764
rect 34885 10755 34943 10761
rect 35342 10752 35348 10764
rect 35400 10752 35406 10804
rect 36633 10795 36691 10801
rect 36633 10761 36645 10795
rect 36679 10792 36691 10795
rect 36722 10792 36728 10804
rect 36679 10764 36728 10792
rect 36679 10761 36691 10764
rect 36633 10755 36691 10761
rect 36722 10752 36728 10764
rect 36780 10752 36786 10804
rect 24581 10727 24639 10733
rect 24581 10693 24593 10727
rect 24627 10693 24639 10727
rect 24581 10687 24639 10693
rect 25593 10727 25651 10733
rect 25593 10693 25605 10727
rect 25639 10724 25651 10727
rect 25682 10724 25688 10736
rect 25639 10696 25688 10724
rect 25639 10693 25651 10696
rect 25593 10687 25651 10693
rect 25682 10684 25688 10696
rect 25740 10724 25746 10736
rect 27801 10727 27859 10733
rect 27801 10724 27813 10727
rect 25740 10696 26648 10724
rect 25740 10684 25746 10696
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 23198 10616 23204 10668
rect 23256 10616 23262 10668
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10656 23443 10659
rect 23474 10656 23480 10668
rect 23431 10628 23480 10656
rect 23431 10625 23443 10628
rect 23385 10619 23443 10625
rect 23474 10616 23480 10628
rect 23532 10616 23538 10668
rect 23750 10616 23756 10668
rect 23808 10656 23814 10668
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23808 10628 24225 10656
rect 23808 10616 23814 10628
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 24302 10616 24308 10668
rect 24360 10616 24366 10668
rect 24765 10659 24823 10665
rect 24765 10656 24777 10659
rect 24596 10628 24777 10656
rect 24596 10600 24624 10628
rect 24765 10625 24777 10628
rect 24811 10625 24823 10659
rect 24765 10619 24823 10625
rect 25774 10616 25780 10668
rect 25832 10616 25838 10668
rect 26326 10616 26332 10668
rect 26384 10616 26390 10668
rect 26418 10616 26424 10668
rect 26476 10616 26482 10668
rect 26620 10665 26648 10696
rect 27172 10696 27813 10724
rect 27172 10668 27200 10696
rect 27801 10693 27813 10696
rect 27847 10693 27859 10727
rect 27801 10687 27859 10693
rect 28534 10684 28540 10736
rect 28592 10724 28598 10736
rect 29196 10724 29224 10752
rect 30208 10724 30236 10752
rect 28592 10696 29132 10724
rect 29196 10696 29500 10724
rect 30208 10696 30788 10724
rect 28592 10684 28598 10696
rect 26605 10659 26663 10665
rect 26605 10625 26617 10659
rect 26651 10625 26663 10659
rect 26605 10619 26663 10625
rect 27154 10616 27160 10668
rect 27212 10616 27218 10668
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10625 27675 10659
rect 27617 10619 27675 10625
rect 22462 10548 22468 10600
rect 22520 10548 22526 10600
rect 23293 10591 23351 10597
rect 23293 10557 23305 10591
rect 23339 10557 23351 10591
rect 23293 10551 23351 10557
rect 23937 10591 23995 10597
rect 23937 10557 23949 10591
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 22738 10520 22744 10532
rect 22204 10492 22744 10520
rect 22738 10480 22744 10492
rect 22796 10480 22802 10532
rect 23308 10520 23336 10551
rect 23216 10492 23336 10520
rect 23952 10520 23980 10551
rect 24578 10548 24584 10600
rect 24636 10548 24642 10600
rect 25961 10591 26019 10597
rect 25961 10557 25973 10591
rect 26007 10588 26019 10591
rect 26050 10588 26056 10600
rect 26007 10560 26056 10588
rect 26007 10557 26019 10560
rect 25961 10551 26019 10557
rect 26050 10548 26056 10560
rect 26108 10548 26114 10600
rect 26789 10591 26847 10597
rect 26789 10557 26801 10591
rect 26835 10588 26847 10591
rect 27065 10591 27123 10597
rect 27065 10588 27077 10591
rect 26835 10560 27077 10588
rect 26835 10557 26847 10560
rect 26789 10551 26847 10557
rect 27065 10557 27077 10560
rect 27111 10588 27123 10591
rect 27632 10588 27660 10619
rect 28994 10616 29000 10668
rect 29052 10616 29058 10668
rect 29104 10656 29132 10696
rect 29472 10665 29500 10696
rect 29273 10659 29331 10665
rect 29273 10656 29285 10659
rect 29104 10628 29285 10656
rect 29273 10625 29285 10628
rect 29319 10625 29331 10659
rect 29273 10619 29331 10625
rect 29457 10659 29515 10665
rect 29457 10625 29469 10659
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 30098 10616 30104 10668
rect 30156 10656 30162 10668
rect 30193 10659 30251 10665
rect 30193 10656 30205 10659
rect 30156 10628 30205 10656
rect 30156 10616 30162 10628
rect 30193 10625 30205 10628
rect 30239 10625 30251 10659
rect 30193 10619 30251 10625
rect 30466 10616 30472 10668
rect 30524 10616 30530 10668
rect 30650 10616 30656 10668
rect 30708 10616 30714 10668
rect 30760 10665 30788 10696
rect 32950 10684 32956 10736
rect 33008 10724 33014 10736
rect 33008 10696 33548 10724
rect 33008 10684 33014 10696
rect 30745 10659 30803 10665
rect 30745 10625 30757 10659
rect 30791 10625 30803 10659
rect 30745 10619 30803 10625
rect 30834 10616 30840 10668
rect 30892 10616 30898 10668
rect 31018 10616 31024 10668
rect 31076 10616 31082 10668
rect 32401 10659 32459 10665
rect 32401 10625 32413 10659
rect 32447 10656 32459 10659
rect 33045 10659 33103 10665
rect 32447 10628 32996 10656
rect 32447 10625 32459 10628
rect 32401 10619 32459 10625
rect 27111 10560 27660 10588
rect 28813 10591 28871 10597
rect 27111 10557 27123 10560
rect 27065 10551 27123 10557
rect 28813 10557 28825 10591
rect 28859 10588 28871 10591
rect 29086 10588 29092 10600
rect 28859 10560 29092 10588
rect 28859 10557 28871 10560
rect 28813 10551 28871 10557
rect 29086 10548 29092 10560
rect 29144 10548 29150 10600
rect 29365 10591 29423 10597
rect 29365 10557 29377 10591
rect 29411 10588 29423 10591
rect 30006 10588 30012 10600
rect 29411 10560 30012 10588
rect 29411 10557 29423 10560
rect 29365 10551 29423 10557
rect 30006 10548 30012 10560
rect 30064 10588 30070 10600
rect 30282 10588 30288 10600
rect 30064 10560 30288 10588
rect 30064 10548 30070 10560
rect 30282 10548 30288 10560
rect 30340 10548 30346 10600
rect 30852 10588 30880 10616
rect 31110 10588 31116 10600
rect 30852 10560 31116 10588
rect 31110 10548 31116 10560
rect 31168 10548 31174 10600
rect 32493 10591 32551 10597
rect 32493 10557 32505 10591
rect 32539 10588 32551 10591
rect 32582 10588 32588 10600
rect 32539 10560 32588 10588
rect 32539 10557 32551 10560
rect 32493 10551 32551 10557
rect 32582 10548 32588 10560
rect 32640 10548 32646 10600
rect 32968 10588 32996 10628
rect 33045 10625 33057 10659
rect 33091 10656 33103 10659
rect 33134 10656 33140 10668
rect 33091 10628 33140 10656
rect 33091 10625 33103 10628
rect 33045 10619 33103 10625
rect 33134 10616 33140 10628
rect 33192 10616 33198 10668
rect 33318 10616 33324 10668
rect 33376 10616 33382 10668
rect 33520 10665 33548 10696
rect 33888 10696 34652 10724
rect 33888 10668 33916 10696
rect 33505 10659 33563 10665
rect 33505 10625 33517 10659
rect 33551 10625 33563 10659
rect 33505 10619 33563 10625
rect 33594 10616 33600 10668
rect 33652 10616 33658 10668
rect 33870 10616 33876 10668
rect 33928 10616 33934 10668
rect 34514 10616 34520 10668
rect 34572 10616 34578 10668
rect 34624 10665 34652 10696
rect 36170 10684 36176 10736
rect 36228 10724 36234 10736
rect 36906 10733 36912 10736
rect 36893 10727 36912 10733
rect 36228 10696 36860 10724
rect 36228 10684 36234 10696
rect 34609 10659 34667 10665
rect 34609 10625 34621 10659
rect 34655 10625 34667 10659
rect 34609 10619 34667 10625
rect 34790 10616 34796 10668
rect 34848 10656 34854 10668
rect 36357 10659 36415 10665
rect 36357 10656 36369 10659
rect 34848 10628 36369 10656
rect 34848 10616 34854 10628
rect 36357 10625 36369 10628
rect 36403 10625 36415 10659
rect 36357 10619 36415 10625
rect 36449 10659 36507 10665
rect 36449 10625 36461 10659
rect 36495 10656 36507 10659
rect 36538 10656 36544 10668
rect 36495 10628 36544 10656
rect 36495 10625 36507 10628
rect 36449 10619 36507 10625
rect 36538 10616 36544 10628
rect 36596 10616 36602 10668
rect 36832 10656 36860 10696
rect 36893 10693 36905 10727
rect 36893 10687 36912 10693
rect 36906 10684 36912 10687
rect 36964 10684 36970 10736
rect 37093 10727 37151 10733
rect 37093 10693 37105 10727
rect 37139 10693 37151 10727
rect 37093 10687 37151 10693
rect 37461 10727 37519 10733
rect 37461 10693 37473 10727
rect 37507 10724 37519 10727
rect 37829 10727 37887 10733
rect 37829 10724 37841 10727
rect 37507 10696 37841 10724
rect 37507 10693 37519 10696
rect 37461 10687 37519 10693
rect 37829 10693 37841 10696
rect 37875 10693 37887 10727
rect 37829 10687 37887 10693
rect 36998 10656 37004 10668
rect 36832 10628 37004 10656
rect 36998 10616 37004 10628
rect 37056 10656 37062 10668
rect 37108 10656 37136 10687
rect 37056 10628 37136 10656
rect 37056 10616 37062 10628
rect 37182 10616 37188 10668
rect 37240 10656 37246 10668
rect 37277 10659 37335 10665
rect 37277 10656 37289 10659
rect 37240 10628 37289 10656
rect 37240 10616 37246 10628
rect 37277 10625 37289 10628
rect 37323 10625 37335 10659
rect 37277 10619 37335 10625
rect 37553 10659 37611 10665
rect 37553 10625 37565 10659
rect 37599 10625 37611 10659
rect 37553 10619 37611 10625
rect 33612 10588 33640 10616
rect 34149 10591 34207 10597
rect 34149 10588 34161 10591
rect 32968 10560 34161 10588
rect 34149 10557 34161 10560
rect 34195 10557 34207 10591
rect 34149 10551 34207 10557
rect 36170 10548 36176 10600
rect 36228 10548 36234 10600
rect 36265 10591 36323 10597
rect 36265 10557 36277 10591
rect 36311 10557 36323 10591
rect 36265 10551 36323 10557
rect 24026 10520 24032 10532
rect 23952 10492 24032 10520
rect 8570 10452 8576 10464
rect 8343 10424 8576 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 8757 10455 8815 10461
rect 8757 10452 8769 10455
rect 8720 10424 8769 10452
rect 8720 10412 8726 10424
rect 8757 10421 8769 10424
rect 8803 10421 8815 10455
rect 8757 10415 8815 10421
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11330 10452 11336 10464
rect 11287 10424 11336 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12894 10412 12900 10464
rect 12952 10412 12958 10464
rect 17221 10455 17279 10461
rect 17221 10421 17233 10455
rect 17267 10452 17279 10455
rect 17862 10452 17868 10464
rect 17267 10424 17868 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 18506 10412 18512 10464
rect 18564 10452 18570 10464
rect 19521 10455 19579 10461
rect 19521 10452 19533 10455
rect 18564 10424 19533 10452
rect 18564 10412 18570 10424
rect 19521 10421 19533 10424
rect 19567 10421 19579 10455
rect 19521 10415 19579 10421
rect 21450 10412 21456 10464
rect 21508 10412 21514 10464
rect 21818 10412 21824 10464
rect 21876 10412 21882 10464
rect 22370 10412 22376 10464
rect 22428 10452 22434 10464
rect 23216 10452 23244 10492
rect 24026 10480 24032 10492
rect 24084 10520 24090 10532
rect 26142 10520 26148 10532
rect 24084 10492 26148 10520
rect 24084 10480 24090 10492
rect 26142 10480 26148 10492
rect 26200 10480 26206 10532
rect 27525 10523 27583 10529
rect 27525 10489 27537 10523
rect 27571 10520 27583 10523
rect 27890 10520 27896 10532
rect 27571 10492 27896 10520
rect 27571 10489 27583 10492
rect 27525 10483 27583 10489
rect 27890 10480 27896 10492
rect 27948 10480 27954 10532
rect 32600 10520 32628 10548
rect 33689 10523 33747 10529
rect 33689 10520 33701 10523
rect 32600 10492 33701 10520
rect 33689 10489 33701 10492
rect 33735 10489 33747 10523
rect 33689 10483 33747 10489
rect 36078 10480 36084 10532
rect 36136 10520 36142 10532
rect 36280 10520 36308 10551
rect 36906 10548 36912 10600
rect 36964 10588 36970 10600
rect 37568 10588 37596 10619
rect 36964 10560 37596 10588
rect 36964 10548 36970 10560
rect 38378 10548 38384 10600
rect 38436 10548 38442 10600
rect 36136 10492 36308 10520
rect 36136 10480 36142 10492
rect 22428 10424 23244 10452
rect 24489 10455 24547 10461
rect 22428 10412 22434 10424
rect 24489 10421 24501 10455
rect 24535 10452 24547 10455
rect 24670 10452 24676 10464
rect 24535 10424 24676 10452
rect 24535 10421 24547 10424
rect 24489 10415 24547 10421
rect 24670 10412 24676 10424
rect 24728 10412 24734 10464
rect 27985 10455 28043 10461
rect 27985 10421 27997 10455
rect 28031 10452 28043 10455
rect 28258 10452 28264 10464
rect 28031 10424 28264 10452
rect 28031 10421 28043 10424
rect 27985 10415 28043 10421
rect 28258 10412 28264 10424
rect 28316 10412 28322 10464
rect 30377 10455 30435 10461
rect 30377 10421 30389 10455
rect 30423 10452 30435 10455
rect 30742 10452 30748 10464
rect 30423 10424 30748 10452
rect 30423 10421 30435 10424
rect 30377 10415 30435 10421
rect 30742 10412 30748 10424
rect 30800 10412 30806 10464
rect 31205 10455 31263 10461
rect 31205 10421 31217 10455
rect 31251 10452 31263 10455
rect 32306 10452 32312 10464
rect 31251 10424 32312 10452
rect 31251 10421 31263 10424
rect 31205 10415 31263 10421
rect 32306 10412 32312 10424
rect 32364 10412 32370 10464
rect 32766 10412 32772 10464
rect 32824 10412 32830 10464
rect 32861 10455 32919 10461
rect 32861 10421 32873 10455
rect 32907 10452 32919 10455
rect 32950 10452 32956 10464
rect 32907 10424 32956 10452
rect 32907 10421 32919 10424
rect 32861 10415 32919 10421
rect 32950 10412 32956 10424
rect 33008 10412 33014 10464
rect 33226 10412 33232 10464
rect 33284 10452 33290 10464
rect 34241 10455 34299 10461
rect 34241 10452 34253 10455
rect 33284 10424 34253 10452
rect 33284 10412 33290 10424
rect 34241 10421 34253 10424
rect 34287 10421 34299 10455
rect 34241 10415 34299 10421
rect 34606 10412 34612 10464
rect 34664 10452 34670 10464
rect 35342 10452 35348 10464
rect 34664 10424 35348 10452
rect 34664 10412 34670 10424
rect 35342 10412 35348 10424
rect 35400 10412 35406 10464
rect 36280 10452 36308 10492
rect 36725 10523 36783 10529
rect 36725 10489 36737 10523
rect 36771 10520 36783 10523
rect 37826 10520 37832 10532
rect 36771 10492 37832 10520
rect 36771 10489 36783 10492
rect 36725 10483 36783 10489
rect 37826 10480 37832 10492
rect 37884 10480 37890 10532
rect 36814 10452 36820 10464
rect 36280 10424 36820 10452
rect 36814 10412 36820 10424
rect 36872 10452 36878 10464
rect 36909 10455 36967 10461
rect 36909 10452 36921 10455
rect 36872 10424 36921 10452
rect 36872 10412 36878 10424
rect 36909 10421 36921 10424
rect 36955 10421 36967 10455
rect 36909 10415 36967 10421
rect 37274 10412 37280 10464
rect 37332 10412 37338 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 1673 10251 1731 10257
rect 1673 10248 1685 10251
rect 1360 10220 1685 10248
rect 1360 10208 1366 10220
rect 1673 10217 1685 10220
rect 1719 10217 1731 10251
rect 1673 10211 1731 10217
rect 8113 10251 8171 10257
rect 8113 10217 8125 10251
rect 8159 10248 8171 10251
rect 8386 10248 8392 10260
rect 8159 10220 8392 10248
rect 8159 10217 8171 10220
rect 8113 10211 8171 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8754 10208 8760 10260
rect 8812 10208 8818 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13872 10220 14105 10248
rect 13872 10208 13878 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14829 10251 14887 10257
rect 14829 10248 14841 10251
rect 14516 10220 14841 10248
rect 14516 10208 14522 10220
rect 14829 10217 14841 10220
rect 14875 10217 14887 10251
rect 14829 10211 14887 10217
rect 16945 10251 17003 10257
rect 16945 10217 16957 10251
rect 16991 10248 17003 10251
rect 17589 10251 17647 10257
rect 17589 10248 17601 10251
rect 16991 10220 17601 10248
rect 16991 10217 17003 10220
rect 16945 10211 17003 10217
rect 17589 10217 17601 10220
rect 17635 10248 17647 10251
rect 17954 10248 17960 10260
rect 17635 10220 17960 10248
rect 17635 10217 17647 10220
rect 17589 10211 17647 10217
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18138 10208 18144 10260
rect 18196 10208 18202 10260
rect 20714 10208 20720 10260
rect 20772 10208 20778 10260
rect 23293 10251 23351 10257
rect 23293 10217 23305 10251
rect 23339 10248 23351 10251
rect 23382 10248 23388 10260
rect 23339 10220 23388 10248
rect 23339 10217 23351 10220
rect 23293 10211 23351 10217
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 23658 10208 23664 10260
rect 23716 10208 23722 10260
rect 23934 10248 23940 10260
rect 23768 10220 23940 10248
rect 14918 10140 14924 10192
rect 14976 10180 14982 10192
rect 15105 10183 15163 10189
rect 15105 10180 15117 10183
rect 14976 10152 15117 10180
rect 14976 10140 14982 10152
rect 15105 10149 15117 10152
rect 15151 10149 15163 10183
rect 15105 10143 15163 10149
rect 17126 10140 17132 10192
rect 17184 10180 17190 10192
rect 17681 10183 17739 10189
rect 17681 10180 17693 10183
rect 17184 10152 17693 10180
rect 17184 10140 17190 10152
rect 17681 10149 17693 10152
rect 17727 10149 17739 10183
rect 21818 10180 21824 10192
rect 17681 10143 17739 10149
rect 21192 10152 21824 10180
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 4856 10084 4997 10112
rect 4856 10072 4862 10084
rect 4985 10081 4997 10084
rect 5031 10112 5043 10115
rect 6546 10112 6552 10124
rect 5031 10084 6552 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 8478 10072 8484 10124
rect 8536 10072 8542 10124
rect 8570 10072 8576 10124
rect 8628 10112 8634 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 8628 10084 9505 10112
rect 8628 10072 8634 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 11054 10112 11060 10124
rect 10551 10084 11060 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 11606 10112 11612 10124
rect 11379 10084 11612 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 13170 10112 13176 10124
rect 12676 10084 13176 10112
rect 12676 10072 12682 10084
rect 13170 10072 13176 10084
rect 13228 10112 13234 10124
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13228 10084 13737 10112
rect 13228 10072 13234 10084
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 15197 10115 15255 10121
rect 15197 10081 15209 10115
rect 15243 10112 15255 10115
rect 15378 10112 15384 10124
rect 15243 10084 15384 10112
rect 15243 10081 15255 10084
rect 15197 10075 15255 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 17037 10115 17095 10121
rect 16439 10084 16620 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6748 10016 7389 10044
rect 5258 9936 5264 9988
rect 5316 9936 5322 9988
rect 5368 9948 5750 9976
rect 934 9868 940 9920
rect 992 9908 998 9920
rect 1397 9911 1455 9917
rect 1397 9908 1409 9911
rect 992 9880 1409 9908
rect 992 9868 998 9880
rect 1397 9877 1409 9880
rect 1443 9877 1455 9911
rect 1397 9871 1455 9877
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 5368 9908 5396 9948
rect 6748 9920 6776 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10044 8171 10047
rect 8294 10044 8300 10056
rect 8159 10016 8300 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 7944 9976 7972 10007
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 10318 10044 10324 10056
rect 8435 10016 10324 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 10870 10044 10876 10056
rect 10735 10016 10876 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 12894 10044 12900 10056
rect 12742 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10044 12958 10056
rect 13446 10044 13452 10056
rect 12952 10016 13452 10044
rect 12952 10004 12958 10016
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 14240 10016 14289 10044
rect 14240 10004 14246 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14550 10004 14556 10056
rect 14608 10004 14614 10056
rect 14642 10004 14648 10056
rect 14700 10044 14706 10056
rect 14737 10047 14795 10053
rect 14737 10044 14749 10047
rect 14700 10016 14749 10044
rect 14700 10004 14706 10016
rect 14737 10013 14749 10016
rect 14783 10044 14795 10047
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 14783 10016 15025 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 15286 10004 15292 10056
rect 15344 10004 15350 10056
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 7944 9948 8953 9976
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 11609 9979 11667 9985
rect 11609 9945 11621 9979
rect 11655 9976 11667 9979
rect 11882 9976 11888 9988
rect 11655 9948 11888 9976
rect 11655 9945 11667 9948
rect 11609 9939 11667 9945
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 13633 9979 13691 9985
rect 13633 9976 13645 9979
rect 13096 9948 13645 9976
rect 13096 9920 13124 9948
rect 13633 9945 13645 9948
rect 13679 9976 13691 9979
rect 13998 9976 14004 9988
rect 13679 9948 14004 9976
rect 13679 9945 13691 9948
rect 13633 9939 13691 9945
rect 13998 9936 14004 9948
rect 14056 9936 14062 9988
rect 16316 9976 16344 10007
rect 16482 10004 16488 10056
rect 16540 10004 16546 10056
rect 16592 10044 16620 10084
rect 17037 10081 17049 10115
rect 17083 10112 17095 10115
rect 17218 10112 17224 10124
rect 17083 10084 17224 10112
rect 17083 10081 17095 10084
rect 17037 10075 17095 10081
rect 17218 10072 17224 10084
rect 17276 10112 17282 10124
rect 17770 10112 17776 10124
rect 17276 10084 17776 10112
rect 17276 10072 17282 10084
rect 17328 10053 17356 10084
rect 17770 10072 17776 10084
rect 17828 10112 17834 10124
rect 17828 10084 18552 10112
rect 17828 10072 17834 10084
rect 18524 10056 18552 10084
rect 18690 10072 18696 10124
rect 18748 10072 18754 10124
rect 21192 10121 21220 10152
rect 21818 10140 21824 10152
rect 21876 10140 21882 10192
rect 21910 10140 21916 10192
rect 21968 10180 21974 10192
rect 23768 10180 23796 10220
rect 23934 10208 23940 10220
rect 23992 10208 23998 10260
rect 24026 10208 24032 10260
rect 24084 10208 24090 10260
rect 26329 10251 26387 10257
rect 26329 10217 26341 10251
rect 26375 10248 26387 10251
rect 27154 10248 27160 10260
rect 26375 10220 27160 10248
rect 26375 10217 26387 10220
rect 26329 10211 26387 10217
rect 27154 10208 27160 10220
rect 27212 10208 27218 10260
rect 28077 10251 28135 10257
rect 28077 10217 28089 10251
rect 28123 10248 28135 10251
rect 28534 10248 28540 10260
rect 28123 10220 28540 10248
rect 28123 10217 28135 10220
rect 28077 10211 28135 10217
rect 28534 10208 28540 10220
rect 28592 10208 28598 10260
rect 28813 10251 28871 10257
rect 28813 10217 28825 10251
rect 28859 10248 28871 10251
rect 28994 10248 29000 10260
rect 28859 10220 29000 10248
rect 28859 10217 28871 10220
rect 28813 10211 28871 10217
rect 28994 10208 29000 10220
rect 29052 10208 29058 10260
rect 30098 10208 30104 10260
rect 30156 10208 30162 10260
rect 30745 10251 30803 10257
rect 30745 10217 30757 10251
rect 30791 10248 30803 10251
rect 31018 10248 31024 10260
rect 30791 10220 31024 10248
rect 30791 10217 30803 10220
rect 30745 10211 30803 10217
rect 31018 10208 31024 10220
rect 31076 10208 31082 10260
rect 34333 10251 34391 10257
rect 34333 10217 34345 10251
rect 34379 10217 34391 10251
rect 34333 10211 34391 10217
rect 25225 10183 25283 10189
rect 25225 10180 25237 10183
rect 21968 10152 23244 10180
rect 21968 10140 21974 10152
rect 21177 10115 21235 10121
rect 21177 10081 21189 10115
rect 21223 10081 21235 10115
rect 21177 10075 21235 10081
rect 21358 10072 21364 10124
rect 21416 10112 21422 10124
rect 22097 10115 22155 10121
rect 22097 10112 22109 10115
rect 21416 10084 22109 10112
rect 21416 10072 21422 10084
rect 22097 10081 22109 10084
rect 22143 10081 22155 10115
rect 22097 10075 22155 10081
rect 16761 10047 16819 10053
rect 16592 10038 16712 10044
rect 16761 10038 16773 10047
rect 16592 10016 16773 10038
rect 16684 10013 16773 10016
rect 16807 10013 16819 10047
rect 16684 10010 16819 10013
rect 16761 10007 16819 10010
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17681 10047 17739 10053
rect 17681 10044 17693 10047
rect 17451 10016 17693 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 17681 10013 17693 10016
rect 17727 10013 17739 10047
rect 17681 10007 17739 10013
rect 17420 9976 17448 10007
rect 16316 9948 17448 9976
rect 17589 9979 17647 9985
rect 17589 9945 17601 9979
rect 17635 9945 17647 9979
rect 17696 9976 17724 10007
rect 17862 10004 17868 10056
rect 17920 10004 17926 10056
rect 17954 10004 17960 10056
rect 18012 10004 18018 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10044 21143 10047
rect 21450 10044 21456 10056
rect 21131 10016 21456 10044
rect 21131 10013 21143 10016
rect 21085 10007 21143 10013
rect 21450 10004 21456 10016
rect 21508 10044 21514 10056
rect 22557 10047 22615 10053
rect 21508 10016 22094 10044
rect 21508 10004 21514 10016
rect 18322 9976 18328 9988
rect 17696 9948 18328 9976
rect 17589 9939 17647 9945
rect 3936 9880 5396 9908
rect 3936 9868 3942 9880
rect 6730 9868 6736 9920
rect 6788 9868 6794 9920
rect 6822 9868 6828 9920
rect 6880 9868 6886 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 9732 9880 9873 9908
rect 9732 9868 9738 9880
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 9861 9871 9919 9877
rect 11238 9868 11244 9920
rect 11296 9868 11302 9920
rect 13078 9868 13084 9920
rect 13136 9868 13142 9920
rect 13170 9868 13176 9920
rect 13228 9868 13234 9920
rect 13538 9868 13544 9920
rect 13596 9868 13602 9920
rect 16577 9911 16635 9917
rect 16577 9877 16589 9911
rect 16623 9908 16635 9911
rect 16666 9908 16672 9920
rect 16623 9880 16672 9908
rect 16623 9877 16635 9880
rect 16577 9871 16635 9877
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 16850 9868 16856 9920
rect 16908 9908 16914 9920
rect 17129 9911 17187 9917
rect 17129 9908 17141 9911
rect 16908 9880 17141 9908
rect 16908 9868 16914 9880
rect 17129 9877 17141 9880
rect 17175 9877 17187 9911
rect 17129 9871 17187 9877
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 17604 9908 17632 9939
rect 18322 9936 18328 9948
rect 18380 9976 18386 9988
rect 18601 9979 18659 9985
rect 18601 9976 18613 9979
rect 18380 9948 18613 9976
rect 18380 9936 18386 9948
rect 18601 9945 18613 9948
rect 18647 9976 18659 9979
rect 19242 9976 19248 9988
rect 18647 9948 19248 9976
rect 18647 9945 18659 9948
rect 18601 9939 18659 9945
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 22066 9976 22094 10016
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 22664 10044 22692 10152
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10112 22799 10115
rect 23106 10112 23112 10124
rect 22787 10084 23112 10112
rect 22787 10081 22799 10084
rect 22741 10075 22799 10081
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 23216 10112 23244 10152
rect 23676 10152 23796 10180
rect 24780 10152 25237 10180
rect 23676 10112 23704 10152
rect 24780 10124 24808 10152
rect 25225 10149 25237 10152
rect 25271 10149 25283 10183
rect 25225 10143 25283 10149
rect 27798 10140 27804 10192
rect 27856 10180 27862 10192
rect 27893 10183 27951 10189
rect 27893 10180 27905 10183
rect 27856 10152 27905 10180
rect 27856 10140 27862 10152
rect 27893 10149 27905 10152
rect 27939 10149 27951 10183
rect 27893 10143 27951 10149
rect 28629 10183 28687 10189
rect 28629 10149 28641 10183
rect 28675 10180 28687 10183
rect 29086 10180 29092 10192
rect 28675 10152 29092 10180
rect 28675 10149 28687 10152
rect 28629 10143 28687 10149
rect 29086 10140 29092 10152
rect 29144 10140 29150 10192
rect 23216 10084 23704 10112
rect 22603 10016 22692 10044
rect 22925 10047 22983 10053
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 22925 10013 22937 10047
rect 22971 10044 22983 10047
rect 23198 10044 23204 10056
rect 22971 10016 23204 10044
rect 22971 10013 22983 10016
rect 22925 10007 22983 10013
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 23290 10004 23296 10056
rect 23348 10004 23354 10056
rect 23584 10053 23612 10084
rect 24670 10072 24676 10124
rect 24728 10072 24734 10124
rect 24762 10072 24768 10124
rect 24820 10072 24826 10124
rect 25682 10072 25688 10124
rect 25740 10072 25746 10124
rect 26142 10072 26148 10124
rect 26200 10072 26206 10124
rect 29638 10072 29644 10124
rect 29696 10072 29702 10124
rect 23385 10047 23443 10053
rect 23385 10013 23397 10047
rect 23431 10013 23443 10047
rect 23385 10007 23443 10013
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 22373 9979 22431 9985
rect 22373 9976 22385 9979
rect 22066 9948 22385 9976
rect 22373 9945 22385 9948
rect 22419 9945 22431 9979
rect 23400 9976 23428 10007
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 23839 10047 23897 10053
rect 23839 10022 23851 10047
rect 23885 10022 23897 10047
rect 23937 10047 23995 10053
rect 23839 10007 23848 10022
rect 22373 9939 22431 9945
rect 22664 9948 23428 9976
rect 23842 9970 23848 10007
rect 23900 9970 23906 10022
rect 23937 10013 23949 10047
rect 23983 10038 23995 10047
rect 23983 10013 24072 10038
rect 23937 10010 24072 10013
rect 23937 10007 23995 10010
rect 24044 9976 24072 10010
rect 24118 10004 24124 10056
rect 24176 10004 24182 10056
rect 24394 10004 24400 10056
rect 24452 10004 24458 10056
rect 24486 10004 24492 10056
rect 24544 10044 24550 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24544 10016 24593 10044
rect 24544 10004 24550 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10044 25007 10047
rect 25130 10044 25136 10056
rect 24995 10016 25136 10044
rect 24995 10013 25007 10016
rect 24949 10007 25007 10013
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25593 10047 25651 10053
rect 25593 10013 25605 10047
rect 25639 10044 25651 10047
rect 25639 10016 25912 10044
rect 25639 10013 25651 10016
rect 25593 10007 25651 10013
rect 25774 9976 25780 9988
rect 24044 9948 25780 9976
rect 17368 9880 17632 9908
rect 17368 9868 17374 9880
rect 21542 9868 21548 9920
rect 21600 9868 21606 9920
rect 21910 9868 21916 9920
rect 21968 9868 21974 9920
rect 22005 9911 22063 9917
rect 22005 9877 22017 9911
rect 22051 9908 22063 9911
rect 22186 9908 22192 9920
rect 22051 9880 22192 9908
rect 22051 9877 22063 9880
rect 22005 9871 22063 9877
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 22388 9908 22416 9939
rect 22664 9908 22692 9948
rect 22388 9880 22692 9908
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 23017 9911 23075 9917
rect 23017 9908 23029 9911
rect 22980 9880 23029 9908
rect 22980 9868 22986 9880
rect 23017 9877 23029 9880
rect 23063 9908 23075 9911
rect 23569 9911 23627 9917
rect 23569 9908 23581 9911
rect 23063 9880 23581 9908
rect 23063 9877 23075 9880
rect 23017 9871 23075 9877
rect 23569 9877 23581 9880
rect 23615 9908 23627 9911
rect 24044 9908 24072 9948
rect 25774 9936 25780 9948
rect 25832 9936 25838 9988
rect 25884 9976 25912 10016
rect 25958 10004 25964 10056
rect 26016 10044 26022 10056
rect 26053 10047 26111 10053
rect 26053 10044 26065 10047
rect 26016 10016 26065 10044
rect 26016 10004 26022 10016
rect 26053 10013 26065 10016
rect 26099 10013 26111 10047
rect 26053 10007 26111 10013
rect 28258 10004 28264 10056
rect 28316 10044 28322 10056
rect 28721 10047 28779 10053
rect 28721 10044 28733 10047
rect 28316 10016 28733 10044
rect 28316 10004 28322 10016
rect 28721 10013 28733 10016
rect 28767 10013 28779 10047
rect 28721 10007 28779 10013
rect 28905 10047 28963 10053
rect 28905 10013 28917 10047
rect 28951 10013 28963 10047
rect 28905 10007 28963 10013
rect 27430 9976 27436 9988
rect 25884 9948 27436 9976
rect 27430 9936 27436 9948
rect 27488 9976 27494 9988
rect 27617 9979 27675 9985
rect 27617 9976 27629 9979
rect 27488 9948 27629 9976
rect 27488 9936 27494 9948
rect 27617 9945 27629 9948
rect 27663 9945 27675 9979
rect 27617 9939 27675 9945
rect 28442 9936 28448 9988
rect 28500 9976 28506 9988
rect 28920 9976 28948 10007
rect 29730 10004 29736 10056
rect 29788 10004 29794 10056
rect 30116 10044 30144 10208
rect 30282 10140 30288 10192
rect 30340 10180 30346 10192
rect 30340 10152 30512 10180
rect 30340 10140 30346 10152
rect 30484 10053 30512 10152
rect 30285 10047 30343 10053
rect 30285 10044 30297 10047
rect 30116 10016 30297 10044
rect 30285 10013 30297 10016
rect 30331 10013 30343 10047
rect 30285 10007 30343 10013
rect 30469 10047 30527 10053
rect 30469 10013 30481 10047
rect 30515 10013 30527 10047
rect 30469 10007 30527 10013
rect 30742 10004 30748 10056
rect 30800 10004 30806 10056
rect 30923 10047 30981 10053
rect 30923 10044 30935 10047
rect 30852 10016 30935 10044
rect 28500 9948 28948 9976
rect 30377 9979 30435 9985
rect 28500 9936 28506 9948
rect 30377 9945 30389 9979
rect 30423 9976 30435 9979
rect 30852 9976 30880 10016
rect 30923 10013 30935 10016
rect 30969 10013 30981 10047
rect 30923 10007 30981 10013
rect 30423 9948 30880 9976
rect 31036 9976 31064 10208
rect 31757 10183 31815 10189
rect 31757 10149 31769 10183
rect 31803 10180 31815 10183
rect 32398 10180 32404 10192
rect 31803 10152 32404 10180
rect 31803 10149 31815 10152
rect 31757 10143 31815 10149
rect 32398 10140 32404 10152
rect 32456 10140 32462 10192
rect 34348 10180 34376 10211
rect 34514 10208 34520 10260
rect 34572 10248 34578 10260
rect 34974 10248 34980 10260
rect 34572 10220 34980 10248
rect 34572 10208 34578 10220
rect 34974 10208 34980 10220
rect 35032 10248 35038 10260
rect 36449 10251 36507 10257
rect 36449 10248 36461 10251
rect 35032 10220 36461 10248
rect 35032 10208 35038 10220
rect 36449 10217 36461 10220
rect 36495 10217 36507 10251
rect 36449 10211 36507 10217
rect 34606 10180 34612 10192
rect 34348 10152 34612 10180
rect 34606 10140 34612 10152
rect 34664 10140 34670 10192
rect 31110 10072 31116 10124
rect 31168 10072 31174 10124
rect 34701 10115 34759 10121
rect 31588 10084 32168 10112
rect 31588 10056 31616 10084
rect 31570 10004 31576 10056
rect 31628 10004 31634 10056
rect 32140 10053 32168 10084
rect 34701 10081 34713 10115
rect 34747 10112 34759 10115
rect 36909 10115 36967 10121
rect 34747 10084 36676 10112
rect 34747 10081 34759 10084
rect 34701 10075 34759 10081
rect 36648 10056 36676 10084
rect 36909 10081 36921 10115
rect 36955 10112 36967 10115
rect 37274 10112 37280 10124
rect 36955 10084 37280 10112
rect 36955 10081 36967 10084
rect 36909 10075 36967 10081
rect 37274 10072 37280 10084
rect 37332 10072 37338 10124
rect 31849 10047 31907 10053
rect 31849 10044 31861 10047
rect 31726 10016 31861 10044
rect 31251 9979 31309 9985
rect 31251 9976 31263 9979
rect 31036 9948 31263 9976
rect 30423 9945 30435 9948
rect 30377 9939 30435 9945
rect 23615 9880 24072 9908
rect 23615 9877 23627 9880
rect 23569 9871 23627 9877
rect 25130 9868 25136 9920
rect 25188 9868 25194 9920
rect 30852 9908 30880 9948
rect 31251 9945 31263 9948
rect 31297 9945 31309 9979
rect 31251 9939 31309 9945
rect 31389 9979 31447 9985
rect 31389 9945 31401 9979
rect 31435 9945 31447 9979
rect 31389 9939 31447 9945
rect 30926 9908 30932 9920
rect 30852 9880 30932 9908
rect 30926 9868 30932 9880
rect 30984 9868 30990 9920
rect 31404 9908 31432 9939
rect 31478 9936 31484 9988
rect 31536 9976 31542 9988
rect 31726 9976 31754 10016
rect 31849 10013 31861 10016
rect 31895 10013 31907 10047
rect 31849 10007 31907 10013
rect 32125 10047 32183 10053
rect 32125 10013 32137 10047
rect 32171 10013 32183 10047
rect 32125 10007 32183 10013
rect 33965 10047 34023 10053
rect 33965 10013 33977 10047
rect 34011 10044 34023 10047
rect 34606 10044 34612 10056
rect 34011 10016 34612 10044
rect 34011 10013 34023 10016
rect 33965 10007 34023 10013
rect 34606 10004 34612 10016
rect 34664 10004 34670 10056
rect 36630 10004 36636 10056
rect 36688 10004 36694 10056
rect 31536 9948 31754 9976
rect 34977 9979 35035 9985
rect 31536 9936 31542 9948
rect 34977 9945 34989 9979
rect 35023 9945 35035 9979
rect 35434 9976 35440 9988
rect 34977 9939 35035 9945
rect 35360 9948 35440 9976
rect 31662 9908 31668 9920
rect 31404 9880 31668 9908
rect 31662 9868 31668 9880
rect 31720 9908 31726 9920
rect 31941 9911 31999 9917
rect 31941 9908 31953 9911
rect 31720 9880 31953 9908
rect 31720 9868 31726 9880
rect 31941 9877 31953 9880
rect 31987 9877 31999 9911
rect 31941 9871 31999 9877
rect 32122 9868 32128 9920
rect 32180 9908 32186 9920
rect 32309 9911 32367 9917
rect 32309 9908 32321 9911
rect 32180 9880 32321 9908
rect 32180 9868 32186 9880
rect 32309 9877 32321 9880
rect 32355 9877 32367 9911
rect 32309 9871 32367 9877
rect 34330 9868 34336 9920
rect 34388 9868 34394 9920
rect 34517 9911 34575 9917
rect 34517 9877 34529 9911
rect 34563 9908 34575 9911
rect 34992 9908 35020 9939
rect 34563 9880 35020 9908
rect 35360 9908 35388 9948
rect 35434 9936 35440 9948
rect 35492 9936 35498 9988
rect 37366 9976 37372 9988
rect 36280 9948 37372 9976
rect 36280 9908 36308 9948
rect 37366 9936 37372 9948
rect 37424 9936 37430 9988
rect 35360 9880 36308 9908
rect 34563 9877 34575 9880
rect 34517 9871 34575 9877
rect 36814 9868 36820 9920
rect 36872 9908 36878 9920
rect 38378 9908 38384 9920
rect 36872 9880 38384 9908
rect 36872 9868 36878 9880
rect 38378 9868 38384 9880
rect 38436 9868 38442 9920
rect 1104 9818 38824 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 38824 9818
rect 1104 9744 38824 9766
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11057 9707 11115 9713
rect 11057 9704 11069 9707
rect 11020 9676 11069 9704
rect 11020 9664 11026 9676
rect 11057 9673 11069 9676
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 11977 9707 12035 9713
rect 11977 9704 11989 9707
rect 11940 9676 11989 9704
rect 11940 9664 11946 9676
rect 11977 9673 11989 9676
rect 12023 9673 12035 9707
rect 11977 9667 12035 9673
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 13354 9704 13360 9716
rect 12483 9676 13360 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 13633 9707 13691 9713
rect 13633 9704 13645 9707
rect 13596 9676 13645 9704
rect 13596 9664 13602 9676
rect 13633 9673 13645 9676
rect 13679 9673 13691 9707
rect 13633 9667 13691 9673
rect 7561 9639 7619 9645
rect 7561 9605 7573 9639
rect 7607 9636 7619 9639
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7607 9608 7849 9636
rect 7607 9605 7619 9608
rect 7561 9599 7619 9605
rect 7837 9605 7849 9608
rect 7883 9605 7895 9639
rect 7837 9599 7895 9605
rect 9858 9596 9864 9648
rect 9916 9596 9922 9648
rect 11238 9596 11244 9648
rect 11296 9596 11302 9648
rect 12345 9639 12403 9645
rect 12345 9605 12357 9639
rect 12391 9636 12403 9639
rect 13078 9636 13084 9648
rect 12391 9608 13084 9636
rect 12391 9605 12403 9608
rect 12345 9599 12403 9605
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 13648 9636 13676 9667
rect 15378 9664 15384 9716
rect 15436 9664 15442 9716
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 17310 9704 17316 9716
rect 16540 9676 17316 9704
rect 16540 9664 16546 9676
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 18230 9664 18236 9716
rect 18288 9664 18294 9716
rect 23014 9664 23020 9716
rect 23072 9704 23078 9716
rect 23474 9704 23480 9716
rect 23072 9676 23480 9704
rect 23072 9664 23078 9676
rect 23474 9664 23480 9676
rect 23532 9704 23538 9716
rect 23658 9704 23664 9716
rect 23532 9676 23664 9704
rect 23532 9664 23538 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 23845 9707 23903 9713
rect 23845 9673 23857 9707
rect 23891 9704 23903 9707
rect 24394 9704 24400 9716
rect 23891 9676 24400 9704
rect 23891 9673 23903 9676
rect 23845 9667 23903 9673
rect 24394 9664 24400 9676
rect 24452 9664 24458 9716
rect 25958 9704 25964 9716
rect 25056 9676 25964 9704
rect 14001 9639 14059 9645
rect 14001 9636 14013 9639
rect 13648 9608 14013 9636
rect 14001 9605 14013 9608
rect 14047 9605 14059 9639
rect 14001 9599 14059 9605
rect 14274 9596 14280 9648
rect 14332 9636 14338 9648
rect 14642 9636 14648 9648
rect 14332 9608 14648 9636
rect 14332 9596 14338 9608
rect 14642 9596 14648 9608
rect 14700 9636 14706 9648
rect 16666 9636 16672 9648
rect 14700 9608 15056 9636
rect 14700 9596 14706 9608
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 6822 9568 6828 9580
rect 4939 9540 6828 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7248 9540 7389 9568
rect 7248 9528 7254 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 8478 9568 8484 9580
rect 7699 9540 8484 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 10686 9528 10692 9580
rect 10744 9568 10750 9580
rect 15028 9577 15056 9608
rect 15764 9608 16672 9636
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10744 9540 10977 9568
rect 10744 9528 10750 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 14737 9571 14795 9577
rect 14737 9568 14749 9571
rect 13587 9540 13952 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 4798 9460 4804 9512
rect 4856 9460 4862 9512
rect 5258 9460 5264 9512
rect 5316 9460 5322 9512
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8168 9472 8401 9500
rect 8168 9460 8174 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6696 9336 7205 9364
rect 6696 9324 6702 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 9140 9364 9168 9463
rect 9398 9460 9404 9512
rect 9456 9460 9462 9512
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 12676 9472 13737 9500
rect 12676 9460 12682 9472
rect 13725 9469 13737 9472
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11241 9435 11299 9441
rect 11241 9432 11253 9435
rect 11112 9404 11253 9432
rect 11112 9392 11118 9404
rect 11241 9401 11253 9404
rect 11287 9401 11299 9435
rect 13924 9432 13952 9540
rect 14016 9540 14749 9568
rect 14016 9512 14044 9540
rect 14737 9537 14749 9540
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 15654 9568 15660 9580
rect 15611 9540 15660 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 15764 9577 15792 9608
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 18248 9636 18276 9664
rect 20990 9636 20996 9648
rect 18248 9608 18354 9636
rect 20838 9608 20996 9636
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 21269 9639 21327 9645
rect 21269 9605 21281 9639
rect 21315 9636 21327 9639
rect 21910 9636 21916 9648
rect 21315 9608 21916 9636
rect 21315 9605 21327 9608
rect 21269 9599 21327 9605
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 22186 9596 22192 9648
rect 22244 9596 22250 9648
rect 23934 9636 23940 9648
rect 22480 9608 22876 9636
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 13998 9460 14004 9512
rect 14056 9460 14062 9512
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14240 9472 14565 9500
rect 14240 9460 14246 9472
rect 14553 9469 14565 9472
rect 14599 9500 14611 9503
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14599 9472 14841 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 14918 9460 14924 9512
rect 14976 9500 14982 9512
rect 15856 9500 15884 9531
rect 14976 9472 15884 9500
rect 16040 9500 16068 9531
rect 16390 9528 16396 9580
rect 16448 9528 16454 9580
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16540 9540 16865 9568
rect 16540 9528 16546 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 17310 9528 17316 9580
rect 17368 9528 17374 9580
rect 17586 9528 17592 9580
rect 17644 9528 17650 9580
rect 22370 9528 22376 9580
rect 22428 9528 22434 9580
rect 22480 9577 22508 9608
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9537 22523 9571
rect 22741 9571 22799 9577
rect 22741 9566 22753 9571
rect 22465 9531 22523 9537
rect 22738 9537 22753 9566
rect 22787 9537 22799 9571
rect 22738 9531 22799 9537
rect 16117 9503 16175 9509
rect 16117 9500 16129 9503
rect 16040 9472 16129 9500
rect 14976 9460 14982 9472
rect 16117 9469 16129 9472
rect 16163 9500 16175 9503
rect 16942 9500 16948 9512
rect 16163 9472 16948 9500
rect 16163 9469 16175 9472
rect 16117 9463 16175 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17865 9503 17923 9509
rect 17865 9469 17877 9503
rect 17911 9500 17923 9503
rect 17954 9500 17960 9512
rect 17911 9472 17960 9500
rect 17911 9469 17923 9472
rect 17865 9463 17923 9469
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 18892 9472 19441 9500
rect 14274 9432 14280 9444
rect 13924 9404 14280 9432
rect 11241 9395 11299 9401
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 15194 9392 15200 9444
rect 15252 9392 15258 9444
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9432 15715 9435
rect 16390 9432 16396 9444
rect 15703 9404 16396 9432
rect 15703 9401 15715 9404
rect 15657 9395 15715 9401
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 10502 9364 10508 9376
rect 9140 9336 10508 9364
rect 7193 9327 7251 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10870 9324 10876 9376
rect 10928 9324 10934 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 12860 9336 13185 9364
rect 12860 9324 12866 9336
rect 13173 9333 13185 9336
rect 13219 9333 13231 9367
rect 13173 9327 13231 9333
rect 15010 9324 15016 9376
rect 15068 9324 15074 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 15344 9336 16221 9364
rect 15344 9324 15350 9336
rect 16209 9333 16221 9336
rect 16255 9333 16267 9367
rect 16209 9327 16267 9333
rect 16301 9367 16359 9373
rect 16301 9333 16313 9367
rect 16347 9364 16359 9367
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 16347 9336 16681 9364
rect 16347 9333 16359 9336
rect 16301 9327 16359 9333
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 16669 9327 16727 9333
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 18892 9364 18920 9472
rect 19429 9469 19441 9472
rect 19475 9500 19487 9503
rect 19702 9500 19708 9512
rect 19475 9472 19708 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 19702 9460 19708 9472
rect 19760 9460 19766 9512
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9500 19855 9503
rect 21542 9500 21548 9512
rect 19843 9472 21548 9500
rect 19843 9469 19855 9472
rect 19797 9463 19855 9469
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 19337 9435 19395 9441
rect 19337 9432 19349 9435
rect 19300 9404 19349 9432
rect 19300 9392 19306 9404
rect 19337 9401 19349 9404
rect 19383 9401 19395 9435
rect 22738 9432 22766 9531
rect 22848 9509 22876 9608
rect 23584 9608 23940 9636
rect 22922 9528 22928 9580
rect 22980 9568 22986 9580
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 22980 9540 23121 9568
rect 22980 9528 22986 9540
rect 23109 9537 23121 9540
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 23198 9528 23204 9580
rect 23256 9528 23262 9580
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9568 23351 9571
rect 23584 9568 23612 9608
rect 23934 9596 23940 9608
rect 23992 9596 23998 9648
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 25056 9636 25084 9676
rect 25958 9664 25964 9676
rect 26016 9664 26022 9716
rect 28169 9707 28227 9713
rect 28169 9673 28181 9707
rect 28215 9704 28227 9707
rect 28442 9704 28448 9716
rect 28215 9676 28448 9704
rect 28215 9673 28227 9676
rect 28169 9667 28227 9673
rect 28442 9664 28448 9676
rect 28500 9664 28506 9716
rect 29457 9707 29515 9713
rect 29457 9673 29469 9707
rect 29503 9704 29515 9707
rect 29638 9704 29644 9716
rect 29503 9676 29644 9704
rect 29503 9673 29515 9676
rect 29457 9667 29515 9673
rect 29638 9664 29644 9676
rect 29696 9664 29702 9716
rect 31297 9707 31355 9713
rect 31297 9673 31309 9707
rect 31343 9704 31355 9707
rect 31478 9704 31484 9716
rect 31343 9676 31484 9704
rect 31343 9673 31355 9676
rect 31297 9667 31355 9673
rect 31478 9664 31484 9676
rect 31536 9664 31542 9716
rect 31662 9664 31668 9716
rect 31720 9664 31726 9716
rect 34330 9664 34336 9716
rect 34388 9704 34394 9716
rect 34425 9707 34483 9713
rect 34425 9704 34437 9707
rect 34388 9676 34437 9704
rect 34388 9664 34394 9676
rect 34425 9673 34437 9676
rect 34471 9673 34483 9707
rect 34425 9667 34483 9673
rect 34606 9664 34612 9716
rect 34664 9704 34670 9716
rect 36265 9707 36323 9713
rect 36265 9704 36277 9707
rect 34664 9676 36277 9704
rect 34664 9664 34670 9676
rect 36265 9673 36277 9676
rect 36311 9704 36323 9707
rect 36906 9704 36912 9716
rect 36311 9676 36912 9704
rect 36311 9673 36323 9676
rect 36265 9667 36323 9673
rect 36906 9664 36912 9676
rect 36964 9664 36970 9716
rect 24912 9608 25084 9636
rect 24912 9596 24918 9608
rect 23339 9540 23612 9568
rect 23339 9537 23351 9540
rect 23293 9531 23351 9537
rect 23658 9528 23664 9580
rect 23716 9528 23722 9580
rect 23845 9571 23903 9577
rect 23845 9537 23857 9571
rect 23891 9568 23903 9571
rect 24946 9568 24952 9580
rect 23891 9540 24952 9568
rect 23891 9537 23903 9540
rect 23845 9531 23903 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 25056 9577 25084 9608
rect 25682 9596 25688 9648
rect 25740 9596 25746 9648
rect 25869 9639 25927 9645
rect 25869 9605 25881 9639
rect 25915 9636 25927 9639
rect 26053 9639 26111 9645
rect 26053 9636 26065 9639
rect 25915 9608 26065 9636
rect 25915 9605 25927 9608
rect 25869 9599 25927 9605
rect 26053 9605 26065 9608
rect 26099 9636 26111 9639
rect 27798 9636 27804 9648
rect 26099 9608 27804 9636
rect 26099 9605 26111 9608
rect 26053 9599 26111 9605
rect 27798 9596 27804 9608
rect 27856 9596 27862 9648
rect 29288 9608 29592 9636
rect 25041 9571 25099 9577
rect 25041 9537 25053 9571
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 25961 9571 26019 9577
rect 25961 9568 25973 9571
rect 25832 9540 25973 9568
rect 25832 9528 25838 9540
rect 25961 9537 25973 9540
rect 26007 9537 26019 9571
rect 25961 9531 26019 9537
rect 26145 9571 26203 9577
rect 26145 9537 26157 9571
rect 26191 9568 26203 9571
rect 26234 9568 26240 9580
rect 26191 9540 26240 9568
rect 26191 9537 26203 9540
rect 26145 9531 26203 9537
rect 22833 9503 22891 9509
rect 22833 9469 22845 9503
rect 22879 9469 22891 9503
rect 22833 9463 22891 9469
rect 23014 9460 23020 9512
rect 23072 9460 23078 9512
rect 23676 9500 23704 9528
rect 25501 9503 25559 9509
rect 25501 9500 25513 9503
rect 23676 9472 25513 9500
rect 25501 9469 25513 9472
rect 25547 9469 25559 9503
rect 25501 9463 25559 9469
rect 26050 9460 26056 9512
rect 26108 9500 26114 9512
rect 26160 9500 26188 9531
rect 26234 9528 26240 9540
rect 26292 9528 26298 9580
rect 28077 9571 28135 9577
rect 28077 9537 28089 9571
rect 28123 9568 28135 9571
rect 28166 9568 28172 9580
rect 28123 9540 28172 9568
rect 28123 9537 28135 9540
rect 28077 9531 28135 9537
rect 28166 9528 28172 9540
rect 28224 9528 28230 9580
rect 28261 9571 28319 9577
rect 28261 9537 28273 9571
rect 28307 9568 28319 9571
rect 28350 9568 28356 9580
rect 28307 9540 28356 9568
rect 28307 9537 28319 9540
rect 28261 9531 28319 9537
rect 28350 9528 28356 9540
rect 28408 9528 28414 9580
rect 29086 9528 29092 9580
rect 29144 9568 29150 9580
rect 29288 9577 29316 9608
rect 29564 9577 29592 9608
rect 31018 9596 31024 9648
rect 31076 9636 31082 9648
rect 32861 9639 32919 9645
rect 31076 9608 31432 9636
rect 31076 9596 31082 9608
rect 29273 9571 29331 9577
rect 29273 9568 29285 9571
rect 29144 9540 29285 9568
rect 29144 9528 29150 9540
rect 29273 9537 29285 9540
rect 29319 9537 29331 9571
rect 29273 9531 29331 9537
rect 29457 9571 29515 9577
rect 29457 9537 29469 9571
rect 29503 9537 29515 9571
rect 29457 9531 29515 9537
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9537 29607 9571
rect 29549 9531 29607 9537
rect 26108 9472 26188 9500
rect 28184 9500 28212 9528
rect 29472 9500 29500 9531
rect 29730 9528 29736 9580
rect 29788 9528 29794 9580
rect 31404 9577 31432 9608
rect 32861 9605 32873 9639
rect 32907 9636 32919 9639
rect 32907 9608 33272 9636
rect 32907 9605 32919 9608
rect 32861 9599 32919 9605
rect 30929 9571 30987 9577
rect 30929 9537 30941 9571
rect 30975 9537 30987 9571
rect 30929 9531 30987 9537
rect 31389 9571 31447 9577
rect 31389 9537 31401 9571
rect 31435 9537 31447 9571
rect 31389 9531 31447 9537
rect 28184 9472 29500 9500
rect 29641 9503 29699 9509
rect 26108 9460 26114 9472
rect 29641 9469 29653 9503
rect 29687 9500 29699 9503
rect 30944 9500 30972 9531
rect 32122 9528 32128 9580
rect 32180 9528 32186 9580
rect 32306 9528 32312 9580
rect 32364 9528 32370 9580
rect 32398 9528 32404 9580
rect 32456 9528 32462 9580
rect 32674 9528 32680 9580
rect 32732 9528 32738 9580
rect 32766 9528 32772 9580
rect 32824 9568 32830 9580
rect 33244 9577 33272 9608
rect 34716 9608 35280 9636
rect 34716 9577 34744 9608
rect 35207 9605 35280 9608
rect 32953 9571 33011 9577
rect 32953 9568 32965 9571
rect 32824 9540 32965 9568
rect 32824 9528 32830 9540
rect 32953 9537 32965 9540
rect 32999 9537 33011 9571
rect 32953 9531 33011 9537
rect 33045 9571 33103 9577
rect 33045 9537 33057 9571
rect 33091 9537 33103 9571
rect 33045 9531 33103 9537
rect 33229 9571 33287 9577
rect 33229 9537 33241 9571
rect 33275 9537 33287 9571
rect 33229 9531 33287 9537
rect 34701 9571 34759 9577
rect 34701 9537 34713 9571
rect 34747 9537 34759 9571
rect 34701 9531 34759 9537
rect 34885 9571 34943 9577
rect 34885 9537 34897 9571
rect 34931 9568 34943 9571
rect 34974 9568 34980 9580
rect 34931 9540 34980 9568
rect 34931 9537 34943 9540
rect 34885 9531 34943 9537
rect 29687 9472 30972 9500
rect 29687 9469 29699 9472
rect 29641 9463 29699 9469
rect 24026 9432 24032 9444
rect 22738 9404 24032 9432
rect 19337 9395 19395 9401
rect 24026 9392 24032 9404
rect 24084 9392 24090 9444
rect 30944 9432 30972 9472
rect 31018 9460 31024 9512
rect 31076 9500 31082 9512
rect 31665 9503 31723 9509
rect 31665 9500 31677 9503
rect 31076 9472 31677 9500
rect 31076 9460 31082 9472
rect 31665 9469 31677 9472
rect 31711 9469 31723 9503
rect 31665 9463 31723 9469
rect 32493 9503 32551 9509
rect 32493 9469 32505 9503
rect 32539 9500 32551 9503
rect 32784 9500 32812 9528
rect 33060 9500 33088 9531
rect 34974 9528 34980 9540
rect 35032 9528 35038 9580
rect 35207 9571 35219 9605
rect 35253 9571 35280 9605
rect 35434 9596 35440 9648
rect 35492 9636 35498 9648
rect 35897 9639 35955 9645
rect 35897 9636 35909 9639
rect 35492 9608 35909 9636
rect 35492 9596 35498 9608
rect 35897 9605 35909 9608
rect 35943 9605 35955 9639
rect 35897 9599 35955 9605
rect 36113 9639 36171 9645
rect 36113 9605 36125 9639
rect 36159 9636 36171 9639
rect 36357 9639 36415 9645
rect 36357 9636 36369 9639
rect 36159 9608 36369 9636
rect 36159 9605 36171 9608
rect 36113 9599 36171 9605
rect 36357 9605 36369 9608
rect 36403 9636 36415 9639
rect 37093 9639 37151 9645
rect 36403 9608 37044 9636
rect 36403 9605 36415 9608
rect 36357 9599 36415 9605
rect 35207 9568 35280 9571
rect 35526 9568 35532 9580
rect 35207 9565 35532 9568
rect 35252 9540 35532 9565
rect 35526 9528 35532 9540
rect 35584 9568 35590 9580
rect 35584 9540 35940 9568
rect 35584 9528 35590 9540
rect 32539 9472 32812 9500
rect 32968 9472 33088 9500
rect 32539 9469 32551 9472
rect 32493 9463 32551 9469
rect 31481 9435 31539 9441
rect 31481 9432 31493 9435
rect 30944 9404 31493 9432
rect 31481 9401 31493 9404
rect 31527 9401 31539 9435
rect 31481 9395 31539 9401
rect 32674 9392 32680 9444
rect 32732 9432 32738 9444
rect 32968 9432 32996 9472
rect 34422 9460 34428 9512
rect 34480 9500 34486 9512
rect 34606 9500 34612 9512
rect 34480 9472 34612 9500
rect 34480 9460 34486 9472
rect 34606 9460 34612 9472
rect 34664 9460 34670 9512
rect 34793 9503 34851 9509
rect 34793 9469 34805 9503
rect 34839 9500 34851 9503
rect 35434 9500 35440 9512
rect 34839 9472 35440 9500
rect 34839 9469 34851 9472
rect 34793 9463 34851 9469
rect 32732 9404 32996 9432
rect 32732 9392 32738 9404
rect 17644 9336 18920 9364
rect 22649 9367 22707 9373
rect 17644 9324 17650 9336
rect 22649 9333 22661 9367
rect 22695 9364 22707 9367
rect 22922 9364 22928 9376
rect 22695 9336 22928 9364
rect 22695 9333 22707 9336
rect 22649 9327 22707 9333
rect 22922 9324 22928 9336
rect 22980 9324 22986 9376
rect 24578 9324 24584 9376
rect 24636 9364 24642 9376
rect 25133 9367 25191 9373
rect 25133 9364 25145 9367
rect 24636 9336 25145 9364
rect 24636 9324 24642 9336
rect 25133 9333 25145 9336
rect 25179 9364 25191 9367
rect 26418 9364 26424 9376
rect 25179 9336 26424 9364
rect 25179 9333 25191 9336
rect 25133 9327 25191 9333
rect 26418 9324 26424 9336
rect 26476 9364 26482 9376
rect 29086 9364 29092 9376
rect 26476 9336 29092 9364
rect 26476 9324 26482 9336
rect 29086 9324 29092 9336
rect 29144 9324 29150 9376
rect 30926 9324 30932 9376
rect 30984 9324 30990 9376
rect 33410 9324 33416 9376
rect 33468 9324 33474 9376
rect 34698 9324 34704 9376
rect 34756 9364 34762 9376
rect 34808 9364 34836 9463
rect 35434 9460 35440 9472
rect 35492 9460 35498 9512
rect 35618 9460 35624 9512
rect 35676 9460 35682 9512
rect 35802 9460 35808 9512
rect 35860 9460 35866 9512
rect 35912 9500 35940 9540
rect 36538 9528 36544 9580
rect 36596 9528 36602 9580
rect 36814 9528 36820 9580
rect 36872 9528 36878 9580
rect 36906 9528 36912 9580
rect 36964 9528 36970 9580
rect 37016 9568 37044 9608
rect 37093 9605 37105 9639
rect 37139 9636 37151 9639
rect 37182 9636 37188 9648
rect 37139 9608 37188 9636
rect 37139 9605 37151 9608
rect 37093 9599 37151 9605
rect 37182 9596 37188 9608
rect 37240 9596 37246 9648
rect 37274 9568 37280 9580
rect 37016 9540 37280 9568
rect 37274 9528 37280 9540
rect 37332 9528 37338 9580
rect 36722 9500 36728 9512
rect 35912 9472 36728 9500
rect 36722 9460 36728 9472
rect 36780 9460 36786 9512
rect 37093 9503 37151 9509
rect 37093 9469 37105 9503
rect 37139 9500 37151 9503
rect 37458 9500 37464 9512
rect 37139 9472 37464 9500
rect 37139 9469 37151 9472
rect 37093 9463 37151 9469
rect 34974 9392 34980 9444
rect 35032 9432 35038 9444
rect 35032 9404 36032 9432
rect 35032 9392 35038 9404
rect 34756 9336 34836 9364
rect 34756 9324 34762 9336
rect 34882 9324 34888 9376
rect 34940 9364 34946 9376
rect 35268 9373 35296 9404
rect 35069 9367 35127 9373
rect 35069 9364 35081 9367
rect 34940 9336 35081 9364
rect 34940 9324 34946 9336
rect 35069 9333 35081 9336
rect 35115 9333 35127 9367
rect 35069 9327 35127 9333
rect 35253 9367 35311 9373
rect 35253 9333 35265 9367
rect 35299 9333 35311 9367
rect 35253 9327 35311 9333
rect 35713 9367 35771 9373
rect 35713 9333 35725 9367
rect 35759 9364 35771 9367
rect 35894 9364 35900 9376
rect 35759 9336 35900 9364
rect 35759 9333 35771 9336
rect 35713 9327 35771 9333
rect 35894 9324 35900 9336
rect 35952 9324 35958 9376
rect 36004 9364 36032 9404
rect 36170 9392 36176 9444
rect 36228 9432 36234 9444
rect 36998 9432 37004 9444
rect 36228 9404 37004 9432
rect 36228 9392 36234 9404
rect 36998 9392 37004 9404
rect 37056 9432 37062 9444
rect 37108 9432 37136 9463
rect 37458 9460 37464 9472
rect 37516 9460 37522 9512
rect 37056 9404 37136 9432
rect 37056 9392 37062 9404
rect 36081 9367 36139 9373
rect 36081 9364 36093 9367
rect 36004 9336 36093 9364
rect 36081 9333 36093 9336
rect 36127 9333 36139 9367
rect 36081 9327 36139 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 8110 9120 8116 9172
rect 8168 9120 8174 9172
rect 9398 9120 9404 9172
rect 9456 9160 9462 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9456 9132 9689 9160
rect 9456 9120 9462 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 10229 9163 10287 9169
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 10962 9160 10968 9172
rect 10275 9132 10968 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 14608 9132 15025 9160
rect 14608 9120 14614 9132
rect 15013 9129 15025 9132
rect 15059 9129 15071 9163
rect 15013 9123 15071 9129
rect 16390 9120 16396 9172
rect 16448 9120 16454 9172
rect 16758 9120 16764 9172
rect 16816 9120 16822 9172
rect 16942 9120 16948 9172
rect 17000 9120 17006 9172
rect 17954 9120 17960 9172
rect 18012 9120 18018 9172
rect 26142 9120 26148 9172
rect 26200 9160 26206 9172
rect 26237 9163 26295 9169
rect 26237 9160 26249 9163
rect 26200 9132 26249 9160
rect 26200 9120 26206 9132
rect 26237 9129 26249 9132
rect 26283 9129 26295 9163
rect 26237 9123 26295 9129
rect 28166 9120 28172 9172
rect 28224 9120 28230 9172
rect 28350 9120 28356 9172
rect 28408 9120 28414 9172
rect 30009 9163 30067 9169
rect 30009 9160 30021 9163
rect 29656 9132 30021 9160
rect 14277 9095 14335 9101
rect 14277 9061 14289 9095
rect 14323 9092 14335 9095
rect 15378 9092 15384 9104
rect 14323 9064 15384 9092
rect 14323 9061 14335 9064
rect 14277 9055 14335 9061
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 21637 9095 21695 9101
rect 21637 9061 21649 9095
rect 21683 9092 21695 9095
rect 21726 9092 21732 9104
rect 21683 9064 21732 9092
rect 21683 9061 21695 9064
rect 21637 9055 21695 9061
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 25774 9092 25780 9104
rect 25056 9064 25780 9092
rect 6638 8984 6644 9036
rect 6696 8984 6702 9036
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 13170 9024 13176 9036
rect 11931 8996 13176 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8925 6423 8959
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 7774 8928 8677 8956
rect 6365 8919 6423 8925
rect 8665 8925 8677 8928
rect 8711 8956 8723 8959
rect 9490 8956 9496 8968
rect 8711 8928 9496 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 6380 8888 6408 8919
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 9674 8916 9680 8968
rect 9732 8916 9738 8968
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 9950 8956 9956 8968
rect 9907 8928 9956 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 11606 8956 11612 8968
rect 10560 8928 11612 8956
rect 10560 8916 10566 8928
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 13372 8956 13400 8987
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 18601 9027 18659 9033
rect 14056 8996 14320 9024
rect 14056 8984 14062 8996
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13372 8928 14105 8956
rect 14093 8925 14105 8928
rect 14139 8956 14151 8959
rect 14182 8956 14188 8968
rect 14139 8928 14188 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 14292 8965 14320 8996
rect 16500 8996 16896 9024
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15197 8959 15255 8965
rect 15197 8956 15209 8959
rect 14976 8928 15209 8956
rect 14976 8916 14982 8928
rect 15197 8925 15209 8928
rect 15243 8925 15255 8959
rect 15197 8919 15255 8925
rect 15286 8916 15292 8968
rect 15344 8916 15350 8968
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 16500 8965 16528 8996
rect 16868 8965 16896 8996
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 18690 9024 18696 9036
rect 18647 8996 18696 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 18690 8984 18696 8996
rect 18748 8984 18754 9036
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15896 8928 16129 8956
rect 15896 8916 15902 8928
rect 16117 8925 16129 8928
rect 16163 8956 16175 8959
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 16163 8928 16497 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 6546 8888 6552 8900
rect 5500 8860 6552 8888
rect 5500 8848 5506 8860
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 8294 8848 8300 8900
rect 8352 8848 8358 8900
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 10413 8891 10471 8897
rect 8628 8860 10272 8888
rect 8628 8848 8634 8860
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 8312 8820 8340 8848
rect 10244 8829 10272 8860
rect 10413 8857 10425 8891
rect 10459 8888 10471 8891
rect 10870 8888 10876 8900
rect 10459 8860 10876 8888
rect 10459 8857 10471 8860
rect 10413 8851 10471 8857
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 13446 8888 13452 8900
rect 13110 8860 13452 8888
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 15010 8848 15016 8900
rect 15068 8848 15074 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 15120 8860 16313 8888
rect 15120 8832 15148 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 16592 8888 16620 8919
rect 18322 8916 18328 8968
rect 18380 8916 18386 8968
rect 21913 8959 21971 8965
rect 21913 8925 21925 8959
rect 21959 8956 21971 8959
rect 23198 8956 23204 8968
rect 21959 8928 23204 8956
rect 21959 8925 21971 8928
rect 21913 8919 21971 8925
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 25056 8965 25084 9064
rect 25774 9052 25780 9064
rect 25832 9052 25838 9104
rect 25869 9095 25927 9101
rect 25869 9061 25881 9095
rect 25915 9092 25927 9095
rect 28184 9092 28212 9120
rect 25915 9064 27384 9092
rect 28184 9064 29132 9092
rect 25915 9061 25927 9064
rect 25869 9055 25927 9061
rect 26050 8984 26056 9036
rect 26108 9024 26114 9036
rect 26108 8996 26188 9024
rect 26108 8984 26114 8996
rect 25041 8959 25099 8965
rect 25041 8925 25053 8959
rect 25087 8925 25099 8959
rect 25041 8919 25099 8925
rect 25222 8916 25228 8968
rect 25280 8916 25286 8968
rect 26160 8965 26188 8996
rect 25317 8959 25375 8965
rect 25317 8925 25329 8959
rect 25363 8925 25375 8959
rect 25317 8919 25375 8925
rect 26145 8959 26203 8965
rect 26145 8925 26157 8959
rect 26191 8925 26203 8959
rect 26145 8919 26203 8925
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8956 26295 8959
rect 26326 8956 26332 8968
rect 26283 8928 26332 8956
rect 26283 8925 26295 8928
rect 26237 8919 26295 8925
rect 16301 8851 16359 8857
rect 16500 8860 16620 8888
rect 16500 8832 16528 8860
rect 21634 8848 21640 8900
rect 21692 8888 21698 8900
rect 25332 8888 25360 8919
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 26421 8959 26479 8965
rect 26421 8925 26433 8959
rect 26467 8925 26479 8959
rect 27356 8956 27384 9064
rect 27816 8996 28488 9024
rect 27816 8965 27844 8996
rect 28460 8965 28488 8996
rect 27801 8959 27859 8965
rect 27801 8956 27813 8959
rect 27356 8928 27813 8956
rect 26421 8919 26479 8925
rect 27801 8925 27813 8928
rect 27847 8925 27859 8959
rect 27801 8919 27859 8925
rect 28261 8959 28319 8965
rect 28261 8925 28273 8959
rect 28307 8925 28319 8959
rect 28261 8919 28319 8925
rect 28445 8959 28503 8965
rect 28445 8925 28457 8959
rect 28491 8925 28503 8959
rect 29104 8956 29132 9064
rect 29656 8965 29684 9132
rect 30009 9129 30021 9132
rect 30055 9129 30067 9163
rect 30009 9123 30067 9129
rect 30929 9163 30987 9169
rect 30929 9129 30941 9163
rect 30975 9160 30987 9163
rect 31018 9160 31024 9172
rect 30975 9132 31024 9160
rect 30975 9129 30987 9132
rect 30929 9123 30987 9129
rect 31018 9120 31024 9132
rect 31076 9120 31082 9172
rect 31849 9163 31907 9169
rect 31849 9129 31861 9163
rect 31895 9160 31907 9163
rect 32674 9160 32680 9172
rect 31895 9132 32680 9160
rect 31895 9129 31907 9132
rect 31849 9123 31907 9129
rect 32674 9120 32680 9132
rect 32732 9120 32738 9172
rect 35342 9120 35348 9172
rect 35400 9160 35406 9172
rect 35802 9160 35808 9172
rect 35400 9132 35808 9160
rect 35400 9120 35406 9132
rect 35802 9120 35808 9132
rect 35860 9160 35866 9172
rect 36170 9160 36176 9172
rect 35860 9132 36176 9160
rect 35860 9120 35866 9132
rect 36170 9120 36176 9132
rect 36228 9120 36234 9172
rect 36722 9120 36728 9172
rect 36780 9160 36786 9172
rect 38381 9163 38439 9169
rect 38381 9160 38393 9163
rect 36780 9132 38393 9160
rect 36780 9120 36786 9132
rect 38381 9129 38393 9132
rect 38427 9129 38439 9163
rect 38381 9123 38439 9129
rect 30377 9095 30435 9101
rect 30377 9061 30389 9095
rect 30423 9092 30435 9095
rect 30423 9064 30604 9092
rect 30423 9061 30435 9064
rect 30377 9055 30435 9061
rect 30576 9033 30604 9064
rect 33962 9052 33968 9104
rect 34020 9092 34026 9104
rect 34020 9064 35112 9092
rect 34020 9052 34026 9064
rect 29917 9027 29975 9033
rect 29917 8993 29929 9027
rect 29963 9024 29975 9027
rect 30561 9027 30619 9033
rect 29963 8996 30144 9024
rect 29963 8993 29975 8996
rect 29917 8987 29975 8993
rect 30116 8968 30144 8996
rect 30561 8993 30573 9027
rect 30607 9024 30619 9027
rect 31294 9024 31300 9036
rect 30607 8996 31300 9024
rect 30607 8993 30619 8996
rect 30561 8987 30619 8993
rect 31294 8984 31300 8996
rect 31352 8984 31358 9036
rect 34514 8984 34520 9036
rect 34572 9024 34578 9036
rect 35084 9033 35112 9064
rect 34793 9027 34851 9033
rect 34793 9024 34805 9027
rect 34572 8996 34805 9024
rect 34572 8984 34578 8996
rect 34793 8993 34805 8996
rect 34839 8993 34851 9027
rect 34793 8987 34851 8993
rect 35069 9027 35127 9033
rect 35069 8993 35081 9027
rect 35115 8993 35127 9027
rect 35069 8987 35127 8993
rect 36630 8984 36636 9036
rect 36688 8984 36694 9036
rect 29641 8959 29699 8965
rect 29641 8956 29653 8959
rect 29104 8928 29653 8956
rect 28445 8919 28503 8925
rect 29641 8925 29653 8928
rect 29687 8925 29699 8959
rect 29641 8919 29699 8925
rect 21692 8860 25360 8888
rect 21692 8848 21698 8860
rect 25590 8848 25596 8900
rect 25648 8888 25654 8900
rect 25869 8891 25927 8897
rect 25869 8888 25881 8891
rect 25648 8860 25881 8888
rect 25648 8848 25654 8860
rect 25869 8857 25881 8860
rect 25915 8857 25927 8891
rect 25869 8851 25927 8857
rect 7064 8792 8340 8820
rect 10229 8823 10287 8829
rect 7064 8780 7070 8792
rect 10229 8789 10241 8823
rect 10275 8820 10287 8823
rect 10686 8820 10692 8832
rect 10275 8792 10692 8820
rect 10275 8789 10287 8792
rect 10229 8783 10287 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 14829 8823 14887 8829
rect 14829 8789 14841 8823
rect 14875 8820 14887 8823
rect 15102 8820 15108 8832
rect 14875 8792 15108 8820
rect 14875 8789 14887 8792
rect 14829 8783 14887 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15562 8780 15568 8832
rect 15620 8780 15626 8832
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 16482 8820 16488 8832
rect 15712 8792 16488 8820
rect 15712 8780 15718 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 18417 8823 18475 8829
rect 18417 8789 18429 8823
rect 18463 8820 18475 8823
rect 18690 8820 18696 8832
rect 18463 8792 18696 8820
rect 18463 8789 18475 8792
rect 18417 8783 18475 8789
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 21818 8780 21824 8832
rect 21876 8780 21882 8832
rect 25225 8823 25283 8829
rect 25225 8789 25237 8823
rect 25271 8820 25283 8823
rect 25406 8820 25412 8832
rect 25271 8792 25412 8820
rect 25271 8789 25283 8792
rect 25225 8783 25283 8789
rect 25406 8780 25412 8792
rect 25464 8780 25470 8832
rect 25498 8780 25504 8832
rect 25556 8780 25562 8832
rect 25884 8820 25912 8851
rect 25958 8848 25964 8900
rect 26016 8888 26022 8900
rect 26053 8891 26111 8897
rect 26053 8888 26065 8891
rect 26016 8860 26065 8888
rect 26016 8848 26022 8860
rect 26053 8857 26065 8860
rect 26099 8857 26111 8891
rect 26053 8851 26111 8857
rect 26436 8820 26464 8919
rect 27982 8848 27988 8900
rect 28040 8888 28046 8900
rect 28276 8888 28304 8919
rect 29730 8916 29736 8968
rect 29788 8956 29794 8968
rect 30009 8959 30067 8965
rect 30009 8956 30021 8959
rect 29788 8928 30021 8956
rect 29788 8916 29794 8928
rect 30009 8925 30021 8928
rect 30055 8925 30067 8959
rect 30009 8919 30067 8925
rect 30098 8916 30104 8968
rect 30156 8916 30162 8968
rect 30745 8959 30803 8965
rect 30745 8925 30757 8959
rect 30791 8925 30803 8959
rect 30745 8919 30803 8925
rect 31665 8959 31723 8965
rect 31665 8925 31677 8959
rect 31711 8956 31723 8959
rect 31754 8956 31760 8968
rect 31711 8928 31760 8956
rect 31711 8925 31723 8928
rect 31665 8919 31723 8925
rect 28040 8860 28304 8888
rect 29917 8891 29975 8897
rect 28040 8848 28046 8860
rect 29917 8857 29929 8891
rect 29963 8888 29975 8891
rect 30760 8888 30788 8919
rect 31754 8916 31760 8928
rect 31812 8916 31818 8968
rect 31846 8916 31852 8968
rect 31904 8916 31910 8968
rect 34698 8916 34704 8968
rect 34756 8956 34762 8968
rect 34885 8959 34943 8965
rect 34885 8956 34897 8959
rect 34756 8928 34897 8956
rect 34756 8916 34762 8928
rect 34885 8925 34897 8928
rect 34931 8925 34943 8959
rect 34885 8919 34943 8925
rect 34977 8959 35035 8965
rect 34977 8925 34989 8959
rect 35023 8956 35035 8959
rect 35526 8956 35532 8968
rect 35023 8928 35532 8956
rect 35023 8925 35035 8928
rect 34977 8919 35035 8925
rect 29963 8860 30788 8888
rect 29963 8857 29975 8860
rect 29917 8851 29975 8857
rect 34330 8848 34336 8900
rect 34388 8888 34394 8900
rect 34992 8888 35020 8919
rect 35526 8916 35532 8928
rect 35584 8916 35590 8968
rect 36446 8916 36452 8968
rect 36504 8916 36510 8968
rect 34388 8860 35020 8888
rect 34388 8848 34394 8860
rect 36906 8848 36912 8900
rect 36964 8848 36970 8900
rect 37366 8848 37372 8900
rect 37424 8848 37430 8900
rect 25884 8792 26464 8820
rect 35250 8780 35256 8832
rect 35308 8780 35314 8832
rect 36170 8780 36176 8832
rect 36228 8820 36234 8832
rect 36265 8823 36323 8829
rect 36265 8820 36277 8823
rect 36228 8792 36277 8820
rect 36228 8780 36234 8792
rect 36265 8789 36277 8792
rect 36311 8789 36323 8823
rect 36265 8783 36323 8789
rect 1104 8730 38824 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 38824 8730
rect 1104 8656 38824 8678
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5408 8588 5457 8616
rect 5408 8576 5414 8588
rect 5445 8585 5457 8588
rect 5491 8616 5503 8619
rect 5491 8588 7328 8616
rect 5491 8585 5503 8588
rect 5445 8579 5503 8585
rect 4798 8548 4804 8560
rect 3988 8520 4804 8548
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 3988 8489 4016 8520
rect 4798 8508 4804 8520
rect 4856 8548 4862 8560
rect 5608 8551 5666 8557
rect 5608 8548 5620 8551
rect 4856 8520 5620 8548
rect 4856 8508 4862 8520
rect 5608 8517 5620 8520
rect 5654 8548 5666 8551
rect 5813 8551 5871 8557
rect 5654 8517 5672 8548
rect 5608 8511 5672 8517
rect 5813 8517 5825 8551
rect 5859 8548 5871 8551
rect 6822 8548 6828 8560
rect 5859 8520 6828 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3936 8452 3985 8480
rect 3936 8440 3942 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4706 8480 4712 8492
rect 4203 8452 4712 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5184 8344 5212 8443
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5644 8480 5672 8511
rect 6822 8508 6828 8520
rect 6880 8548 6886 8560
rect 6880 8520 7144 8548
rect 6880 8508 6886 8520
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5644 8452 5917 8480
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 7116 8489 7144 8520
rect 7300 8492 7328 8588
rect 7760 8588 9628 8616
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6227 8452 6561 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7760 8489 7788 8588
rect 8021 8551 8079 8557
rect 8021 8517 8033 8551
rect 8067 8548 8079 8551
rect 8294 8548 8300 8560
rect 8067 8520 8300 8548
rect 8067 8517 8079 8520
rect 8021 8511 8079 8517
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 9490 8548 9496 8560
rect 9246 8520 9496 8548
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7484 8356 7512 8443
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 8570 8412 8576 8424
rect 7699 8384 8576 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 9600 8421 9628 8588
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 14458 8616 14464 8628
rect 11664 8588 14464 8616
rect 11664 8576 11670 8588
rect 9766 8508 9772 8560
rect 9824 8548 9830 8560
rect 9824 8520 10350 8548
rect 9824 8508 9830 8520
rect 12544 8489 12572 8588
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15562 8616 15568 8628
rect 15243 8588 15568 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15562 8576 15568 8588
rect 15620 8616 15626 8628
rect 16117 8619 16175 8625
rect 16117 8616 16129 8619
rect 15620 8588 16129 8616
rect 15620 8576 15626 8588
rect 16117 8585 16129 8588
rect 16163 8585 16175 8619
rect 16117 8579 16175 8585
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17681 8619 17739 8625
rect 17681 8616 17693 8619
rect 17368 8588 17693 8616
rect 17368 8576 17374 8588
rect 17681 8585 17693 8588
rect 17727 8616 17739 8619
rect 18690 8616 18696 8628
rect 17727 8588 18696 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 22278 8576 22284 8628
rect 22336 8616 22342 8628
rect 23201 8619 23259 8625
rect 23201 8616 23213 8619
rect 22336 8588 23213 8616
rect 22336 8576 22342 8588
rect 23201 8585 23213 8588
rect 23247 8585 23259 8619
rect 24854 8616 24860 8628
rect 23201 8579 23259 8585
rect 23952 8588 24860 8616
rect 20996 8560 21048 8566
rect 12802 8508 12808 8560
rect 12860 8508 12866 8560
rect 13446 8508 13452 8560
rect 13504 8508 13510 8560
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 15289 8551 15347 8557
rect 15289 8548 15301 8551
rect 15160 8520 15301 8548
rect 15160 8508 15166 8520
rect 15289 8517 15301 8520
rect 15335 8517 15347 8551
rect 15289 8511 15347 8517
rect 16025 8551 16083 8557
rect 16025 8517 16037 8551
rect 16071 8548 16083 8551
rect 16390 8548 16396 8560
rect 16071 8520 16396 8548
rect 16071 8517 16083 8520
rect 16025 8511 16083 8517
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 21453 8551 21511 8557
rect 21453 8517 21465 8551
rect 21499 8548 21511 8551
rect 21818 8548 21824 8560
rect 21499 8520 21824 8548
rect 21499 8517 21511 8520
rect 21453 8511 21511 8517
rect 21818 8508 21824 8520
rect 21876 8548 21882 8560
rect 21876 8520 23796 8548
rect 21876 8508 21882 8520
rect 20996 8502 21048 8508
rect 22480 8492 22508 8520
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 16224 8452 18000 8480
rect 16224 8424 16252 8452
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9631 8384 9720 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 5184 8316 6193 8344
rect 6181 8313 6193 8316
rect 6227 8313 6239 8347
rect 6181 8307 6239 8313
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 7524 8316 7880 8344
rect 7524 8304 7530 8316
rect 2866 8236 2872 8288
rect 2924 8276 2930 8288
rect 3973 8279 4031 8285
rect 3973 8276 3985 8279
rect 2924 8248 3985 8276
rect 2924 8236 2930 8248
rect 3973 8245 3985 8248
rect 4019 8245 4031 8279
rect 3973 8239 4031 8245
rect 5350 8236 5356 8288
rect 5408 8236 5414 8288
rect 5629 8279 5687 8285
rect 5629 8245 5641 8279
rect 5675 8276 5687 8279
rect 5994 8276 6000 8288
rect 5675 8248 6000 8276
rect 5675 8245 5687 8248
rect 5629 8239 5687 8245
rect 5994 8236 6000 8248
rect 6052 8276 6058 8288
rect 6730 8276 6736 8288
rect 6052 8248 6736 8276
rect 6052 8236 6058 8248
rect 6730 8236 6736 8248
rect 6788 8276 6794 8288
rect 7742 8276 7748 8288
rect 6788 8248 7748 8276
rect 6788 8236 6794 8248
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 7852 8276 7880 8316
rect 9122 8276 9128 8288
rect 7852 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8276 9186 8288
rect 9493 8279 9551 8285
rect 9493 8276 9505 8279
rect 9180 8248 9505 8276
rect 9180 8236 9186 8248
rect 9493 8245 9505 8248
rect 9539 8245 9551 8279
rect 9692 8276 9720 8384
rect 9858 8372 9864 8424
rect 9916 8372 9922 8424
rect 11333 8415 11391 8421
rect 11333 8381 11345 8415
rect 11379 8412 11391 8415
rect 11698 8412 11704 8424
rect 11379 8384 11704 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 11698 8372 11704 8384
rect 11756 8412 11762 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 11756 8384 12081 8412
rect 11756 8372 11762 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 14274 8372 14280 8424
rect 14332 8372 14338 8424
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 16206 8412 16212 8424
rect 15519 8384 16212 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 17770 8372 17776 8424
rect 17828 8372 17834 8424
rect 17972 8421 18000 8452
rect 22462 8440 22468 8492
rect 22520 8440 22526 8492
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8480 22891 8483
rect 23198 8480 23204 8492
rect 22879 8452 23204 8480
rect 22879 8449 22891 8452
rect 22833 8443 22891 8449
rect 23198 8440 23204 8452
rect 23256 8480 23262 8492
rect 23385 8483 23443 8489
rect 23385 8480 23397 8483
rect 23256 8452 23397 8480
rect 23256 8440 23262 8452
rect 23385 8449 23397 8452
rect 23431 8449 23443 8483
rect 23385 8443 23443 8449
rect 17957 8415 18015 8421
rect 17957 8381 17969 8415
rect 18003 8412 18015 8415
rect 18598 8412 18604 8424
rect 18003 8384 18604 8412
rect 18003 8381 18015 8384
rect 17957 8375 18015 8381
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 19610 8372 19616 8424
rect 19668 8372 19674 8424
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20027 8384 21036 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 21008 8344 21036 8384
rect 21450 8372 21456 8424
rect 21508 8412 21514 8424
rect 21913 8415 21971 8421
rect 21913 8412 21925 8415
rect 21508 8384 21925 8412
rect 21508 8372 21514 8384
rect 21913 8381 21925 8384
rect 21959 8412 21971 8415
rect 23400 8412 23428 8443
rect 23474 8440 23480 8492
rect 23532 8440 23538 8492
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8449 23719 8483
rect 23661 8443 23719 8449
rect 23676 8412 23704 8443
rect 21959 8384 23336 8412
rect 23400 8384 23704 8412
rect 23768 8412 23796 8520
rect 23842 8440 23848 8492
rect 23900 8440 23906 8492
rect 23952 8489 23980 8588
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 25777 8619 25835 8625
rect 25777 8616 25789 8619
rect 25280 8588 25789 8616
rect 25280 8576 25286 8588
rect 25777 8585 25789 8588
rect 25823 8616 25835 8619
rect 26326 8616 26332 8628
rect 25823 8588 26332 8616
rect 25823 8585 25835 8588
rect 25777 8579 25835 8585
rect 26326 8576 26332 8588
rect 26384 8576 26390 8628
rect 27525 8619 27583 8625
rect 27525 8585 27537 8619
rect 27571 8616 27583 8619
rect 27982 8616 27988 8628
rect 27571 8588 27988 8616
rect 27571 8585 27583 8588
rect 27525 8579 27583 8585
rect 27982 8576 27988 8588
rect 28040 8576 28046 8628
rect 29181 8619 29239 8625
rect 29181 8585 29193 8619
rect 29227 8616 29239 8619
rect 29730 8616 29736 8628
rect 29227 8588 29736 8616
rect 29227 8585 29239 8588
rect 29181 8579 29239 8585
rect 29730 8576 29736 8588
rect 29788 8576 29794 8628
rect 31294 8576 31300 8628
rect 31352 8576 31358 8628
rect 31662 8576 31668 8628
rect 31720 8625 31726 8628
rect 31720 8619 31739 8625
rect 31727 8585 31739 8619
rect 31720 8579 31739 8585
rect 31720 8576 31726 8579
rect 31846 8576 31852 8628
rect 31904 8576 31910 8628
rect 35250 8576 35256 8628
rect 35308 8576 35314 8628
rect 36725 8619 36783 8625
rect 36725 8585 36737 8619
rect 36771 8616 36783 8619
rect 36906 8616 36912 8628
rect 36771 8588 36912 8616
rect 36771 8585 36783 8588
rect 36725 8579 36783 8585
rect 36906 8576 36912 8588
rect 36964 8576 36970 8628
rect 25590 8548 25596 8560
rect 25240 8520 25596 8548
rect 25240 8492 25268 8520
rect 25590 8508 25596 8520
rect 25648 8508 25654 8560
rect 27430 8548 27436 8560
rect 25700 8520 27436 8548
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24029 8483 24087 8489
rect 24029 8449 24041 8483
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 24578 8480 24584 8492
rect 24443 8452 24584 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24044 8412 24072 8443
rect 24578 8440 24584 8452
rect 24636 8440 24642 8492
rect 25222 8440 25228 8492
rect 25280 8440 25286 8492
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 25424 8412 25452 8443
rect 25498 8440 25504 8492
rect 25556 8480 25562 8492
rect 25700 8489 25728 8520
rect 27430 8508 27436 8520
rect 27488 8508 27494 8560
rect 28169 8551 28227 8557
rect 28169 8517 28181 8551
rect 28215 8548 28227 8551
rect 28626 8548 28632 8560
rect 28215 8520 28632 8548
rect 28215 8517 28227 8520
rect 28169 8511 28227 8517
rect 28626 8508 28632 8520
rect 28684 8548 28690 8560
rect 28997 8551 29055 8557
rect 28997 8548 29009 8551
rect 28684 8520 29009 8548
rect 28684 8508 28690 8520
rect 28997 8517 29009 8520
rect 29043 8517 29055 8551
rect 31481 8551 31539 8557
rect 31481 8548 31493 8551
rect 28997 8511 29055 8517
rect 31128 8520 31493 8548
rect 31128 8492 31156 8520
rect 31481 8517 31493 8520
rect 31527 8517 31539 8551
rect 31481 8511 31539 8517
rect 25685 8483 25743 8489
rect 25685 8480 25697 8483
rect 25556 8452 25697 8480
rect 25556 8440 25562 8452
rect 25685 8449 25697 8452
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25869 8483 25927 8489
rect 25869 8449 25881 8483
rect 25915 8480 25927 8483
rect 25961 8483 26019 8489
rect 25961 8480 25973 8483
rect 25915 8452 25973 8480
rect 25915 8449 25927 8452
rect 25869 8443 25927 8449
rect 25961 8449 25973 8452
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 26053 8483 26111 8489
rect 26053 8449 26065 8483
rect 26099 8480 26111 8483
rect 26234 8480 26240 8492
rect 26099 8452 26240 8480
rect 26099 8449 26111 8452
rect 26053 8443 26111 8449
rect 25884 8412 25912 8443
rect 26234 8440 26240 8452
rect 26292 8480 26298 8492
rect 27154 8480 27160 8492
rect 26292 8452 27160 8480
rect 26292 8440 26298 8452
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 28074 8440 28080 8492
rect 28132 8440 28138 8492
rect 28258 8440 28264 8492
rect 28316 8480 28322 8492
rect 28537 8483 28595 8489
rect 28537 8480 28549 8483
rect 28316 8452 28549 8480
rect 28316 8440 28322 8452
rect 28537 8449 28549 8452
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 28721 8483 28779 8489
rect 28721 8449 28733 8483
rect 28767 8480 28779 8483
rect 28813 8483 28871 8489
rect 28813 8480 28825 8483
rect 28767 8452 28825 8480
rect 28767 8449 28779 8452
rect 28721 8443 28779 8449
rect 28813 8449 28825 8452
rect 28859 8449 28871 8483
rect 28813 8443 28871 8449
rect 31110 8440 31116 8492
rect 31168 8440 31174 8492
rect 31389 8483 31447 8489
rect 31389 8449 31401 8483
rect 31435 8480 31447 8483
rect 31680 8480 31708 8576
rect 33873 8551 33931 8557
rect 33873 8517 33885 8551
rect 33919 8548 33931 8551
rect 33962 8548 33968 8560
rect 33919 8520 33968 8548
rect 33919 8517 33931 8520
rect 33873 8511 33931 8517
rect 33962 8508 33968 8520
rect 34020 8548 34026 8560
rect 34020 8520 34560 8548
rect 34020 8508 34026 8520
rect 31435 8452 31708 8480
rect 34057 8483 34115 8489
rect 31435 8449 31447 8452
rect 31389 8443 31447 8449
rect 34057 8449 34069 8483
rect 34103 8480 34115 8483
rect 34330 8480 34336 8492
rect 34103 8452 34336 8480
rect 34103 8449 34115 8452
rect 34057 8443 34115 8449
rect 34330 8440 34336 8452
rect 34388 8440 34394 8492
rect 34532 8489 34560 8520
rect 34517 8483 34575 8489
rect 34517 8449 34529 8483
rect 34563 8480 34575 8483
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 34563 8452 34897 8480
rect 34563 8449 34575 8452
rect 34517 8443 34575 8449
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 34885 8443 34943 8449
rect 35986 8440 35992 8492
rect 36044 8480 36050 8492
rect 36633 8483 36691 8489
rect 36633 8480 36645 8483
rect 36044 8452 36645 8480
rect 36044 8440 36050 8452
rect 36633 8449 36645 8452
rect 36679 8449 36691 8483
rect 36633 8443 36691 8449
rect 36817 8483 36875 8489
rect 36817 8449 36829 8483
rect 36863 8480 36875 8483
rect 37274 8480 37280 8492
rect 36863 8452 37280 8480
rect 36863 8449 36875 8452
rect 36817 8443 36875 8449
rect 37274 8440 37280 8452
rect 37332 8440 37338 8492
rect 23768 8384 25912 8412
rect 21959 8381 21971 8384
rect 21913 8375 21971 8381
rect 22370 8344 22376 8356
rect 21008 8316 22376 8344
rect 22370 8304 22376 8316
rect 22428 8304 22434 8356
rect 23308 8344 23336 8384
rect 27062 8372 27068 8424
rect 27120 8372 27126 8424
rect 28092 8412 28120 8440
rect 28353 8415 28411 8421
rect 28353 8412 28365 8415
rect 28092 8384 28365 8412
rect 28353 8381 28365 8384
rect 28399 8381 28411 8415
rect 28353 8375 28411 8381
rect 34606 8372 34612 8424
rect 34664 8372 34670 8424
rect 34790 8372 34796 8424
rect 34848 8372 34854 8424
rect 24489 8347 24547 8353
rect 23308 8316 24440 8344
rect 10502 8276 10508 8288
rect 9692 8248 10508 8276
rect 9493 8239 9551 8245
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 11514 8236 11520 8288
rect 11572 8236 11578 8288
rect 14366 8236 14372 8288
rect 14424 8276 14430 8288
rect 14829 8279 14887 8285
rect 14829 8276 14841 8279
rect 14424 8248 14841 8276
rect 14424 8236 14430 8248
rect 14829 8245 14841 8248
rect 14875 8245 14887 8279
rect 14829 8239 14887 8245
rect 15654 8236 15660 8288
rect 15712 8236 15718 8288
rect 17218 8236 17224 8288
rect 17276 8276 17282 8288
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 17276 8248 17325 8276
rect 17276 8236 17282 8248
rect 17313 8245 17325 8248
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 24302 8236 24308 8288
rect 24360 8236 24366 8288
rect 24412 8276 24440 8316
rect 24489 8313 24501 8347
rect 24535 8344 24547 8347
rect 24854 8344 24860 8356
rect 24535 8316 24860 8344
rect 24535 8313 24547 8316
rect 24489 8307 24547 8313
rect 24854 8304 24860 8316
rect 24912 8304 24918 8356
rect 31113 8347 31171 8353
rect 31113 8313 31125 8347
rect 31159 8344 31171 8347
rect 31754 8344 31760 8356
rect 31159 8316 31760 8344
rect 31159 8313 31171 8316
rect 31113 8307 31171 8313
rect 31754 8304 31760 8316
rect 31812 8304 31818 8356
rect 34241 8347 34299 8353
rect 34241 8313 34253 8347
rect 34287 8344 34299 8347
rect 34287 8316 34836 8344
rect 34287 8313 34299 8316
rect 34241 8307 34299 8313
rect 34808 8288 34836 8316
rect 24946 8276 24952 8288
rect 24412 8248 24952 8276
rect 24946 8236 24952 8248
rect 25004 8276 25010 8288
rect 26602 8276 26608 8288
rect 25004 8248 26608 8276
rect 25004 8236 25010 8248
rect 26602 8236 26608 8248
rect 26660 8236 26666 8288
rect 31294 8236 31300 8288
rect 31352 8276 31358 8288
rect 31665 8279 31723 8285
rect 31665 8276 31677 8279
rect 31352 8248 31677 8276
rect 31352 8236 31358 8248
rect 31665 8245 31677 8248
rect 31711 8245 31723 8279
rect 31665 8239 31723 8245
rect 34422 8236 34428 8288
rect 34480 8236 34486 8288
rect 34790 8236 34796 8288
rect 34848 8236 34854 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 3878 8032 3884 8084
rect 3936 8032 3942 8084
rect 6822 8032 6828 8084
rect 6880 8032 6886 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7190 8072 7196 8084
rect 7147 8044 7196 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7466 8072 7472 8084
rect 7331 8044 7472 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 7742 8032 7748 8084
rect 7800 8032 7806 8084
rect 8294 8032 8300 8084
rect 8352 8032 8358 8084
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 9858 8072 9864 8084
rect 9723 8044 9864 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 18690 8032 18696 8084
rect 18748 8032 18754 8084
rect 23014 8032 23020 8084
rect 23072 8072 23078 8084
rect 23290 8072 23296 8084
rect 23072 8044 23296 8072
rect 23072 8032 23078 8044
rect 23290 8032 23296 8044
rect 23348 8072 23354 8084
rect 26881 8075 26939 8081
rect 23348 8044 25360 8072
rect 23348 8032 23354 8044
rect 8205 8007 8263 8013
rect 8205 7973 8217 8007
rect 8251 8004 8263 8007
rect 9582 8004 9588 8016
rect 8251 7976 9588 8004
rect 8251 7973 8263 7976
rect 8205 7967 8263 7973
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 21174 7964 21180 8016
rect 21232 8004 21238 8016
rect 21358 8004 21364 8016
rect 21232 7976 21364 8004
rect 21232 7964 21238 7976
rect 21358 7964 21364 7976
rect 21416 7964 21422 8016
rect 21637 8007 21695 8013
rect 21637 7973 21649 8007
rect 21683 8004 21695 8007
rect 24670 8004 24676 8016
rect 21683 7976 22094 8004
rect 21683 7973 21695 7976
rect 21637 7967 21695 7973
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5442 7936 5448 7948
rect 5123 7908 5448 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 7699 7908 7941 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 7929 7905 7941 7908
rect 7975 7936 7987 7939
rect 8110 7936 8116 7948
rect 7975 7908 8116 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8496 7908 9045 7936
rect 8496 7880 8524 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 9033 7899 9091 7905
rect 9950 7896 9956 7948
rect 10008 7896 10014 7948
rect 11514 7936 11520 7948
rect 10060 7908 11520 7936
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4430 7868 4436 7880
rect 4295 7840 4436 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 6880 7840 8033 7868
rect 6880 7828 6886 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 3970 7800 3976 7812
rect 3476 7772 3976 7800
rect 3476 7760 3482 7772
rect 3970 7760 3976 7772
rect 4028 7800 4034 7812
rect 4028 7772 5304 7800
rect 4028 7760 4034 7772
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 4856 7704 4997 7732
rect 4856 7692 4862 7704
rect 4985 7701 4997 7704
rect 5031 7701 5043 7735
rect 5276 7732 5304 7772
rect 5350 7760 5356 7812
rect 5408 7760 5414 7812
rect 7745 7803 7803 7809
rect 5736 7772 5842 7800
rect 5736 7732 5764 7772
rect 7745 7769 7757 7803
rect 7791 7800 7803 7803
rect 8846 7800 8852 7812
rect 7791 7772 8852 7800
rect 7791 7769 7803 7772
rect 7745 7763 7803 7769
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 7006 7732 7012 7744
rect 5276 7704 7012 7732
rect 4985 7695 5043 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 8956 7732 8984 7831
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 10060 7877 10088 7908
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 14090 7896 14096 7948
rect 14148 7896 14154 7948
rect 14366 7896 14372 7948
rect 14424 7896 14430 7948
rect 16206 7896 16212 7948
rect 16264 7896 16270 7948
rect 16390 7896 16396 7948
rect 16448 7896 16454 7948
rect 17218 7896 17224 7948
rect 17276 7896 17282 7948
rect 22066 7936 22094 7976
rect 23860 7976 24676 8004
rect 22066 7908 22784 7936
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 16945 7871 17003 7877
rect 16945 7868 16957 7871
rect 16724 7840 16957 7868
rect 16724 7828 16730 7840
rect 16945 7837 16957 7840
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 21358 7828 21364 7880
rect 21416 7828 21422 7880
rect 21450 7828 21456 7880
rect 21508 7828 21514 7880
rect 21726 7828 21732 7880
rect 21784 7828 21790 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 21836 7840 22385 7868
rect 21836 7812 21864 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 22462 7828 22468 7880
rect 22520 7828 22526 7880
rect 22756 7877 22784 7908
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 23014 7828 23020 7880
rect 23072 7828 23078 7880
rect 23290 7828 23296 7880
rect 23348 7868 23354 7880
rect 23860 7877 23888 7976
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 24946 8004 24952 8016
rect 24781 7976 24952 8004
rect 24210 7936 24216 7948
rect 24044 7908 24216 7936
rect 24044 7877 24072 7908
rect 24210 7896 24216 7908
rect 24268 7896 24274 7948
rect 23753 7871 23811 7877
rect 23753 7868 23765 7871
rect 23348 7840 23765 7868
rect 23348 7828 23354 7840
rect 23753 7837 23765 7840
rect 23799 7837 23811 7871
rect 23753 7831 23811 7837
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7837 23903 7871
rect 23845 7831 23903 7837
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24118 7828 24124 7880
rect 24176 7828 24182 7880
rect 24302 7828 24308 7880
rect 24360 7868 24366 7880
rect 24781 7877 24809 7976
rect 24946 7964 24952 7976
rect 25004 7964 25010 8016
rect 25133 8007 25191 8013
rect 25133 7973 25145 8007
rect 25179 8004 25191 8007
rect 25222 8004 25228 8016
rect 25179 7976 25228 8004
rect 25179 7973 25191 7976
rect 25133 7967 25191 7973
rect 25222 7964 25228 7976
rect 25280 7964 25286 8016
rect 25332 7936 25360 8044
rect 26881 8041 26893 8075
rect 26927 8072 26939 8075
rect 27062 8072 27068 8084
rect 26927 8044 27068 8072
rect 26927 8041 26939 8044
rect 26881 8035 26939 8041
rect 27062 8032 27068 8044
rect 27120 8072 27126 8084
rect 27157 8075 27215 8081
rect 27157 8072 27169 8075
rect 27120 8044 27169 8072
rect 27120 8032 27126 8044
rect 27157 8041 27169 8044
rect 27203 8041 27215 8075
rect 27157 8035 27215 8041
rect 31110 8032 31116 8084
rect 31168 8032 31174 8084
rect 34698 8072 34704 8084
rect 34348 8044 34704 8072
rect 28169 8007 28227 8013
rect 28169 7973 28181 8007
rect 28215 8004 28227 8007
rect 28258 8004 28264 8016
rect 28215 7976 28264 8004
rect 28215 7973 28227 7976
rect 28169 7967 28227 7973
rect 28258 7964 28264 7976
rect 28316 7964 28322 8016
rect 30098 7964 30104 8016
rect 30156 7964 30162 8016
rect 34348 8004 34376 8044
rect 34698 8032 34704 8044
rect 34756 8072 34762 8084
rect 34756 8044 36952 8072
rect 34756 8032 34762 8044
rect 34256 7976 34376 8004
rect 36357 8007 36415 8013
rect 27525 7939 27583 7945
rect 25240 7908 25360 7936
rect 26988 7908 27384 7936
rect 24404 7871 24462 7877
rect 24404 7868 24416 7871
rect 24360 7840 24416 7868
rect 24360 7828 24366 7840
rect 24404 7837 24416 7840
rect 24450 7837 24462 7871
rect 24404 7831 24462 7837
rect 24545 7871 24603 7877
rect 24545 7837 24557 7871
rect 24591 7837 24603 7871
rect 24545 7831 24603 7837
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 10318 7760 10324 7812
rect 10376 7800 10382 7812
rect 10781 7803 10839 7809
rect 10781 7800 10793 7803
rect 10376 7772 10793 7800
rect 10376 7760 10382 7772
rect 10781 7769 10793 7772
rect 10827 7769 10839 7803
rect 10781 7763 10839 7769
rect 11330 7760 11336 7812
rect 11388 7760 11394 7812
rect 15378 7760 15384 7812
rect 15436 7760 15442 7812
rect 18230 7760 18236 7812
rect 18288 7760 18294 7812
rect 21637 7803 21695 7809
rect 21637 7769 21649 7803
rect 21683 7800 21695 7803
rect 21818 7800 21824 7812
rect 21683 7772 21824 7800
rect 21683 7769 21695 7772
rect 21637 7763 21695 7769
rect 21818 7760 21824 7772
rect 21876 7760 21882 7812
rect 21913 7803 21971 7809
rect 21913 7769 21925 7803
rect 21959 7800 21971 7803
rect 22002 7800 22008 7812
rect 21959 7772 22008 7800
rect 21959 7769 21971 7772
rect 21913 7763 21971 7769
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 22557 7803 22615 7809
rect 22557 7769 22569 7803
rect 22603 7800 22615 7803
rect 22833 7803 22891 7809
rect 22833 7800 22845 7803
rect 22603 7772 22845 7800
rect 22603 7769 22615 7772
rect 22557 7763 22615 7769
rect 22833 7769 22845 7772
rect 22879 7769 22891 7803
rect 22833 7763 22891 7769
rect 23201 7803 23259 7809
rect 23201 7769 23213 7803
rect 23247 7800 23259 7803
rect 23658 7800 23664 7812
rect 23247 7772 23664 7800
rect 23247 7769 23259 7772
rect 23201 7763 23259 7769
rect 23658 7760 23664 7772
rect 23716 7760 23722 7812
rect 24210 7760 24216 7812
rect 24268 7800 24274 7812
rect 24560 7800 24588 7831
rect 24854 7828 24860 7880
rect 24912 7877 24918 7880
rect 24912 7831 24920 7877
rect 25133 7871 25191 7877
rect 25133 7837 25145 7871
rect 25179 7870 25191 7871
rect 25240 7870 25268 7908
rect 25179 7842 25268 7870
rect 25179 7837 25191 7842
rect 25133 7831 25191 7837
rect 24912 7828 24918 7831
rect 25314 7828 25320 7880
rect 25372 7828 25378 7880
rect 26786 7828 26792 7880
rect 26844 7828 26850 7880
rect 26988 7877 27016 7908
rect 27356 7880 27384 7908
rect 27525 7905 27537 7939
rect 27571 7936 27583 7939
rect 27893 7939 27951 7945
rect 27893 7936 27905 7939
rect 27571 7908 27905 7936
rect 27571 7905 27583 7908
rect 27525 7899 27583 7905
rect 27893 7905 27905 7908
rect 27939 7936 27951 7939
rect 28905 7939 28963 7945
rect 27939 7908 28488 7936
rect 27939 7905 27951 7908
rect 27893 7899 27951 7905
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 24268 7772 24588 7800
rect 24673 7803 24731 7809
rect 24268 7760 24274 7772
rect 24673 7769 24685 7803
rect 24719 7800 24731 7803
rect 24946 7800 24952 7812
rect 24719 7772 24952 7800
rect 24719 7769 24731 7772
rect 24673 7763 24731 7769
rect 24946 7760 24952 7772
rect 25004 7800 25010 7812
rect 25332 7800 25360 7828
rect 25004 7772 25360 7800
rect 27080 7800 27108 7831
rect 27338 7828 27344 7880
rect 27396 7828 27402 7880
rect 27798 7828 27804 7880
rect 27856 7868 27862 7880
rect 28460 7877 28488 7908
rect 28905 7905 28917 7939
rect 28951 7936 28963 7939
rect 29641 7939 29699 7945
rect 29641 7936 29653 7939
rect 28951 7908 29653 7936
rect 28951 7905 28963 7908
rect 28905 7899 28963 7905
rect 29641 7905 29653 7908
rect 29687 7936 29699 7939
rect 30929 7939 30987 7945
rect 29687 7908 30236 7936
rect 29687 7905 29699 7908
rect 29641 7899 29699 7905
rect 28261 7871 28319 7877
rect 28261 7868 28273 7871
rect 27856 7840 28273 7868
rect 27856 7828 27862 7840
rect 28261 7837 28273 7840
rect 28307 7837 28319 7871
rect 28261 7831 28319 7837
rect 28445 7871 28503 7877
rect 28445 7837 28457 7871
rect 28491 7837 28503 7871
rect 28445 7831 28503 7837
rect 28626 7828 28632 7880
rect 28684 7868 28690 7880
rect 30208 7877 30236 7908
rect 30929 7905 30941 7939
rect 30975 7936 30987 7939
rect 30975 7908 31432 7936
rect 30975 7905 30987 7908
rect 30929 7899 30987 7905
rect 31404 7880 31432 7908
rect 33778 7896 33784 7948
rect 33836 7936 33842 7948
rect 33873 7939 33931 7945
rect 33873 7936 33885 7939
rect 33836 7908 33885 7936
rect 33836 7896 33842 7908
rect 33873 7905 33885 7908
rect 33919 7905 33931 7939
rect 33873 7899 33931 7905
rect 28721 7871 28779 7877
rect 28721 7868 28733 7871
rect 28684 7840 28733 7868
rect 28684 7828 28690 7840
rect 28721 7837 28733 7840
rect 28767 7837 28779 7871
rect 28721 7831 28779 7837
rect 29733 7871 29791 7877
rect 29733 7837 29745 7871
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 30193 7871 30251 7877
rect 30193 7837 30205 7871
rect 30239 7837 30251 7871
rect 30193 7831 30251 7837
rect 30561 7871 30619 7877
rect 30561 7837 30573 7871
rect 30607 7868 30619 7871
rect 30837 7871 30895 7877
rect 30837 7868 30849 7871
rect 30607 7840 30849 7868
rect 30607 7837 30619 7840
rect 30561 7831 30619 7837
rect 30837 7837 30849 7840
rect 30883 7868 30895 7871
rect 31297 7871 31355 7877
rect 31297 7868 31309 7871
rect 30883 7840 31309 7868
rect 30883 7837 30895 7840
rect 30837 7831 30895 7837
rect 31297 7837 31309 7840
rect 31343 7837 31355 7871
rect 31297 7831 31355 7837
rect 27154 7800 27160 7812
rect 27080 7772 27160 7800
rect 25004 7760 25010 7772
rect 27154 7760 27160 7772
rect 27212 7800 27218 7812
rect 29178 7800 29184 7812
rect 27212 7772 29184 7800
rect 27212 7760 27218 7772
rect 29178 7760 29184 7772
rect 29236 7760 29242 7812
rect 29748 7800 29776 7831
rect 31386 7828 31392 7880
rect 31444 7868 31450 7880
rect 31481 7871 31539 7877
rect 31481 7868 31493 7871
rect 31444 7840 31493 7868
rect 31444 7828 31450 7840
rect 31481 7837 31493 7840
rect 31527 7837 31539 7871
rect 31481 7831 31539 7837
rect 31754 7828 31760 7880
rect 31812 7828 31818 7880
rect 34256 7877 34284 7976
rect 36357 7973 36369 8007
rect 36403 8004 36415 8007
rect 36538 8004 36544 8016
rect 36403 7976 36544 8004
rect 36403 7973 36415 7976
rect 36357 7967 36415 7973
rect 36538 7964 36544 7976
rect 36596 7964 36602 8016
rect 36814 7964 36820 8016
rect 36872 7964 36878 8016
rect 34333 7939 34391 7945
rect 34333 7905 34345 7939
rect 34379 7936 34391 7939
rect 34422 7936 34428 7948
rect 34379 7908 34428 7936
rect 34379 7905 34391 7908
rect 34333 7899 34391 7905
rect 34422 7896 34428 7908
rect 34480 7896 34486 7948
rect 36832 7936 36860 7964
rect 35636 7908 36860 7936
rect 34241 7871 34299 7877
rect 34241 7837 34253 7871
rect 34287 7837 34299 7871
rect 34440 7868 34468 7896
rect 34701 7871 34759 7877
rect 34701 7868 34713 7871
rect 34440 7840 34713 7868
rect 34241 7831 34299 7837
rect 34701 7837 34713 7840
rect 34747 7837 34759 7871
rect 34701 7831 34759 7837
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 34885 7871 34943 7877
rect 34885 7868 34897 7871
rect 34848 7840 34897 7868
rect 34848 7828 34854 7840
rect 34885 7837 34897 7840
rect 34931 7837 34943 7871
rect 34885 7831 34943 7837
rect 35161 7871 35219 7877
rect 35161 7837 35173 7871
rect 35207 7868 35219 7871
rect 35250 7868 35256 7880
rect 35207 7840 35256 7868
rect 35207 7837 35219 7840
rect 35161 7831 35219 7837
rect 35250 7828 35256 7840
rect 35308 7828 35314 7880
rect 35636 7877 35664 7908
rect 35345 7871 35403 7877
rect 35345 7837 35357 7871
rect 35391 7868 35403 7871
rect 35621 7871 35679 7877
rect 35621 7868 35633 7871
rect 35391 7840 35633 7868
rect 35391 7837 35403 7840
rect 35345 7831 35403 7837
rect 35621 7837 35633 7840
rect 35667 7837 35679 7871
rect 36081 7871 36139 7877
rect 36081 7868 36093 7871
rect 35621 7831 35679 7837
rect 36004 7840 36093 7868
rect 30374 7800 30380 7812
rect 29748 7772 30380 7800
rect 30374 7760 30380 7772
rect 30432 7760 30438 7812
rect 35268 7800 35296 7828
rect 35437 7803 35495 7809
rect 35437 7800 35449 7803
rect 35268 7772 35449 7800
rect 35437 7769 35449 7772
rect 35483 7769 35495 7803
rect 35437 7763 35495 7769
rect 36004 7744 36032 7840
rect 36081 7837 36093 7840
rect 36127 7837 36139 7871
rect 36081 7831 36139 7837
rect 36262 7828 36268 7880
rect 36320 7868 36326 7880
rect 36357 7871 36415 7877
rect 36357 7868 36369 7871
rect 36320 7840 36369 7868
rect 36320 7828 36326 7840
rect 36357 7837 36369 7840
rect 36403 7837 36415 7871
rect 36357 7831 36415 7837
rect 36817 7871 36875 7877
rect 36817 7837 36829 7871
rect 36863 7837 36875 7871
rect 36924 7868 36952 8044
rect 37274 8032 37280 8084
rect 37332 8072 37338 8084
rect 37737 8075 37795 8081
rect 37737 8072 37749 8075
rect 37332 8044 37749 8072
rect 37332 8032 37338 8044
rect 37737 8041 37749 8044
rect 37783 8041 37795 8075
rect 37737 8035 37795 8041
rect 37001 7939 37059 7945
rect 37001 7905 37013 7939
rect 37047 7936 37059 7939
rect 37829 7939 37887 7945
rect 37047 7908 37596 7936
rect 37047 7905 37059 7908
rect 37001 7899 37059 7905
rect 36924 7840 37228 7868
rect 36817 7831 36875 7837
rect 36832 7800 36860 7831
rect 36998 7800 37004 7812
rect 36832 7772 37004 7800
rect 36998 7760 37004 7772
rect 37056 7760 37062 7812
rect 37200 7809 37228 7840
rect 37274 7828 37280 7880
rect 37332 7828 37338 7880
rect 37568 7877 37596 7908
rect 37829 7905 37841 7939
rect 37875 7936 37887 7939
rect 38470 7936 38476 7948
rect 37875 7908 38476 7936
rect 37875 7905 37887 7908
rect 37829 7899 37887 7905
rect 37553 7871 37611 7877
rect 37553 7837 37565 7871
rect 37599 7837 37611 7871
rect 37553 7831 37611 7837
rect 37185 7803 37243 7809
rect 37185 7769 37197 7803
rect 37231 7800 37243 7803
rect 37844 7800 37872 7899
rect 38470 7896 38476 7908
rect 38528 7896 38534 7948
rect 37918 7828 37924 7880
rect 37976 7828 37982 7880
rect 38197 7871 38255 7877
rect 38197 7868 38209 7871
rect 38120 7840 38209 7868
rect 37231 7772 37872 7800
rect 37231 7769 37243 7772
rect 37185 7763 37243 7769
rect 7340 7704 8984 7732
rect 7340 7692 7346 7704
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 11572 7704 12265 7732
rect 11572 7692 11578 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 16482 7692 16488 7744
rect 16540 7692 16546 7744
rect 16853 7735 16911 7741
rect 16853 7701 16865 7735
rect 16899 7732 16911 7735
rect 16942 7732 16948 7744
rect 16899 7704 16948 7732
rect 16899 7701 16911 7704
rect 16853 7695 16911 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 22094 7692 22100 7744
rect 22152 7692 22158 7744
rect 22189 7735 22247 7741
rect 22189 7701 22201 7735
rect 22235 7732 22247 7735
rect 22370 7732 22376 7744
rect 22235 7704 22376 7732
rect 22235 7701 22247 7704
rect 22189 7695 22247 7701
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 23290 7692 23296 7744
rect 23348 7732 23354 7744
rect 23569 7735 23627 7741
rect 23569 7732 23581 7735
rect 23348 7704 23581 7732
rect 23348 7692 23354 7704
rect 23569 7701 23581 7704
rect 23615 7701 23627 7735
rect 23569 7695 23627 7701
rect 24578 7692 24584 7744
rect 24636 7732 24642 7744
rect 25041 7735 25099 7741
rect 25041 7732 25053 7735
rect 24636 7704 25053 7732
rect 24636 7692 24642 7704
rect 25041 7701 25053 7704
rect 25087 7701 25099 7735
rect 25041 7695 25099 7701
rect 31938 7692 31944 7744
rect 31996 7692 32002 7744
rect 33502 7692 33508 7744
rect 33560 7732 33566 7744
rect 34701 7735 34759 7741
rect 34701 7732 34713 7735
rect 33560 7704 34713 7732
rect 33560 7692 33566 7704
rect 34701 7701 34713 7704
rect 34747 7701 34759 7735
rect 34701 7695 34759 7701
rect 35342 7692 35348 7744
rect 35400 7692 35406 7744
rect 35805 7735 35863 7741
rect 35805 7701 35817 7735
rect 35851 7732 35863 7735
rect 35986 7732 35992 7744
rect 35851 7704 35992 7732
rect 35851 7701 35863 7704
rect 35805 7695 35863 7701
rect 35986 7692 35992 7704
rect 36044 7692 36050 7744
rect 36078 7692 36084 7744
rect 36136 7732 36142 7744
rect 36173 7735 36231 7741
rect 36173 7732 36185 7735
rect 36136 7704 36185 7732
rect 36136 7692 36142 7704
rect 36173 7701 36185 7704
rect 36219 7701 36231 7735
rect 36173 7695 36231 7701
rect 37366 7692 37372 7744
rect 37424 7692 37430 7744
rect 38120 7741 38148 7840
rect 38197 7837 38209 7840
rect 38243 7837 38255 7871
rect 38197 7831 38255 7837
rect 38105 7735 38163 7741
rect 38105 7701 38117 7735
rect 38151 7701 38163 7735
rect 38105 7695 38163 7701
rect 38378 7692 38384 7744
rect 38436 7692 38442 7744
rect 1104 7642 38824 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 38824 7642
rect 1104 7568 38824 7590
rect 4706 7488 4712 7540
rect 4764 7488 4770 7540
rect 10318 7488 10324 7540
rect 10376 7488 10382 7540
rect 11146 7528 11152 7540
rect 10428 7500 11152 7528
rect 10428 7472 10456 7500
rect 11146 7488 11152 7500
rect 11204 7528 11210 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11204 7500 11529 7528
rect 11204 7488 11210 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 15654 7528 15660 7540
rect 11517 7491 11575 7497
rect 14752 7500 15660 7528
rect 2866 7420 2872 7472
rect 2924 7420 2930 7472
rect 9953 7463 10011 7469
rect 9953 7429 9965 7463
rect 9999 7429 10011 7463
rect 9953 7423 10011 7429
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4080 7364 4629 7392
rect 4080 7336 4108 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 842 7284 848 7336
rect 900 7324 906 7336
rect 1397 7327 1455 7333
rect 1397 7324 1409 7327
rect 900 7296 1409 7324
rect 900 7284 906 7296
rect 1397 7293 1409 7296
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 2590 7284 2596 7336
rect 2648 7284 2654 7336
rect 4062 7284 4068 7336
rect 4120 7284 4126 7336
rect 4632 7324 4660 7355
rect 4798 7352 4804 7404
rect 4856 7352 4862 7404
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5258 7392 5264 7404
rect 5123 7364 5264 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 4908 7324 4936 7355
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 7558 7352 7564 7404
rect 7616 7392 7622 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 7616 7364 8217 7392
rect 7616 7352 7622 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 9968 7392 9996 7423
rect 10134 7420 10140 7472
rect 10192 7469 10198 7472
rect 10192 7463 10211 7469
rect 10199 7429 10211 7463
rect 10192 7423 10211 7429
rect 10192 7420 10198 7423
rect 10410 7420 10416 7472
rect 10468 7420 10474 7472
rect 14752 7469 14780 7500
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 16390 7528 16396 7540
rect 16255 7500 16396 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16482 7488 16488 7540
rect 16540 7528 16546 7540
rect 17770 7528 17776 7540
rect 16540 7500 17776 7528
rect 16540 7488 16546 7500
rect 17770 7488 17776 7500
rect 17828 7528 17834 7540
rect 18417 7531 18475 7537
rect 18417 7528 18429 7531
rect 17828 7500 18429 7528
rect 17828 7488 17834 7500
rect 18417 7497 18429 7500
rect 18463 7497 18475 7531
rect 18417 7491 18475 7497
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 22738 7528 22744 7540
rect 21416 7500 22744 7528
rect 21416 7488 21422 7500
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 24210 7528 24216 7540
rect 22848 7500 24216 7528
rect 14737 7463 14795 7469
rect 14737 7429 14749 7463
rect 14783 7429 14795 7463
rect 14737 7423 14795 7429
rect 15194 7420 15200 7472
rect 15252 7420 15258 7472
rect 16942 7420 16948 7472
rect 17000 7420 17006 7472
rect 18230 7460 18236 7472
rect 18170 7432 18236 7460
rect 18230 7420 18236 7432
rect 18288 7460 18294 7472
rect 19978 7460 19984 7472
rect 18288 7432 19984 7460
rect 18288 7420 18294 7432
rect 19978 7420 19984 7432
rect 20036 7420 20042 7472
rect 22557 7463 22615 7469
rect 22557 7460 22569 7463
rect 20916 7432 22569 7460
rect 11330 7392 11336 7404
rect 9968 7364 11336 7392
rect 8205 7355 8263 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 20916 7401 20944 7432
rect 22557 7429 22569 7432
rect 22603 7429 22615 7463
rect 22557 7423 22615 7429
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 21174 7352 21180 7404
rect 21232 7352 21238 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21407 7364 21833 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22848 7401 22876 7500
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 25038 7528 25044 7540
rect 24596 7500 25044 7528
rect 23290 7460 23296 7472
rect 23032 7432 23296 7460
rect 22833 7395 22891 7401
rect 22833 7392 22845 7395
rect 22152 7364 22845 7392
rect 22152 7352 22158 7364
rect 22833 7361 22845 7364
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 22922 7352 22928 7404
rect 22980 7352 22986 7404
rect 23032 7401 23060 7432
rect 23290 7420 23296 7432
rect 23348 7420 23354 7472
rect 24228 7401 24256 7488
rect 24596 7460 24624 7500
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 25130 7488 25136 7540
rect 25188 7488 25194 7540
rect 26786 7488 26792 7540
rect 26844 7528 26850 7540
rect 26973 7531 27031 7537
rect 26973 7528 26985 7531
rect 26844 7500 26985 7528
rect 26844 7488 26850 7500
rect 26973 7497 26985 7500
rect 27019 7497 27031 7531
rect 26973 7491 27031 7497
rect 27338 7488 27344 7540
rect 27396 7528 27402 7540
rect 27433 7531 27491 7537
rect 27433 7528 27445 7531
rect 27396 7500 27445 7528
rect 27396 7488 27402 7500
rect 27433 7497 27445 7500
rect 27479 7497 27491 7531
rect 27433 7491 27491 7497
rect 36817 7531 36875 7537
rect 36817 7497 36829 7531
rect 36863 7528 36875 7531
rect 37918 7528 37924 7540
rect 36863 7500 37924 7528
rect 36863 7497 36875 7500
rect 36817 7491 36875 7497
rect 37918 7488 37924 7500
rect 37976 7488 37982 7540
rect 25148 7460 25176 7488
rect 24320 7432 24624 7460
rect 24688 7432 25176 7460
rect 27157 7463 27215 7469
rect 24320 7401 24348 7432
rect 23017 7395 23075 7401
rect 23017 7361 23029 7395
rect 23063 7361 23075 7395
rect 23017 7355 23075 7361
rect 23201 7395 23259 7401
rect 23201 7361 23213 7395
rect 23247 7361 23259 7395
rect 23201 7355 23259 7361
rect 24029 7395 24087 7401
rect 24029 7361 24041 7395
rect 24075 7392 24087 7395
rect 24213 7395 24271 7401
rect 24075 7364 24164 7392
rect 24075 7361 24087 7364
rect 24029 7355 24087 7361
rect 4632 7296 4936 7324
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7324 8447 7327
rect 8570 7324 8576 7336
rect 8435 7296 8576 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 11054 7324 11060 7336
rect 10560 7296 11060 7324
rect 10560 7284 10566 7296
rect 11054 7284 11060 7296
rect 11112 7324 11118 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 11112 7296 11161 7324
rect 11112 7284 11118 7296
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 21192 7256 21220 7352
rect 21450 7284 21456 7336
rect 21508 7324 21514 7336
rect 21634 7324 21640 7336
rect 21508 7296 21640 7324
rect 21508 7284 21514 7296
rect 21634 7284 21640 7296
rect 21692 7324 21698 7336
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 21692 7296 22385 7324
rect 21692 7284 21698 7296
rect 22373 7293 22385 7296
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 21726 7256 21732 7268
rect 21192 7228 21732 7256
rect 21726 7216 21732 7228
rect 21784 7256 21790 7268
rect 23216 7256 23244 7355
rect 23290 7256 23296 7268
rect 21784 7228 23296 7256
rect 21784 7216 21790 7228
rect 23290 7216 23296 7228
rect 23348 7216 23354 7268
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4430 7188 4436 7200
rect 4387 7160 4436 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4430 7148 4436 7160
rect 4488 7188 4494 7200
rect 4798 7188 4804 7200
rect 4488 7160 4804 7188
rect 4488 7148 4494 7160
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 4890 7148 4896 7200
rect 4948 7148 4954 7200
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7800 7160 8033 7188
rect 7800 7148 7806 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 10137 7191 10195 7197
rect 10137 7157 10149 7191
rect 10183 7188 10195 7191
rect 10778 7188 10784 7200
rect 10183 7160 10784 7188
rect 10183 7157 10195 7160
rect 10137 7151 10195 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 20714 7148 20720 7200
rect 20772 7148 20778 7200
rect 23842 7148 23848 7200
rect 23900 7148 23906 7200
rect 24136 7188 24164 7364
rect 24213 7361 24225 7395
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 24412 7324 24440 7355
rect 24578 7352 24584 7404
rect 24636 7352 24642 7404
rect 24688 7401 24716 7432
rect 27157 7429 27169 7463
rect 27203 7460 27215 7463
rect 36998 7460 37004 7472
rect 27203 7432 27476 7460
rect 27203 7429 27215 7432
rect 27157 7423 27215 7429
rect 24673 7395 24731 7401
rect 24673 7361 24685 7395
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24762 7352 24768 7404
rect 24820 7392 24826 7404
rect 24820 7364 24865 7392
rect 24820 7352 24826 7364
rect 24946 7352 24952 7404
rect 25004 7352 25010 7404
rect 25038 7352 25044 7404
rect 25096 7352 25102 7404
rect 25130 7352 25136 7404
rect 25188 7401 25194 7404
rect 27448 7401 27476 7432
rect 36372 7432 37004 7460
rect 25188 7355 25196 7401
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7361 27399 7395
rect 27341 7355 27399 7361
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7392 27491 7395
rect 27522 7392 27528 7404
rect 27479 7364 27528 7392
rect 27479 7361 27491 7364
rect 27433 7355 27491 7361
rect 25188 7352 25194 7355
rect 27356 7324 27384 7355
rect 27522 7352 27528 7364
rect 27580 7352 27586 7404
rect 27617 7395 27675 7401
rect 27617 7361 27629 7395
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 27632 7324 27660 7355
rect 32306 7352 32312 7404
rect 32364 7352 32370 7404
rect 32769 7395 32827 7401
rect 32769 7392 32781 7395
rect 32692 7364 32781 7392
rect 24412 7296 24716 7324
rect 27356 7296 27660 7324
rect 24688 7268 24716 7296
rect 27448 7268 27476 7296
rect 31938 7284 31944 7336
rect 31996 7324 32002 7336
rect 32217 7327 32275 7333
rect 32217 7324 32229 7327
rect 31996 7296 32229 7324
rect 31996 7284 32002 7296
rect 32217 7293 32229 7296
rect 32263 7293 32275 7327
rect 32217 7287 32275 7293
rect 32692 7268 32720 7364
rect 32769 7361 32781 7364
rect 32815 7361 32827 7395
rect 32769 7355 32827 7361
rect 32950 7352 32956 7404
rect 33008 7352 33014 7404
rect 33134 7352 33140 7404
rect 33192 7352 33198 7404
rect 33321 7395 33379 7401
rect 33321 7361 33333 7395
rect 33367 7361 33379 7395
rect 33321 7355 33379 7361
rect 32861 7327 32919 7333
rect 32861 7293 32873 7327
rect 32907 7324 32919 7327
rect 33336 7324 33364 7355
rect 33410 7352 33416 7404
rect 33468 7352 33474 7404
rect 33502 7352 33508 7404
rect 33560 7352 33566 7404
rect 33686 7352 33692 7404
rect 33744 7352 33750 7404
rect 35713 7395 35771 7401
rect 35713 7361 35725 7395
rect 35759 7392 35771 7395
rect 36078 7392 36084 7404
rect 35759 7364 36084 7392
rect 35759 7361 35771 7364
rect 35713 7355 35771 7361
rect 36078 7352 36084 7364
rect 36136 7352 36142 7404
rect 36170 7352 36176 7404
rect 36228 7352 36234 7404
rect 36372 7401 36400 7432
rect 36998 7420 37004 7432
rect 37056 7420 37062 7472
rect 36357 7395 36415 7401
rect 36357 7361 36369 7395
rect 36403 7361 36415 7395
rect 36357 7355 36415 7361
rect 36446 7352 36452 7404
rect 36504 7352 36510 7404
rect 36538 7352 36544 7404
rect 36596 7352 36602 7404
rect 32907 7296 33364 7324
rect 32907 7293 32919 7296
rect 32861 7287 32919 7293
rect 35802 7284 35808 7336
rect 35860 7284 35866 7336
rect 24670 7216 24676 7268
rect 24728 7216 24734 7268
rect 27430 7216 27436 7268
rect 27488 7216 27494 7268
rect 32674 7216 32680 7268
rect 32732 7216 32738 7268
rect 24946 7188 24952 7200
rect 24136 7160 24952 7188
rect 24946 7148 24952 7160
rect 25004 7148 25010 7200
rect 25317 7191 25375 7197
rect 25317 7157 25329 7191
rect 25363 7188 25375 7191
rect 25498 7188 25504 7200
rect 25363 7160 25504 7188
rect 25363 7157 25375 7160
rect 25317 7151 25375 7157
rect 25498 7148 25504 7160
rect 25556 7148 25562 7200
rect 33410 7148 33416 7200
rect 33468 7188 33474 7200
rect 33873 7191 33931 7197
rect 33873 7188 33885 7191
rect 33468 7160 33885 7188
rect 33468 7148 33474 7160
rect 33873 7157 33885 7160
rect 33919 7157 33931 7191
rect 33873 7151 33931 7157
rect 35437 7191 35495 7197
rect 35437 7157 35449 7191
rect 35483 7188 35495 7191
rect 35710 7188 35716 7200
rect 35483 7160 35716 7188
rect 35483 7157 35495 7160
rect 35437 7151 35495 7157
rect 35710 7148 35716 7160
rect 35768 7148 35774 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 3970 6984 3976 6996
rect 3467 6956 3976 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 5457 6987 5515 6993
rect 5457 6984 5469 6987
rect 4948 6956 5469 6984
rect 4948 6944 4954 6956
rect 5457 6953 5469 6956
rect 5503 6953 5515 6987
rect 5457 6947 5515 6953
rect 6444 6987 6502 6993
rect 6444 6953 6456 6987
rect 6490 6984 6502 6987
rect 7190 6984 7196 6996
rect 6490 6956 7196 6984
rect 6490 6953 6502 6956
rect 6444 6947 6502 6953
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 19968 6987 20026 6993
rect 19968 6953 19980 6987
rect 20014 6984 20026 6987
rect 20714 6984 20720 6996
rect 20014 6956 20720 6984
rect 20014 6953 20026 6956
rect 19968 6947 20026 6953
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 21450 6944 21456 6996
rect 21508 6944 21514 6996
rect 27798 6944 27804 6996
rect 27856 6944 27862 6996
rect 30374 6944 30380 6996
rect 30432 6944 30438 6996
rect 36712 6987 36770 6993
rect 36712 6953 36724 6987
rect 36758 6984 36770 6987
rect 37366 6984 37372 6996
rect 36758 6956 37372 6984
rect 36758 6953 36770 6956
rect 36712 6947 36770 6953
rect 37366 6944 37372 6956
rect 37424 6944 37430 6996
rect 3605 6919 3663 6925
rect 3605 6885 3617 6919
rect 3651 6916 3663 6919
rect 4062 6916 4068 6928
rect 3651 6888 4068 6916
rect 3651 6885 3663 6888
rect 3605 6879 3663 6885
rect 4062 6876 4068 6888
rect 4120 6876 4126 6928
rect 15194 6916 15200 6928
rect 15120 6888 15200 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2682 6848 2688 6860
rect 1443 6820 2688 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2682 6808 2688 6820
rect 2740 6848 2746 6860
rect 4154 6848 4160 6860
rect 2740 6820 4160 6848
rect 2740 6808 2746 6820
rect 4154 6808 4160 6820
rect 4212 6848 4218 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 4212 6820 5733 6848
rect 4212 6808 4218 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 6227 6820 8953 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 8941 6817 8953 6820
rect 8987 6848 8999 6851
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 8987 6820 12173 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 3142 6780 3148 6792
rect 2806 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6780 3206 6792
rect 3200 6752 3832 6780
rect 3200 6740 3206 6752
rect 3804 6724 3832 6752
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 1670 6672 1676 6724
rect 1728 6672 1734 6724
rect 3234 6672 3240 6724
rect 3292 6672 3298 6724
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 7834 6712 7840 6724
rect 3844 6684 4278 6712
rect 7682 6684 7840 6712
rect 3844 6672 3850 6684
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 8588 6712 8616 6740
rect 7944 6684 8616 6712
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3252 6644 3280 6672
rect 3191 6616 3280 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 3447 6647 3505 6653
rect 3447 6644 3459 6647
rect 3384 6616 3459 6644
rect 3384 6604 3390 6616
rect 3447 6613 3459 6616
rect 3493 6644 3505 6647
rect 5534 6644 5540 6656
rect 3493 6616 5540 6644
rect 3493 6613 3505 6616
rect 3447 6607 3505 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 7944 6653 7972 6684
rect 9214 6672 9220 6724
rect 9272 6672 9278 6724
rect 9766 6672 9772 6724
rect 9824 6672 9830 6724
rect 10888 6721 10916 6820
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13446 6848 13452 6860
rect 12952 6820 13452 6848
rect 12952 6808 12958 6820
rect 13446 6808 13452 6820
rect 13504 6848 13510 6860
rect 15120 6848 15148 6888
rect 15194 6876 15200 6888
rect 15252 6876 15258 6928
rect 13504 6820 15148 6848
rect 13504 6808 13510 6820
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 26237 6851 26295 6857
rect 26237 6848 26249 6851
rect 21048 6820 21312 6848
rect 21048 6808 21054 6820
rect 11330 6740 11336 6792
rect 11388 6740 11394 6792
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11698 6740 11704 6792
rect 11756 6740 11762 6792
rect 11790 6740 11796 6792
rect 11848 6740 11854 6792
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 13924 6752 14657 6780
rect 10873 6715 10931 6721
rect 10873 6681 10885 6715
rect 10919 6712 10931 6715
rect 11054 6712 11060 6724
rect 10919 6684 11060 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 11716 6712 11744 6740
rect 12066 6712 12072 6724
rect 11716 6684 12072 6712
rect 12066 6672 12072 6684
rect 12124 6672 12130 6724
rect 12434 6672 12440 6724
rect 12492 6672 12498 6724
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 12894 6712 12900 6724
rect 12768 6684 12900 6712
rect 12768 6672 12774 6684
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8018 6604 8024 6656
rect 8076 6604 8082 6656
rect 10502 6604 10508 6656
rect 10560 6644 10566 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10560 6616 10701 6644
rect 10560 6604 10566 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 13924 6653 13952 6752
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 16632 6752 17693 6780
rect 16632 6740 16638 6752
rect 17681 6749 17693 6752
rect 17727 6780 17739 6783
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 17727 6752 17785 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 17773 6749 17785 6752
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 18506 6672 18512 6724
rect 18564 6712 18570 6724
rect 19610 6712 19616 6724
rect 18564 6684 19616 6712
rect 18564 6672 18570 6684
rect 19610 6672 19616 6684
rect 19668 6712 19674 6724
rect 19720 6712 19748 6743
rect 21284 6712 21312 6820
rect 25884 6820 26249 6848
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 23474 6780 23480 6792
rect 22879 6752 23480 6780
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 23474 6740 23480 6752
rect 23532 6740 23538 6792
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6780 24915 6783
rect 25130 6780 25136 6792
rect 24903 6752 25136 6780
rect 24903 6749 24915 6752
rect 24857 6743 24915 6749
rect 25130 6740 25136 6752
rect 25188 6780 25194 6792
rect 25884 6789 25912 6820
rect 26237 6817 26249 6820
rect 26283 6817 26295 6851
rect 26237 6811 26295 6817
rect 27246 6808 27252 6860
rect 27304 6848 27310 6860
rect 27433 6851 27491 6857
rect 27433 6848 27445 6851
rect 27304 6820 27445 6848
rect 27304 6808 27310 6820
rect 27433 6817 27445 6820
rect 27479 6817 27491 6851
rect 32769 6851 32827 6857
rect 27433 6811 27491 6817
rect 29288 6820 29776 6848
rect 29288 6792 29316 6820
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 25188 6752 25697 6780
rect 25188 6740 25194 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 25869 6783 25927 6789
rect 25869 6749 25881 6783
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 26050 6740 26056 6792
rect 26108 6740 26114 6792
rect 26142 6740 26148 6792
rect 26200 6740 26206 6792
rect 26329 6783 26387 6789
rect 26329 6749 26341 6783
rect 26375 6749 26387 6783
rect 26329 6743 26387 6749
rect 27525 6783 27583 6789
rect 27525 6749 27537 6783
rect 27571 6749 27583 6783
rect 27525 6743 27583 6749
rect 21358 6712 21364 6724
rect 19668 6684 19748 6712
rect 21206 6684 21364 6712
rect 19668 6672 19674 6684
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 25406 6672 25412 6724
rect 25464 6712 25470 6724
rect 26344 6712 26372 6743
rect 25464 6684 26372 6712
rect 25464 6672 25470 6684
rect 27430 6672 27436 6724
rect 27488 6712 27494 6724
rect 27540 6712 27568 6743
rect 29086 6740 29092 6792
rect 29144 6740 29150 6792
rect 29270 6740 29276 6792
rect 29328 6740 29334 6792
rect 29748 6789 29776 6820
rect 32769 6817 32781 6851
rect 32815 6848 32827 6851
rect 33134 6848 33140 6860
rect 32815 6820 33140 6848
rect 32815 6817 32827 6820
rect 32769 6811 32827 6817
rect 33134 6808 33140 6820
rect 33192 6808 33198 6860
rect 34701 6851 34759 6857
rect 34701 6848 34713 6851
rect 33796 6820 34713 6848
rect 33796 6792 33824 6820
rect 34701 6817 34713 6820
rect 34747 6817 34759 6851
rect 34701 6811 34759 6817
rect 35802 6808 35808 6860
rect 35860 6808 35866 6860
rect 36354 6808 36360 6860
rect 36412 6848 36418 6860
rect 36449 6851 36507 6857
rect 36449 6848 36461 6851
rect 36412 6820 36461 6848
rect 36412 6808 36418 6820
rect 36449 6817 36461 6820
rect 36495 6817 36507 6851
rect 36449 6811 36507 6817
rect 38470 6808 38476 6860
rect 38528 6808 38534 6860
rect 29549 6783 29607 6789
rect 29549 6749 29561 6783
rect 29595 6749 29607 6783
rect 29549 6743 29607 6749
rect 29733 6783 29791 6789
rect 29733 6749 29745 6783
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 27488 6684 27568 6712
rect 29104 6712 29132 6740
rect 29564 6712 29592 6743
rect 31938 6740 31944 6792
rect 31996 6780 32002 6792
rect 32125 6783 32183 6789
rect 32125 6780 32137 6783
rect 31996 6752 32137 6780
rect 31996 6740 32002 6752
rect 32125 6749 32137 6752
rect 32171 6749 32183 6783
rect 32125 6743 32183 6749
rect 32674 6740 32680 6792
rect 32732 6740 32738 6792
rect 32861 6783 32919 6789
rect 32861 6749 32873 6783
rect 32907 6780 32919 6783
rect 32950 6780 32956 6792
rect 32907 6752 32956 6780
rect 32907 6749 32919 6752
rect 32861 6743 32919 6749
rect 32950 6740 32956 6752
rect 33008 6740 33014 6792
rect 33410 6740 33416 6792
rect 33468 6740 33474 6792
rect 33502 6740 33508 6792
rect 33560 6780 33566 6792
rect 33560 6752 33605 6780
rect 33560 6740 33566 6752
rect 33778 6740 33784 6792
rect 33836 6740 33842 6792
rect 33870 6740 33876 6792
rect 33928 6789 33934 6792
rect 33928 6783 33977 6789
rect 33928 6749 33931 6783
rect 33965 6780 33977 6783
rect 34793 6783 34851 6789
rect 34793 6780 34805 6783
rect 33965 6752 34805 6780
rect 33965 6749 33977 6752
rect 33928 6743 33977 6749
rect 34793 6749 34805 6752
rect 34839 6749 34851 6783
rect 34793 6743 34851 6749
rect 34977 6783 35035 6789
rect 34977 6749 34989 6783
rect 35023 6749 35035 6783
rect 34977 6743 35035 6749
rect 33928 6740 33934 6743
rect 29104 6684 29592 6712
rect 29917 6715 29975 6721
rect 27488 6672 27494 6684
rect 29917 6681 29929 6715
rect 29963 6712 29975 6715
rect 30009 6715 30067 6721
rect 30009 6712 30021 6715
rect 29963 6684 30021 6712
rect 29963 6681 29975 6684
rect 29917 6675 29975 6681
rect 30009 6681 30021 6684
rect 30055 6681 30067 6715
rect 30009 6675 30067 6681
rect 30193 6715 30251 6721
rect 30193 6681 30205 6715
rect 30239 6681 30251 6715
rect 30193 6675 30251 6681
rect 13909 6647 13967 6653
rect 13909 6644 13921 6647
rect 12216 6616 13921 6644
rect 12216 6604 12222 6616
rect 13909 6613 13921 6616
rect 13955 6613 13967 6647
rect 13909 6607 13967 6613
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 22554 6604 22560 6656
rect 22612 6644 22618 6656
rect 22741 6647 22799 6653
rect 22741 6644 22753 6647
rect 22612 6616 22753 6644
rect 22612 6604 22618 6616
rect 22741 6613 22753 6616
rect 22787 6613 22799 6647
rect 22741 6607 22799 6613
rect 24394 6604 24400 6656
rect 24452 6644 24458 6656
rect 24765 6647 24823 6653
rect 24765 6644 24777 6647
rect 24452 6616 24777 6644
rect 24452 6604 24458 6616
rect 24765 6613 24777 6616
rect 24811 6613 24823 6647
rect 24765 6607 24823 6613
rect 29181 6647 29239 6653
rect 29181 6613 29193 6647
rect 29227 6644 29239 6647
rect 29362 6644 29368 6656
rect 29227 6616 29368 6644
rect 29227 6613 29239 6616
rect 29181 6607 29239 6613
rect 29362 6604 29368 6616
rect 29420 6644 29426 6656
rect 30208 6644 30236 6675
rect 32306 6672 32312 6724
rect 32364 6672 32370 6724
rect 33318 6672 33324 6724
rect 33376 6712 33382 6724
rect 33686 6712 33692 6724
rect 33376 6684 33692 6712
rect 33376 6672 33382 6684
rect 33686 6672 33692 6684
rect 33744 6672 33750 6724
rect 34992 6712 35020 6743
rect 35342 6740 35348 6792
rect 35400 6780 35406 6792
rect 35621 6783 35679 6789
rect 35621 6780 35633 6783
rect 35400 6752 35633 6780
rect 35400 6740 35406 6752
rect 35621 6749 35633 6752
rect 35667 6749 35679 6783
rect 35621 6743 35679 6749
rect 34072 6684 35020 6712
rect 29420 6616 30236 6644
rect 29420 6604 29426 6616
rect 32398 6604 32404 6656
rect 32456 6644 32462 6656
rect 34072 6653 34100 6684
rect 37458 6672 37464 6724
rect 37516 6672 37522 6724
rect 32493 6647 32551 6653
rect 32493 6644 32505 6647
rect 32456 6616 32505 6644
rect 32456 6604 32462 6616
rect 32493 6613 32505 6616
rect 32539 6613 32551 6647
rect 32493 6607 32551 6613
rect 34057 6647 34115 6653
rect 34057 6613 34069 6647
rect 34103 6613 34115 6647
rect 34057 6607 34115 6613
rect 34790 6604 34796 6656
rect 34848 6644 34854 6656
rect 35161 6647 35219 6653
rect 35161 6644 35173 6647
rect 34848 6616 35173 6644
rect 34848 6604 34854 6616
rect 35161 6613 35173 6616
rect 35207 6613 35219 6647
rect 35161 6607 35219 6613
rect 35434 6604 35440 6656
rect 35492 6604 35498 6656
rect 1104 6554 38824 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 38824 6554
rect 1104 6480 38824 6502
rect 7190 6400 7196 6452
rect 7248 6400 7254 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8021 6443 8079 6449
rect 7800 6412 7972 6440
rect 7800 6400 7806 6412
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6372 4675 6375
rect 5261 6375 5319 6381
rect 5261 6372 5273 6375
rect 4663 6344 5273 6372
rect 4663 6341 4675 6344
rect 4617 6335 4675 6341
rect 5261 6341 5273 6344
rect 5307 6341 5319 6375
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 5261 6335 5319 6341
rect 7392 6344 7849 6372
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2731 6276 2973 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 3326 6304 3332 6316
rect 2961 6267 3019 6273
rect 3160 6276 3332 6304
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 1728 6208 2329 6236
rect 1728 6196 1734 6208
rect 2317 6205 2329 6208
rect 2363 6205 2375 6239
rect 2317 6199 2375 6205
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 2866 6236 2872 6248
rect 2823 6208 2872 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 2866 6196 2872 6208
rect 2924 6236 2930 6248
rect 3160 6236 3188 6276
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4709 6307 4767 6313
rect 4709 6304 4721 6307
rect 4028 6276 4721 6304
rect 4028 6264 4034 6276
rect 4709 6273 4721 6276
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 5031 6276 5457 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 2924 6208 3188 6236
rect 2924 6196 2930 6208
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3605 6239 3663 6245
rect 3605 6236 3617 6239
rect 3292 6208 3617 6236
rect 3292 6196 3298 6208
rect 3605 6205 3617 6208
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 3620 6168 3648 6199
rect 4798 6196 4804 6248
rect 4856 6196 4862 6248
rect 5000 6168 5028 6267
rect 5534 6264 5540 6316
rect 5592 6264 5598 6316
rect 7392 6313 7420 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 7944 6372 7972 6412
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 9214 6440 9220 6452
rect 8067 6412 9220 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10321 6443 10379 6449
rect 10008 6412 10272 6440
rect 10008 6400 10014 6412
rect 10134 6372 10140 6384
rect 7944 6344 8432 6372
rect 7837 6335 7895 6341
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8110 6304 8116 6316
rect 7975 6276 8116 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8404 6313 8432 6344
rect 8680 6344 10140 6372
rect 8680 6313 8708 6344
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 10244 6372 10272 6412
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10870 6440 10876 6452
rect 10367 6412 10876 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 10870 6400 10876 6412
rect 10928 6440 10934 6452
rect 11698 6440 11704 6452
rect 10928 6412 11704 6440
rect 10928 6400 10934 6412
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 11992 6412 12480 6440
rect 10689 6375 10747 6381
rect 10689 6372 10701 6375
rect 10244 6344 10701 6372
rect 10689 6341 10701 6344
rect 10735 6372 10747 6375
rect 11790 6372 11796 6384
rect 10735 6344 11796 6372
rect 10735 6341 10747 6344
rect 10689 6335 10747 6341
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 8018 6236 8024 6248
rect 7699 6208 8024 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8312 6236 8340 6267
rect 8496 6236 8524 6267
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 10502 6304 10508 6316
rect 10152 6276 10508 6304
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8312 6208 8432 6236
rect 8496 6208 8861 6236
rect 3620 6140 5028 6168
rect 5258 6128 5264 6180
rect 5316 6128 5322 6180
rect 8294 6168 8300 6180
rect 8128 6140 8300 6168
rect 4706 6060 4712 6112
rect 4764 6060 4770 6112
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 8128 6100 8156 6140
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 8404 6168 8432 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 10152 6245 10180 6276
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 11256 6313 11284 6344
rect 11790 6332 11796 6344
rect 11848 6332 11854 6384
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6302 11023 6307
rect 11241 6307 11299 6313
rect 11011 6274 11100 6302
rect 11011 6273 11023 6274
rect 10965 6267 11023 6273
rect 10112 6239 10180 6245
rect 10112 6236 10124 6239
rect 9180 6208 10124 6236
rect 9180 6196 9186 6208
rect 10112 6205 10124 6208
rect 10158 6208 10180 6239
rect 10229 6239 10287 6245
rect 10158 6205 10170 6208
rect 10112 6199 10170 6205
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6236 10655 6239
rect 11072 6236 11100 6274
rect 11241 6273 11253 6307
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 11514 6264 11520 6316
rect 11572 6304 11578 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11572 6276 11713 6304
rect 11572 6264 11578 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 11992 6304 12020 6412
rect 12066 6332 12072 6384
rect 12124 6372 12130 6384
rect 12452 6381 12480 6412
rect 23014 6400 23020 6452
rect 23072 6440 23078 6452
rect 23201 6443 23259 6449
rect 23201 6440 23213 6443
rect 23072 6412 23213 6440
rect 23072 6400 23078 6412
rect 23201 6409 23213 6412
rect 23247 6409 23259 6443
rect 23201 6403 23259 6409
rect 23474 6400 23480 6452
rect 23532 6400 23538 6452
rect 24394 6400 24400 6452
rect 24452 6400 24458 6452
rect 24486 6400 24492 6452
rect 24544 6440 24550 6452
rect 24544 6412 25268 6440
rect 24544 6400 24550 6412
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 12124 6344 12173 6372
rect 12124 6332 12130 6344
rect 12161 6341 12173 6344
rect 12207 6341 12219 6375
rect 12161 6335 12219 6341
rect 12437 6375 12495 6381
rect 12437 6341 12449 6375
rect 12483 6372 12495 6375
rect 12526 6372 12532 6384
rect 12483 6344 12532 6372
rect 12483 6341 12495 6344
rect 12437 6335 12495 6341
rect 12526 6332 12532 6344
rect 12584 6372 12590 6384
rect 13265 6375 13323 6381
rect 13265 6372 13277 6375
rect 12584 6344 13277 6372
rect 12584 6332 12590 6344
rect 13265 6341 13277 6344
rect 13311 6341 13323 6375
rect 13265 6335 13323 6341
rect 22925 6375 22983 6381
rect 22925 6341 22937 6375
rect 22971 6372 22983 6375
rect 23492 6372 23520 6400
rect 24670 6372 24676 6384
rect 22971 6344 24676 6372
rect 22971 6341 22983 6344
rect 22925 6335 22983 6341
rect 24670 6332 24676 6344
rect 24728 6332 24734 6384
rect 25240 6316 25268 6412
rect 26050 6400 26056 6452
rect 26108 6440 26114 6452
rect 26145 6443 26203 6449
rect 26145 6440 26157 6443
rect 26108 6412 26157 6440
rect 26108 6400 26114 6412
rect 26145 6409 26157 6412
rect 26191 6409 26203 6443
rect 26145 6403 26203 6409
rect 27246 6400 27252 6452
rect 27304 6400 27310 6452
rect 28813 6443 28871 6449
rect 28813 6409 28825 6443
rect 28859 6440 28871 6443
rect 29270 6440 29276 6452
rect 28859 6412 29276 6440
rect 28859 6409 28871 6412
rect 28813 6403 28871 6409
rect 29270 6400 29276 6412
rect 29328 6400 29334 6452
rect 30837 6443 30895 6449
rect 30837 6409 30849 6443
rect 30883 6440 30895 6443
rect 30883 6412 31432 6440
rect 30883 6409 30895 6412
rect 30837 6403 30895 6409
rect 25406 6332 25412 6384
rect 25464 6372 25470 6384
rect 25777 6375 25835 6381
rect 25777 6372 25789 6375
rect 25464 6344 25789 6372
rect 25464 6332 25470 6344
rect 25777 6341 25789 6344
rect 25823 6372 25835 6375
rect 25823 6344 26648 6372
rect 25823 6341 25835 6344
rect 25777 6335 25835 6341
rect 11931 6276 12020 6304
rect 12345 6307 12403 6313
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12345 6273 12357 6307
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 12667 6276 12725 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 12713 6273 12725 6276
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 11532 6236 11560 6264
rect 10643 6208 11560 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 9140 6168 9168 6196
rect 8404 6140 9168 6168
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 10244 6168 10272 6199
rect 9364 6140 10272 6168
rect 9364 6128 9370 6140
rect 10778 6128 10784 6180
rect 10836 6168 10842 6180
rect 12250 6168 12256 6180
rect 10836 6140 12256 6168
rect 10836 6128 10842 6140
rect 12250 6128 12256 6140
rect 12308 6168 12314 6180
rect 12360 6168 12388 6267
rect 12802 6264 12808 6316
rect 12860 6304 12866 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12860 6276 12909 6304
rect 12860 6264 12866 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 13044 6276 13093 6304
rect 13044 6264 13050 6276
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 14090 6304 14096 6316
rect 13403 6276 14096 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 16666 6264 16672 6316
rect 16724 6304 16730 6316
rect 17957 6307 18015 6313
rect 17957 6304 17969 6307
rect 16724 6276 17969 6304
rect 16724 6264 16730 6276
rect 17957 6273 17969 6276
rect 18003 6304 18015 6307
rect 18506 6304 18512 6316
rect 18003 6276 18512 6304
rect 18003 6273 18015 6276
rect 17957 6267 18015 6273
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 22002 6264 22008 6316
rect 22060 6304 22066 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 22060 6276 22109 6304
rect 22060 6264 22066 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6273 23351 6307
rect 23293 6267 23351 6273
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6304 23535 6307
rect 24210 6304 24216 6316
rect 23523 6276 24216 6304
rect 23523 6273 23535 6276
rect 23477 6267 23535 6273
rect 22278 6196 22284 6248
rect 22336 6196 22342 6248
rect 23198 6196 23204 6248
rect 23256 6236 23262 6248
rect 23308 6236 23336 6267
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 24305 6307 24363 6313
rect 24305 6273 24317 6307
rect 24351 6304 24363 6307
rect 24854 6304 24860 6316
rect 24351 6276 24860 6304
rect 24351 6273 24363 6276
rect 24305 6267 24363 6273
rect 24854 6264 24860 6276
rect 24912 6304 24918 6316
rect 24949 6307 25007 6313
rect 24949 6304 24961 6307
rect 24912 6276 24961 6304
rect 24912 6264 24918 6276
rect 24949 6273 24961 6276
rect 24995 6304 25007 6307
rect 25038 6304 25044 6316
rect 24995 6276 25044 6304
rect 24995 6273 25007 6276
rect 24949 6267 25007 6273
rect 25038 6264 25044 6276
rect 25096 6264 25102 6316
rect 25130 6264 25136 6316
rect 25188 6264 25194 6316
rect 25222 6264 25228 6316
rect 25280 6264 25286 6316
rect 25314 6264 25320 6316
rect 25372 6264 25378 6316
rect 25498 6264 25504 6316
rect 25556 6264 25562 6316
rect 25958 6264 25964 6316
rect 26016 6304 26022 6316
rect 26142 6304 26148 6316
rect 26016 6276 26148 6304
rect 26016 6264 26022 6276
rect 26142 6264 26148 6276
rect 26200 6264 26206 6316
rect 26620 6313 26648 6344
rect 27430 6332 27436 6384
rect 27488 6372 27494 6384
rect 27893 6375 27951 6381
rect 27893 6372 27905 6375
rect 27488 6344 27905 6372
rect 27488 6332 27494 6344
rect 27893 6341 27905 6344
rect 27939 6341 27951 6375
rect 27893 6335 27951 6341
rect 30668 6344 31156 6372
rect 30668 6316 30696 6344
rect 26605 6307 26663 6313
rect 26605 6273 26617 6307
rect 26651 6273 26663 6307
rect 26605 6267 26663 6273
rect 26786 6264 26792 6316
rect 26844 6264 26850 6316
rect 27801 6307 27859 6313
rect 27801 6304 27813 6307
rect 27356 6276 27813 6304
rect 24581 6239 24639 6245
rect 24581 6236 24593 6239
rect 23256 6208 24593 6236
rect 23256 6196 23262 6208
rect 24581 6205 24593 6208
rect 24627 6236 24639 6239
rect 24762 6236 24768 6248
rect 24627 6208 24768 6236
rect 24627 6205 24639 6208
rect 24581 6199 24639 6205
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 12308 6140 12388 6168
rect 12308 6128 12314 6140
rect 12434 6128 12440 6180
rect 12492 6168 12498 6180
rect 12621 6171 12679 6177
rect 12621 6168 12633 6171
rect 12492 6140 12633 6168
rect 12492 6128 12498 6140
rect 12621 6137 12633 6140
rect 12667 6137 12679 6171
rect 12621 6131 12679 6137
rect 22646 6128 22652 6180
rect 22704 6168 22710 6180
rect 23937 6171 23995 6177
rect 23937 6168 23949 6171
rect 22704 6140 23949 6168
rect 22704 6128 22710 6140
rect 23937 6137 23949 6140
rect 23983 6137 23995 6171
rect 23937 6131 23995 6137
rect 26786 6128 26792 6180
rect 26844 6168 26850 6180
rect 27356 6177 27384 6276
rect 27801 6273 27813 6276
rect 27847 6273 27859 6307
rect 27801 6267 27859 6273
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 28445 6307 28503 6313
rect 28445 6273 28457 6307
rect 28491 6304 28503 6307
rect 28905 6307 28963 6313
rect 28905 6304 28917 6307
rect 28491 6276 28917 6304
rect 28491 6273 28503 6276
rect 28445 6267 28503 6273
rect 28905 6273 28917 6276
rect 28951 6304 28963 6307
rect 28994 6304 29000 6316
rect 28951 6276 29000 6304
rect 28951 6273 28963 6276
rect 28905 6267 28963 6273
rect 27706 6196 27712 6248
rect 27764 6236 27770 6248
rect 28092 6236 28120 6267
rect 28994 6264 29000 6276
rect 29052 6264 29058 6316
rect 29089 6307 29147 6313
rect 29089 6273 29101 6307
rect 29135 6273 29147 6307
rect 29089 6267 29147 6273
rect 27764 6208 28120 6236
rect 28353 6239 28411 6245
rect 27764 6196 27770 6208
rect 28353 6205 28365 6239
rect 28399 6236 28411 6239
rect 29104 6236 29132 6267
rect 29362 6264 29368 6316
rect 29420 6264 29426 6316
rect 29549 6307 29607 6313
rect 29549 6273 29561 6307
rect 29595 6304 29607 6307
rect 30469 6307 30527 6313
rect 30469 6304 30481 6307
rect 29595 6276 30481 6304
rect 29595 6273 29607 6276
rect 29549 6267 29607 6273
rect 30469 6273 30481 6276
rect 30515 6273 30527 6307
rect 30469 6267 30527 6273
rect 28399 6208 29132 6236
rect 30484 6236 30512 6267
rect 30650 6264 30656 6316
rect 30708 6264 30714 6316
rect 31128 6313 31156 6344
rect 31294 6332 31300 6384
rect 31352 6332 31358 6384
rect 31404 6313 31432 6412
rect 33318 6400 33324 6452
rect 33376 6400 33382 6452
rect 36081 6443 36139 6449
rect 36081 6409 36093 6443
rect 36127 6440 36139 6443
rect 36446 6440 36452 6452
rect 36127 6412 36452 6440
rect 36127 6409 36139 6412
rect 36081 6403 36139 6409
rect 36446 6400 36452 6412
rect 36504 6400 36510 6452
rect 31846 6332 31852 6384
rect 31904 6372 31910 6384
rect 31941 6375 31999 6381
rect 31941 6372 31953 6375
rect 31904 6344 31953 6372
rect 31904 6332 31910 6344
rect 31941 6341 31953 6344
rect 31987 6372 31999 6375
rect 32493 6375 32551 6381
rect 32493 6372 32505 6375
rect 31987 6344 32505 6372
rect 31987 6341 31999 6344
rect 31941 6335 31999 6341
rect 32493 6341 32505 6344
rect 32539 6341 32551 6375
rect 35434 6372 35440 6384
rect 32493 6335 32551 6341
rect 35176 6344 35440 6372
rect 30929 6307 30987 6313
rect 30929 6273 30941 6307
rect 30975 6273 30987 6307
rect 30929 6267 30987 6273
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6273 31171 6307
rect 31113 6267 31171 6273
rect 31205 6307 31263 6313
rect 31205 6273 31217 6307
rect 31251 6273 31263 6307
rect 31205 6267 31263 6273
rect 31389 6307 31447 6313
rect 31389 6273 31401 6307
rect 31435 6273 31447 6307
rect 31389 6267 31447 6273
rect 30944 6236 30972 6267
rect 30484 6208 30972 6236
rect 31021 6239 31079 6245
rect 28399 6205 28411 6208
rect 28353 6199 28411 6205
rect 31021 6205 31033 6239
rect 31067 6236 31079 6239
rect 31220 6236 31248 6267
rect 31067 6208 31248 6236
rect 31404 6236 31432 6267
rect 31570 6264 31576 6316
rect 31628 6264 31634 6316
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6304 31815 6307
rect 32125 6307 32183 6313
rect 32125 6304 32137 6307
rect 31803 6276 32137 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 32125 6273 32137 6276
rect 32171 6273 32183 6307
rect 32125 6267 32183 6273
rect 32309 6307 32367 6313
rect 32309 6273 32321 6307
rect 32355 6273 32367 6307
rect 32309 6267 32367 6273
rect 31772 6236 31800 6267
rect 31404 6208 31800 6236
rect 31067 6205 31079 6208
rect 31021 6199 31079 6205
rect 27341 6171 27399 6177
rect 27341 6168 27353 6171
rect 26844 6140 27353 6168
rect 26844 6128 26850 6140
rect 27341 6137 27353 6140
rect 27387 6137 27399 6171
rect 27341 6131 27399 6137
rect 28077 6171 28135 6177
rect 28077 6137 28089 6171
rect 28123 6168 28135 6171
rect 28368 6168 28396 6199
rect 28123 6140 28396 6168
rect 28123 6137 28135 6140
rect 28077 6131 28135 6137
rect 31570 6128 31576 6180
rect 31628 6168 31634 6180
rect 32324 6168 32352 6267
rect 32398 6264 32404 6316
rect 32456 6264 32462 6316
rect 32677 6307 32735 6313
rect 32677 6273 32689 6307
rect 32723 6304 32735 6307
rect 32766 6304 32772 6316
rect 32723 6276 32772 6304
rect 32723 6273 32735 6276
rect 32677 6267 32735 6273
rect 32766 6264 32772 6276
rect 32824 6264 32830 6316
rect 33134 6264 33140 6316
rect 33192 6264 33198 6316
rect 34606 6264 34612 6316
rect 34664 6264 34670 6316
rect 34790 6313 34796 6316
rect 34757 6307 34796 6313
rect 34757 6273 34769 6307
rect 34757 6267 34796 6273
rect 34790 6264 34796 6267
rect 34848 6264 34854 6316
rect 34885 6307 34943 6313
rect 34885 6273 34897 6307
rect 34931 6273 34943 6307
rect 34885 6267 34943 6273
rect 34977 6307 35035 6313
rect 34977 6273 34989 6307
rect 35023 6273 35035 6307
rect 34977 6267 35035 6273
rect 35074 6307 35132 6313
rect 35074 6273 35086 6307
rect 35120 6304 35132 6307
rect 35176 6304 35204 6344
rect 35434 6332 35440 6344
rect 35492 6332 35498 6384
rect 35529 6307 35587 6313
rect 35529 6304 35541 6307
rect 35120 6276 35204 6304
rect 35268 6276 35541 6304
rect 35120 6273 35132 6276
rect 35074 6267 35132 6273
rect 32861 6239 32919 6245
rect 32861 6205 32873 6239
rect 32907 6236 32919 6239
rect 32953 6239 33011 6245
rect 32953 6236 32965 6239
rect 32907 6208 32965 6236
rect 32907 6205 32919 6208
rect 32861 6199 32919 6205
rect 32953 6205 32965 6208
rect 32999 6236 33011 6239
rect 33318 6236 33324 6248
rect 32999 6208 33324 6236
rect 32999 6205 33011 6208
rect 32953 6199 33011 6205
rect 33318 6196 33324 6208
rect 33376 6196 33382 6248
rect 34422 6196 34428 6248
rect 34480 6236 34486 6248
rect 34900 6236 34928 6267
rect 34480 6208 34928 6236
rect 34480 6196 34486 6208
rect 31628 6140 32352 6168
rect 31628 6128 31634 6140
rect 34790 6128 34796 6180
rect 34848 6168 34854 6180
rect 34992 6168 35020 6267
rect 35268 6177 35296 6276
rect 35529 6273 35541 6276
rect 35575 6273 35587 6307
rect 35529 6267 35587 6273
rect 35618 6264 35624 6316
rect 35676 6304 35682 6316
rect 35713 6307 35771 6313
rect 35713 6304 35725 6307
rect 35676 6276 35725 6304
rect 35676 6264 35682 6276
rect 35713 6273 35725 6276
rect 35759 6273 35771 6307
rect 35713 6267 35771 6273
rect 35805 6307 35863 6313
rect 35805 6273 35817 6307
rect 35851 6273 35863 6307
rect 35805 6267 35863 6273
rect 35897 6307 35955 6313
rect 35897 6273 35909 6307
rect 35943 6304 35955 6307
rect 35986 6304 35992 6316
rect 35943 6276 35992 6304
rect 35943 6273 35955 6276
rect 35897 6267 35955 6273
rect 35342 6196 35348 6248
rect 35400 6236 35406 6248
rect 35820 6236 35848 6267
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 35400 6208 35848 6236
rect 35400 6196 35406 6208
rect 34848 6140 35020 6168
rect 35253 6171 35311 6177
rect 34848 6128 34854 6140
rect 35253 6137 35265 6171
rect 35299 6137 35311 6171
rect 35253 6131 35311 6137
rect 5215 6072 8156 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8754 6100 8760 6112
rect 8260 6072 8760 6100
rect 8260 6060 8266 6072
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 9953 6103 10011 6109
rect 9953 6069 9965 6103
rect 9999 6100 10011 6103
rect 10686 6100 10692 6112
rect 9999 6072 10692 6100
rect 9999 6069 10011 6072
rect 9953 6063 10011 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 11020 6072 11161 6100
rect 11020 6060 11026 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11296 6072 11529 6100
rect 11296 6060 11302 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 11974 6060 11980 6112
rect 12032 6060 12038 6112
rect 22738 6060 22744 6112
rect 22796 6100 22802 6112
rect 23017 6103 23075 6109
rect 23017 6100 23029 6103
rect 22796 6072 23029 6100
rect 22796 6060 22802 6072
rect 23017 6069 23029 6072
rect 23063 6069 23075 6103
rect 23017 6063 23075 6069
rect 24765 6103 24823 6109
rect 24765 6069 24777 6103
rect 24811 6100 24823 6103
rect 25038 6100 25044 6112
rect 24811 6072 25044 6100
rect 24811 6069 24823 6072
rect 24765 6063 24823 6069
rect 25038 6060 25044 6072
rect 25096 6060 25102 6112
rect 26418 6060 26424 6112
rect 26476 6100 26482 6112
rect 26605 6103 26663 6109
rect 26605 6100 26617 6103
rect 26476 6072 26617 6100
rect 26476 6060 26482 6072
rect 26605 6069 26617 6072
rect 26651 6069 26663 6103
rect 26605 6063 26663 6069
rect 32030 6060 32036 6112
rect 32088 6100 32094 6112
rect 32217 6103 32275 6109
rect 32217 6100 32229 6103
rect 32088 6072 32229 6100
rect 32088 6060 32094 6072
rect 32217 6069 32229 6072
rect 32263 6069 32275 6103
rect 32217 6063 32275 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5534 5896 5540 5908
rect 5215 5868 5540 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 9122 5896 9128 5908
rect 8435 5868 9128 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 2590 5760 2596 5772
rect 1903 5732 2596 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 3605 5763 3663 5769
rect 3605 5729 3617 5763
rect 3651 5760 3663 5763
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 3651 5732 4629 5760
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 4617 5729 4629 5732
rect 4663 5760 4675 5763
rect 4706 5760 4712 5772
rect 4663 5732 4712 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 4706 5720 4712 5732
rect 4764 5760 4770 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4764 5732 4813 5760
rect 4764 5720 4770 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 7742 5720 7748 5772
rect 7800 5720 7806 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 8404 5760 8432 5859
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9585 5899 9643 5905
rect 9585 5865 9597 5899
rect 9631 5865 9643 5899
rect 9585 5859 9643 5865
rect 9493 5763 9551 5769
rect 7883 5732 8432 5760
rect 8956 5732 9444 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 842 5652 848 5704
rect 900 5692 906 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 900 5664 1409 5692
rect 900 5652 906 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 3878 5692 3884 5704
rect 3835 5664 3884 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 2133 5627 2191 5633
rect 2133 5593 2145 5627
rect 2179 5593 2191 5627
rect 2133 5587 2191 5593
rect 2148 5556 2176 5587
rect 3142 5584 3148 5636
rect 3200 5584 3206 5636
rect 3804 5624 3832 5655
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 4019 5664 4077 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5000 5624 5028 5655
rect 5626 5652 5632 5704
rect 5684 5652 5690 5704
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 5994 5692 6000 5704
rect 5859 5664 6000 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 6641 5695 6699 5701
rect 6641 5692 6653 5695
rect 6604 5664 6653 5692
rect 6604 5652 6610 5664
rect 6641 5661 6653 5664
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5692 8079 5695
rect 8110 5692 8116 5704
rect 8067 5664 8116 5692
rect 8067 5661 8079 5664
rect 8021 5655 8079 5661
rect 8110 5652 8116 5664
rect 8168 5692 8174 5704
rect 8956 5692 8984 5732
rect 8168 5664 8984 5692
rect 8168 5652 8174 5664
rect 9030 5652 9036 5704
rect 9088 5652 9094 5704
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 3804 5596 5028 5624
rect 7576 5624 7604 5652
rect 8357 5627 8415 5633
rect 8357 5624 8369 5627
rect 7576 5596 8369 5624
rect 8357 5593 8369 5596
rect 8403 5593 8415 5627
rect 8357 5587 8415 5593
rect 8570 5584 8576 5636
rect 8628 5584 8634 5636
rect 9214 5584 9220 5636
rect 9272 5584 9278 5636
rect 9306 5584 9312 5636
rect 9364 5584 9370 5636
rect 2958 5556 2964 5568
rect 2148 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3752 5528 3893 5556
rect 3752 5516 3758 5528
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 3881 5519 3939 5525
rect 5718 5516 5724 5568
rect 5776 5516 5782 5568
rect 6086 5516 6092 5568
rect 6144 5516 6150 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 7156 5528 7573 5556
rect 7156 5516 7162 5528
rect 7561 5525 7573 5528
rect 7607 5525 7619 5559
rect 8588 5556 8616 5584
rect 9324 5556 9352 5584
rect 8588 5528 9352 5556
rect 9416 5556 9444 5732
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 9600 5760 9628 5859
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 10505 5899 10563 5905
rect 10505 5865 10517 5899
rect 10551 5896 10563 5899
rect 10551 5868 11284 5896
rect 10551 5865 10563 5868
rect 10505 5859 10563 5865
rect 10045 5831 10103 5837
rect 10045 5797 10057 5831
rect 10091 5797 10103 5831
rect 10045 5791 10103 5797
rect 10781 5831 10839 5837
rect 10781 5797 10793 5831
rect 10827 5828 10839 5831
rect 11146 5828 11152 5840
rect 10827 5800 11152 5828
rect 10827 5797 10839 5800
rect 10781 5791 10839 5797
rect 9539 5732 9628 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 9674 5720 9680 5772
rect 9732 5720 9738 5772
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 9582 5584 9588 5636
rect 9640 5584 9646 5636
rect 10060 5624 10088 5791
rect 11146 5788 11152 5800
rect 11204 5788 11210 5840
rect 11256 5828 11284 5868
rect 11422 5856 11428 5908
rect 11480 5856 11486 5908
rect 22830 5856 22836 5908
rect 22888 5896 22894 5908
rect 23477 5899 23535 5905
rect 23477 5896 23489 5899
rect 22888 5868 23489 5896
rect 22888 5856 22894 5868
rect 23477 5865 23489 5868
rect 23523 5865 23535 5899
rect 23477 5859 23535 5865
rect 26786 5856 26792 5908
rect 26844 5856 26850 5908
rect 27617 5899 27675 5905
rect 27617 5865 27629 5899
rect 27663 5896 27675 5899
rect 27706 5896 27712 5908
rect 27663 5868 27712 5896
rect 27663 5865 27675 5868
rect 27617 5859 27675 5865
rect 27706 5856 27712 5868
rect 27764 5856 27770 5908
rect 30101 5899 30159 5905
rect 30101 5865 30113 5899
rect 30147 5896 30159 5899
rect 30650 5896 30656 5908
rect 30147 5868 30656 5896
rect 30147 5865 30159 5868
rect 30101 5859 30159 5865
rect 30650 5856 30656 5868
rect 30708 5856 30714 5908
rect 31941 5899 31999 5905
rect 31941 5865 31953 5899
rect 31987 5896 31999 5899
rect 32306 5896 32312 5908
rect 31987 5868 32312 5896
rect 31987 5865 31999 5868
rect 31941 5859 31999 5865
rect 32306 5856 32312 5868
rect 32364 5856 32370 5908
rect 32769 5899 32827 5905
rect 32769 5865 32781 5899
rect 32815 5896 32827 5899
rect 33134 5896 33140 5908
rect 32815 5868 33140 5896
rect 32815 5865 32827 5868
rect 32769 5859 32827 5865
rect 33134 5856 33140 5868
rect 33192 5856 33198 5908
rect 33781 5899 33839 5905
rect 33781 5865 33793 5899
rect 33827 5896 33839 5899
rect 33870 5896 33876 5908
rect 33827 5868 33876 5896
rect 33827 5865 33839 5868
rect 33781 5859 33839 5865
rect 33870 5856 33876 5868
rect 33928 5856 33934 5908
rect 34422 5856 34428 5908
rect 34480 5856 34486 5908
rect 34606 5856 34612 5908
rect 34664 5896 34670 5908
rect 34701 5899 34759 5905
rect 34701 5896 34713 5899
rect 34664 5868 34713 5896
rect 34664 5856 34670 5868
rect 34701 5865 34713 5868
rect 34747 5865 34759 5899
rect 34701 5859 34759 5865
rect 35161 5899 35219 5905
rect 35161 5865 35173 5899
rect 35207 5896 35219 5899
rect 35434 5896 35440 5908
rect 35207 5868 35440 5896
rect 35207 5865 35219 5868
rect 35161 5859 35219 5865
rect 35434 5856 35440 5868
rect 35492 5856 35498 5908
rect 35618 5856 35624 5908
rect 35676 5856 35682 5908
rect 11701 5831 11759 5837
rect 11701 5828 11713 5831
rect 11256 5800 11713 5828
rect 11701 5797 11713 5800
rect 11747 5797 11759 5831
rect 11701 5791 11759 5797
rect 22370 5788 22376 5840
rect 22428 5828 22434 5840
rect 22925 5831 22983 5837
rect 22925 5828 22937 5831
rect 22428 5800 22937 5828
rect 22428 5788 22434 5800
rect 22925 5797 22937 5800
rect 22971 5797 22983 5831
rect 22925 5791 22983 5797
rect 23124 5800 25084 5828
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10962 5760 10968 5772
rect 10459 5732 10968 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11471 5732 12081 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 12345 5763 12403 5769
rect 12345 5729 12357 5763
rect 12391 5760 12403 5763
rect 12894 5760 12900 5772
rect 12391 5732 12900 5760
rect 12391 5729 12403 5732
rect 12345 5723 12403 5729
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 13173 5763 13231 5769
rect 13173 5729 13185 5763
rect 13219 5760 13231 5763
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 13219 5732 15577 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 21726 5720 21732 5772
rect 21784 5720 21790 5772
rect 22554 5720 22560 5772
rect 22612 5720 22618 5772
rect 22741 5763 22799 5769
rect 22741 5729 22753 5763
rect 22787 5760 22799 5763
rect 22830 5760 22836 5772
rect 22787 5732 22836 5760
rect 22787 5729 22799 5732
rect 22741 5723 22799 5729
rect 22830 5720 22836 5732
rect 22888 5720 22894 5772
rect 10502 5652 10508 5704
rect 10560 5652 10566 5704
rect 10686 5652 10692 5704
rect 10744 5652 10750 5704
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5692 10931 5695
rect 11146 5692 11152 5704
rect 10919 5664 11152 5692
rect 10919 5661 10931 5664
rect 10873 5655 10931 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5692 11575 5695
rect 11882 5692 11888 5704
rect 11563 5664 11888 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 10597 5627 10655 5633
rect 10597 5624 10609 5627
rect 10060 5596 10609 5624
rect 10597 5593 10609 5596
rect 10643 5593 10655 5627
rect 10704 5624 10732 5652
rect 11057 5627 11115 5633
rect 11057 5624 11069 5627
rect 10704 5596 11069 5624
rect 10597 5587 10655 5593
rect 11057 5593 11069 5596
rect 11103 5593 11115 5627
rect 11057 5587 11115 5593
rect 11422 5584 11428 5636
rect 11480 5624 11486 5636
rect 11992 5624 12020 5655
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 12250 5652 12256 5704
rect 12308 5652 12314 5704
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5692 12495 5695
rect 12526 5692 12532 5704
rect 12483 5664 12532 5692
rect 12483 5661 12495 5664
rect 12437 5655 12495 5661
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 12851 5664 13277 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 13354 5652 13360 5704
rect 13412 5692 13418 5704
rect 13817 5695 13875 5701
rect 13817 5692 13829 5695
rect 13412 5664 13829 5692
rect 13412 5652 13418 5664
rect 13817 5661 13829 5664
rect 13863 5661 13875 5695
rect 13817 5655 13875 5661
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 16666 5692 16672 5704
rect 15896 5664 16672 5692
rect 15896 5652 15902 5664
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 22646 5692 22652 5704
rect 22511 5664 22652 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 22925 5695 22983 5701
rect 22925 5661 22937 5695
rect 22971 5692 22983 5695
rect 23014 5692 23020 5704
rect 22971 5664 23020 5692
rect 22971 5661 22983 5664
rect 22925 5655 22983 5661
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 11480 5596 12020 5624
rect 11480 5584 11486 5596
rect 12710 5584 12716 5636
rect 12768 5624 12774 5636
rect 21545 5627 21603 5633
rect 12768 5596 14398 5624
rect 12768 5584 12774 5596
rect 21545 5593 21557 5627
rect 21591 5624 21603 5627
rect 22002 5624 22008 5636
rect 21591 5596 22008 5624
rect 21591 5593 21603 5596
rect 21545 5587 21603 5593
rect 22002 5584 22008 5596
rect 22060 5584 22066 5636
rect 23124 5633 23152 5800
rect 23290 5720 23296 5772
rect 23348 5720 23354 5772
rect 24302 5760 24308 5772
rect 23584 5732 24308 5760
rect 23198 5652 23204 5704
rect 23256 5652 23262 5704
rect 23474 5652 23480 5704
rect 23532 5692 23538 5704
rect 23584 5701 23612 5732
rect 24302 5720 24308 5732
rect 24360 5760 24366 5772
rect 25056 5760 25084 5800
rect 25130 5788 25136 5840
rect 25188 5788 25194 5840
rect 25314 5760 25320 5772
rect 24360 5732 24905 5760
rect 25056 5732 25320 5760
rect 24360 5720 24366 5732
rect 23569 5695 23627 5701
rect 23569 5692 23581 5695
rect 23532 5664 23581 5692
rect 23532 5652 23538 5664
rect 23569 5661 23581 5664
rect 23615 5661 23627 5695
rect 23569 5655 23627 5661
rect 23842 5652 23848 5704
rect 23900 5692 23906 5704
rect 24877 5701 24905 5732
rect 25314 5720 25320 5732
rect 25372 5760 25378 5772
rect 26329 5763 26387 5769
rect 26329 5760 26341 5763
rect 25372 5732 26341 5760
rect 25372 5720 25378 5732
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 23900 5664 24409 5692
rect 23900 5652 23906 5664
rect 24397 5661 24409 5664
rect 24443 5661 24455 5695
rect 24397 5655 24455 5661
rect 24545 5695 24603 5701
rect 24545 5661 24557 5695
rect 24591 5692 24603 5695
rect 24877 5695 24959 5701
rect 24591 5661 24624 5692
rect 24545 5655 24624 5661
rect 24877 5661 24913 5695
rect 24947 5661 24959 5695
rect 24877 5658 24959 5661
rect 24901 5655 24959 5658
rect 23109 5627 23167 5633
rect 23109 5593 23121 5627
rect 23155 5593 23167 5627
rect 23109 5587 23167 5593
rect 10689 5559 10747 5565
rect 10689 5556 10701 5559
rect 9416 5528 10701 5556
rect 7561 5519 7619 5525
rect 10689 5525 10701 5528
rect 10735 5556 10747 5559
rect 11882 5556 11888 5568
rect 10735 5528 11888 5556
rect 10735 5525 10747 5528
rect 10689 5519 10747 5525
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 13354 5516 13360 5568
rect 13412 5556 13418 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13412 5528 14105 5556
rect 13412 5516 13418 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 21174 5516 21180 5568
rect 21232 5516 21238 5568
rect 21637 5559 21695 5565
rect 21637 5525 21649 5559
rect 21683 5556 21695 5559
rect 22097 5559 22155 5565
rect 22097 5556 22109 5559
rect 21683 5528 22109 5556
rect 21683 5525 21695 5528
rect 21637 5519 21695 5525
rect 22097 5525 22109 5528
rect 22143 5525 22155 5559
rect 22097 5519 22155 5525
rect 23290 5516 23296 5568
rect 23348 5516 23354 5568
rect 24596 5556 24624 5655
rect 25038 5652 25044 5704
rect 25096 5692 25102 5704
rect 25424 5701 25452 5732
rect 26329 5729 26341 5732
rect 26375 5729 26387 5763
rect 26329 5723 26387 5729
rect 26528 5732 27384 5760
rect 25133 5695 25191 5701
rect 25133 5692 25145 5695
rect 25096 5664 25145 5692
rect 25096 5652 25102 5664
rect 25133 5661 25145 5664
rect 25179 5661 25191 5695
rect 25133 5655 25191 5661
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5661 25467 5695
rect 25409 5655 25467 5661
rect 25869 5695 25927 5701
rect 25869 5661 25881 5695
rect 25915 5661 25927 5695
rect 25869 5655 25927 5661
rect 25961 5695 26019 5701
rect 25961 5661 25973 5695
rect 26007 5692 26019 5695
rect 26050 5692 26056 5704
rect 26007 5664 26056 5692
rect 26007 5661 26019 5664
rect 25961 5655 26019 5661
rect 24670 5584 24676 5636
rect 24728 5584 24734 5636
rect 24765 5627 24823 5633
rect 24765 5593 24777 5627
rect 24811 5624 24823 5627
rect 25222 5624 25228 5636
rect 24811 5596 25228 5624
rect 24811 5593 24823 5596
rect 24765 5587 24823 5593
rect 25222 5584 25228 5596
rect 25280 5624 25286 5636
rect 25317 5627 25375 5633
rect 25317 5624 25329 5627
rect 25280 5596 25329 5624
rect 25280 5584 25286 5596
rect 25317 5593 25329 5596
rect 25363 5624 25375 5627
rect 25590 5624 25596 5636
rect 25363 5596 25596 5624
rect 25363 5593 25375 5596
rect 25317 5587 25375 5593
rect 25590 5584 25596 5596
rect 25648 5584 25654 5636
rect 25884 5624 25912 5655
rect 26050 5652 26056 5664
rect 26108 5652 26114 5704
rect 26145 5695 26203 5701
rect 26145 5661 26157 5695
rect 26191 5692 26203 5695
rect 26237 5695 26295 5701
rect 26237 5692 26249 5695
rect 26191 5664 26249 5692
rect 26191 5661 26203 5664
rect 26145 5655 26203 5661
rect 26237 5661 26249 5664
rect 26283 5661 26295 5695
rect 26237 5655 26295 5661
rect 26418 5652 26424 5704
rect 26476 5652 26482 5704
rect 26528 5624 26556 5732
rect 27356 5704 27384 5732
rect 34348 5732 34744 5760
rect 27249 5695 27307 5701
rect 27249 5692 27261 5695
rect 26988 5664 27261 5692
rect 26988 5633 27016 5664
rect 27249 5661 27261 5664
rect 27295 5661 27307 5695
rect 27249 5655 27307 5661
rect 27338 5652 27344 5704
rect 27396 5692 27402 5704
rect 27433 5695 27491 5701
rect 27433 5692 27445 5695
rect 27396 5664 27445 5692
rect 27396 5652 27402 5664
rect 27433 5661 27445 5664
rect 27479 5661 27491 5695
rect 27433 5655 27491 5661
rect 31846 5652 31852 5704
rect 31904 5652 31910 5704
rect 32030 5652 32036 5704
rect 32088 5652 32094 5704
rect 32398 5652 32404 5704
rect 32456 5692 32462 5704
rect 32493 5695 32551 5701
rect 32493 5692 32505 5695
rect 32456 5664 32505 5692
rect 32456 5652 32462 5664
rect 32493 5661 32505 5664
rect 32539 5661 32551 5695
rect 32493 5655 32551 5661
rect 32766 5652 32772 5704
rect 32824 5652 32830 5704
rect 33778 5652 33784 5704
rect 33836 5652 33842 5704
rect 33870 5652 33876 5704
rect 33928 5692 33934 5704
rect 34348 5701 34376 5732
rect 34716 5704 34744 5732
rect 34790 5720 34796 5772
rect 34848 5760 34854 5772
rect 34848 5732 35112 5760
rect 34848 5720 34854 5732
rect 35084 5704 35112 5732
rect 33965 5695 34023 5701
rect 33965 5692 33977 5695
rect 33928 5664 33977 5692
rect 33928 5652 33934 5664
rect 33965 5661 33977 5664
rect 34011 5661 34023 5695
rect 33965 5655 34023 5661
rect 34333 5695 34391 5701
rect 34333 5661 34345 5695
rect 34379 5661 34391 5695
rect 34333 5655 34391 5661
rect 34514 5652 34520 5704
rect 34572 5652 34578 5704
rect 34698 5652 34704 5704
rect 34756 5652 34762 5704
rect 34885 5695 34943 5701
rect 34885 5661 34897 5695
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 25884 5596 26556 5624
rect 26973 5627 27031 5633
rect 26973 5593 26985 5627
rect 27019 5593 27031 5627
rect 26973 5587 27031 5593
rect 24854 5556 24860 5568
rect 24596 5528 24860 5556
rect 24854 5516 24860 5528
rect 24912 5516 24918 5568
rect 25038 5516 25044 5568
rect 25096 5516 25102 5568
rect 25958 5516 25964 5568
rect 26016 5556 26022 5568
rect 26988 5556 27016 5587
rect 27154 5584 27160 5636
rect 27212 5584 27218 5636
rect 29730 5584 29736 5636
rect 29788 5584 29794 5636
rect 29822 5584 29828 5636
rect 29880 5624 29886 5636
rect 29917 5627 29975 5633
rect 29917 5624 29929 5627
rect 29880 5596 29929 5624
rect 29880 5584 29886 5596
rect 29917 5593 29929 5596
rect 29963 5593 29975 5627
rect 31864 5624 31892 5652
rect 32677 5627 32735 5633
rect 32677 5624 32689 5627
rect 31864 5596 32689 5624
rect 29917 5587 29975 5593
rect 32677 5593 32689 5596
rect 32723 5593 32735 5627
rect 34532 5624 34560 5652
rect 34900 5624 34928 5655
rect 35066 5652 35072 5704
rect 35124 5652 35130 5704
rect 35342 5652 35348 5704
rect 35400 5652 35406 5704
rect 35437 5695 35495 5701
rect 35437 5661 35449 5695
rect 35483 5692 35495 5695
rect 35802 5692 35808 5704
rect 35483 5664 35808 5692
rect 35483 5661 35495 5664
rect 35437 5655 35495 5661
rect 35802 5652 35808 5664
rect 35860 5652 35866 5704
rect 34532 5596 34928 5624
rect 32677 5587 32735 5593
rect 26016 5528 27016 5556
rect 26016 5516 26022 5528
rect 1104 5466 38824 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 38824 5466
rect 1104 5392 38824 5414
rect 2958 5312 2964 5364
rect 3016 5312 3022 5364
rect 3786 5312 3792 5364
rect 3844 5352 3850 5364
rect 3844 5324 4568 5352
rect 3844 5312 3850 5324
rect 3881 5287 3939 5293
rect 3881 5253 3893 5287
rect 3927 5284 3939 5287
rect 4154 5284 4160 5296
rect 3927 5256 4160 5284
rect 3927 5253 3939 5256
rect 3881 5247 3939 5253
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 4540 5284 4568 5324
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5684 5324 6377 5352
rect 5684 5312 5690 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6533 5355 6591 5361
rect 6533 5321 6545 5355
rect 6579 5352 6591 5355
rect 6914 5352 6920 5364
rect 6579 5324 6920 5352
rect 6579 5321 6591 5324
rect 6533 5315 6591 5321
rect 6914 5312 6920 5324
rect 6972 5352 6978 5364
rect 7374 5352 7380 5364
rect 6972 5324 7380 5352
rect 6972 5312 6978 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 9585 5355 9643 5361
rect 9585 5321 9597 5355
rect 9631 5352 9643 5355
rect 10502 5352 10508 5364
rect 9631 5324 10508 5352
rect 9631 5321 9643 5324
rect 9585 5315 9643 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 13354 5352 13360 5364
rect 11992 5324 13360 5352
rect 11992 5296 12020 5324
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 22002 5312 22008 5364
rect 22060 5312 22066 5364
rect 22646 5352 22652 5364
rect 22388 5324 22652 5352
rect 4798 5284 4804 5296
rect 4540 5256 4804 5284
rect 4798 5244 4804 5256
rect 4856 5284 4862 5296
rect 6733 5287 6791 5293
rect 4856 5256 5198 5284
rect 4856 5244 4862 5256
rect 6733 5253 6745 5287
rect 6779 5284 6791 5287
rect 6779 5256 7604 5284
rect 6779 5253 6791 5256
rect 6733 5247 6791 5253
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3694 5216 3700 5228
rect 3099 5188 3700 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 4172 5216 4200 5244
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 4172 5188 4445 5216
rect 4433 5185 4445 5188
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6748 5216 6776 5247
rect 6236 5188 6776 5216
rect 6236 5176 6242 5188
rect 7098 5176 7104 5228
rect 7156 5176 7162 5228
rect 7374 5176 7380 5228
rect 7432 5176 7438 5228
rect 7576 5225 7604 5256
rect 11974 5244 11980 5296
rect 12032 5244 12038 5296
rect 12193 5287 12251 5293
rect 12193 5253 12205 5287
rect 12239 5284 12251 5287
rect 12894 5284 12900 5296
rect 12239 5256 12900 5284
rect 12239 5253 12251 5256
rect 12193 5247 12251 5253
rect 12894 5244 12900 5256
rect 12952 5284 12958 5296
rect 21358 5284 21364 5296
rect 12952 5256 13492 5284
rect 21206 5256 21364 5284
rect 12952 5244 12958 5256
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7926 5216 7932 5228
rect 7607 5188 7932 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7926 5176 7932 5188
rect 7984 5216 7990 5228
rect 8294 5216 8300 5228
rect 7984 5188 8300 5216
rect 7984 5176 7990 5188
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 9401 5219 9459 5225
rect 9171 5188 9352 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 842 5108 848 5160
rect 900 5148 906 5160
rect 1397 5151 1455 5157
rect 1397 5148 1409 5151
rect 900 5120 1409 5148
rect 900 5108 906 5120
rect 1397 5117 1409 5120
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 5718 5148 5724 5160
rect 4755 5120 5724 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 7392 5148 7420 5176
rect 8202 5148 8208 5160
rect 7392 5120 8208 5148
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8386 5108 8392 5160
rect 8444 5148 8450 5160
rect 9217 5151 9275 5157
rect 9217 5148 9229 5151
rect 8444 5120 9229 5148
rect 8444 5108 8450 5120
rect 9217 5117 9229 5120
rect 9263 5117 9275 5151
rect 9324 5148 9352 5188
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9490 5216 9496 5228
rect 9447 5188 9496 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 9490 5176 9496 5188
rect 9548 5216 9554 5228
rect 9858 5216 9864 5228
rect 9548 5188 9864 5216
rect 9548 5176 9554 5188
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11238 5216 11244 5228
rect 11195 5188 11244 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 12802 5216 12808 5228
rect 11992 5188 12808 5216
rect 9674 5148 9680 5160
rect 9324 5120 9680 5148
rect 9217 5111 9275 5117
rect 6181 5083 6239 5089
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 9232 5080 9260 5111
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 11992 5148 12020 5188
rect 12802 5176 12808 5188
rect 12860 5216 12866 5228
rect 13464 5225 13492 5256
rect 21358 5244 21364 5256
rect 21416 5284 21422 5296
rect 22388 5284 22416 5324
rect 22646 5312 22652 5324
rect 22704 5312 22710 5364
rect 22922 5312 22928 5364
rect 22980 5312 22986 5364
rect 24302 5312 24308 5364
rect 24360 5352 24366 5364
rect 29549 5355 29607 5361
rect 24360 5324 25452 5352
rect 24360 5312 24366 5324
rect 23290 5284 23296 5296
rect 21416 5256 22416 5284
rect 22480 5256 23296 5284
rect 21416 5244 21422 5256
rect 13081 5219 13139 5225
rect 12860 5188 13032 5216
rect 12860 5176 12866 5188
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 11348 5120 12020 5148
rect 12176 5120 12449 5148
rect 9582 5080 9588 5092
rect 6227 5052 6592 5080
rect 9232 5052 9588 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 6564 5024 6592 5052
rect 9582 5040 9588 5052
rect 9640 5040 9646 5092
rect 11348 5089 11376 5120
rect 11333 5083 11391 5089
rect 11333 5049 11345 5083
rect 11379 5049 11391 5083
rect 11333 5043 11391 5049
rect 12176 5024 12204 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 13004 5148 13032 5188
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 13127 5188 13185 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 18564 5188 19809 5216
rect 18564 5176 18570 5188
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 21591 5219 21649 5225
rect 21591 5185 21603 5219
rect 21637 5216 21649 5219
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21637 5188 21833 5216
rect 21637 5185 21649 5188
rect 21591 5179 21649 5185
rect 21821 5185 21833 5188
rect 21867 5216 21879 5219
rect 21867 5188 22094 5216
rect 21867 5185 21879 5188
rect 21821 5179 21879 5185
rect 13722 5148 13728 5160
rect 13004 5120 13728 5148
rect 12437 5111 12495 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 20165 5151 20223 5157
rect 20165 5117 20177 5151
rect 20211 5148 20223 5151
rect 21174 5148 21180 5160
rect 20211 5120 21180 5148
rect 20211 5117 20223 5120
rect 20165 5111 20223 5117
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 22066 5148 22094 5188
rect 22370 5176 22376 5228
rect 22428 5176 22434 5228
rect 22480 5225 22508 5256
rect 23290 5244 23296 5256
rect 23348 5244 23354 5296
rect 24854 5244 24860 5296
rect 24912 5244 24918 5296
rect 25130 5244 25136 5296
rect 25188 5284 25194 5296
rect 25424 5293 25452 5324
rect 29549 5321 29561 5355
rect 29595 5352 29607 5355
rect 29730 5352 29736 5364
rect 29595 5324 29736 5352
rect 29595 5321 29607 5324
rect 29549 5315 29607 5321
rect 29730 5312 29736 5324
rect 29788 5312 29794 5364
rect 29822 5312 29828 5364
rect 29880 5312 29886 5364
rect 31205 5355 31263 5361
rect 31205 5321 31217 5355
rect 31251 5352 31263 5355
rect 31570 5352 31576 5364
rect 31251 5324 31576 5352
rect 31251 5321 31263 5324
rect 31205 5315 31263 5321
rect 31570 5312 31576 5324
rect 31628 5312 31634 5364
rect 31941 5355 31999 5361
rect 31941 5321 31953 5355
rect 31987 5352 31999 5355
rect 32677 5355 32735 5361
rect 31987 5324 32628 5352
rect 31987 5321 31999 5324
rect 31941 5315 31999 5321
rect 25317 5287 25375 5293
rect 25317 5284 25329 5287
rect 25188 5256 25329 5284
rect 25188 5244 25194 5256
rect 25317 5253 25329 5256
rect 25363 5253 25375 5287
rect 25317 5247 25375 5253
rect 25409 5287 25467 5293
rect 25409 5253 25421 5287
rect 25455 5253 25467 5287
rect 25409 5247 25467 5253
rect 25590 5244 25596 5296
rect 25648 5244 25654 5296
rect 29840 5284 29868 5312
rect 32401 5287 32459 5293
rect 29380 5256 29776 5284
rect 29840 5256 30144 5284
rect 29380 5228 29408 5256
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 22738 5176 22744 5228
rect 22796 5176 22802 5228
rect 22830 5176 22836 5228
rect 22888 5216 22894 5228
rect 23017 5219 23075 5225
rect 23017 5216 23029 5219
rect 22888 5188 23029 5216
rect 22888 5176 22894 5188
rect 23017 5185 23029 5188
rect 23063 5216 23075 5219
rect 23934 5216 23940 5228
rect 23063 5188 23940 5216
rect 23063 5185 23075 5188
rect 23017 5179 23075 5185
rect 23934 5176 23940 5188
rect 23992 5176 23998 5228
rect 25041 5219 25099 5225
rect 25041 5185 25053 5219
rect 25087 5185 25099 5219
rect 25041 5179 25099 5185
rect 25056 5148 25084 5179
rect 25222 5176 25228 5228
rect 25280 5176 25286 5228
rect 29362 5176 29368 5228
rect 29420 5176 29426 5228
rect 29641 5219 29699 5225
rect 29641 5185 29653 5219
rect 29687 5185 29699 5219
rect 29748 5216 29776 5256
rect 30116 5225 30144 5256
rect 31496 5256 32168 5284
rect 29825 5219 29883 5225
rect 29825 5216 29837 5219
rect 29748 5188 29837 5216
rect 29641 5179 29699 5185
rect 29825 5185 29837 5188
rect 29871 5185 29883 5219
rect 29825 5179 29883 5185
rect 29917 5219 29975 5225
rect 29917 5185 29929 5219
rect 29963 5185 29975 5219
rect 29917 5179 29975 5185
rect 30101 5219 30159 5225
rect 30101 5185 30113 5219
rect 30147 5185 30159 5219
rect 30101 5179 30159 5185
rect 25406 5148 25412 5160
rect 22066 5120 24992 5148
rect 25056 5120 25412 5148
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 22649 5083 22707 5089
rect 22649 5080 22661 5083
rect 21784 5052 22661 5080
rect 21784 5040 21790 5052
rect 22649 5049 22661 5052
rect 22695 5080 22707 5083
rect 24486 5080 24492 5092
rect 22695 5052 24492 5080
rect 22695 5049 22707 5052
rect 22649 5043 22707 5049
rect 24486 5040 24492 5052
rect 24544 5040 24550 5092
rect 24964 5080 24992 5120
rect 25406 5108 25412 5120
rect 25464 5108 25470 5160
rect 28166 5108 28172 5160
rect 28224 5148 28230 5160
rect 28629 5151 28687 5157
rect 28629 5148 28641 5151
rect 28224 5120 28641 5148
rect 28224 5108 28230 5120
rect 28629 5117 28641 5120
rect 28675 5117 28687 5151
rect 28629 5111 28687 5117
rect 29178 5108 29184 5160
rect 29236 5148 29242 5160
rect 29656 5148 29684 5179
rect 29932 5148 29960 5179
rect 30834 5176 30840 5228
rect 30892 5176 30898 5228
rect 29236 5120 29684 5148
rect 29748 5120 29960 5148
rect 30009 5151 30067 5157
rect 29236 5108 29242 5120
rect 25958 5080 25964 5092
rect 24964 5052 25964 5080
rect 25958 5040 25964 5052
rect 26016 5040 26022 5092
rect 28905 5083 28963 5089
rect 28905 5049 28917 5083
rect 28951 5049 28963 5083
rect 28905 5043 28963 5049
rect 29089 5083 29147 5089
rect 29089 5049 29101 5083
rect 29135 5080 29147 5083
rect 29748 5080 29776 5120
rect 30009 5117 30021 5151
rect 30055 5148 30067 5151
rect 30745 5151 30803 5157
rect 30745 5148 30757 5151
rect 30055 5120 30757 5148
rect 30055 5117 30067 5120
rect 30009 5111 30067 5117
rect 30745 5117 30757 5120
rect 30791 5117 30803 5151
rect 30852 5148 30880 5176
rect 31496 5148 31524 5256
rect 31570 5176 31576 5228
rect 31628 5216 31634 5228
rect 32140 5225 32168 5256
rect 32401 5253 32413 5287
rect 32447 5284 32459 5287
rect 32447 5256 32536 5284
rect 32447 5253 32459 5256
rect 32401 5247 32459 5253
rect 32508 5225 32536 5256
rect 32125 5219 32183 5225
rect 31628 5188 32076 5216
rect 31628 5176 31634 5188
rect 31665 5151 31723 5157
rect 31665 5148 31677 5151
rect 30852 5120 31677 5148
rect 30745 5111 30803 5117
rect 31665 5117 31677 5120
rect 31711 5117 31723 5151
rect 32048 5148 32076 5188
rect 32125 5185 32137 5219
rect 32171 5185 32183 5219
rect 32125 5179 32183 5185
rect 32493 5219 32551 5225
rect 32493 5185 32505 5219
rect 32539 5185 32551 5219
rect 32600 5216 32628 5324
rect 32677 5321 32689 5355
rect 32723 5352 32735 5355
rect 32766 5352 32772 5364
rect 32723 5324 32772 5352
rect 32723 5321 32735 5324
rect 32677 5315 32735 5321
rect 32766 5312 32772 5324
rect 32824 5312 32830 5364
rect 33318 5312 33324 5364
rect 33376 5361 33382 5364
rect 33376 5355 33395 5361
rect 33383 5321 33395 5355
rect 33376 5315 33395 5321
rect 33505 5355 33563 5361
rect 33505 5321 33517 5355
rect 33551 5352 33563 5355
rect 33778 5352 33784 5364
rect 33551 5324 33784 5352
rect 33551 5321 33563 5324
rect 33505 5315 33563 5321
rect 33376 5312 33382 5315
rect 33778 5312 33784 5324
rect 33836 5312 33842 5364
rect 34609 5355 34667 5361
rect 34609 5321 34621 5355
rect 34655 5352 34667 5355
rect 34698 5352 34704 5364
rect 34655 5324 34704 5352
rect 34655 5321 34667 5324
rect 34609 5315 34667 5321
rect 34698 5312 34704 5324
rect 34756 5312 34762 5364
rect 35066 5312 35072 5364
rect 35124 5352 35130 5364
rect 35345 5355 35403 5361
rect 35345 5352 35357 5355
rect 35124 5324 35357 5352
rect 35124 5312 35130 5324
rect 35345 5321 35357 5324
rect 35391 5321 35403 5355
rect 35345 5315 35403 5321
rect 33134 5244 33140 5296
rect 33192 5284 33198 5296
rect 33873 5287 33931 5293
rect 33873 5284 33885 5287
rect 33192 5256 33885 5284
rect 33192 5244 33198 5256
rect 33873 5253 33885 5256
rect 33919 5253 33931 5287
rect 33873 5247 33931 5253
rect 32677 5219 32735 5225
rect 32677 5216 32689 5219
rect 32600 5188 32689 5216
rect 32493 5179 32551 5185
rect 32677 5185 32689 5188
rect 32723 5185 32735 5219
rect 32677 5179 32735 5185
rect 32401 5151 32459 5157
rect 32401 5148 32413 5151
rect 32048 5120 32413 5148
rect 31665 5111 31723 5117
rect 32401 5117 32413 5120
rect 32447 5117 32459 5151
rect 32401 5111 32459 5117
rect 29135 5052 29776 5080
rect 29135 5049 29147 5052
rect 29089 5043 29147 5049
rect 6546 4972 6552 5024
rect 6604 4972 6610 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 6917 5015 6975 5021
rect 6917 5012 6929 5015
rect 6880 4984 6929 5012
rect 6880 4972 6886 4984
rect 6917 4981 6929 4984
rect 6963 4981 6975 5015
rect 6917 4975 6975 4981
rect 9398 4972 9404 5024
rect 9456 4972 9462 5024
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11296 4984 11713 5012
rect 11296 4972 11302 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 12158 4972 12164 5024
rect 12216 4972 12222 5024
rect 12342 4972 12348 5024
rect 12400 4972 12406 5024
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 13173 5015 13231 5021
rect 13173 5012 13185 5015
rect 12676 4984 13185 5012
rect 12676 4972 12682 4984
rect 13173 4981 13185 4984
rect 13219 4981 13231 5015
rect 13173 4975 13231 4981
rect 22186 4972 22192 5024
rect 22244 4972 22250 5024
rect 25774 4972 25780 5024
rect 25832 4972 25838 5024
rect 28626 4972 28632 5024
rect 28684 5012 28690 5024
rect 28920 5012 28948 5043
rect 29822 5040 29828 5092
rect 29880 5040 29886 5092
rect 30760 5080 30788 5111
rect 32217 5083 32275 5089
rect 32217 5080 32229 5083
rect 30760 5052 32229 5080
rect 31588 5021 31616 5052
rect 32217 5049 32229 5052
rect 32263 5049 32275 5083
rect 32217 5043 32275 5049
rect 28684 4984 28948 5012
rect 31573 5015 31631 5021
rect 28684 4972 28690 4984
rect 31573 4981 31585 5015
rect 31619 4981 31631 5015
rect 32692 5012 32720 5179
rect 33318 5176 33324 5228
rect 33376 5216 33382 5228
rect 33597 5219 33655 5225
rect 33597 5216 33609 5219
rect 33376 5188 33609 5216
rect 33376 5176 33382 5188
rect 33597 5185 33609 5188
rect 33643 5185 33655 5219
rect 33597 5179 33655 5185
rect 33689 5219 33747 5225
rect 33689 5185 33701 5219
rect 33735 5185 33747 5219
rect 33689 5179 33747 5185
rect 33704 5080 33732 5179
rect 34146 5176 34152 5228
rect 34204 5216 34210 5228
rect 34241 5219 34299 5225
rect 34241 5216 34253 5219
rect 34204 5188 34253 5216
rect 34204 5176 34210 5188
rect 34241 5185 34253 5188
rect 34287 5185 34299 5219
rect 34241 5179 34299 5185
rect 34425 5219 34483 5225
rect 34425 5185 34437 5219
rect 34471 5185 34483 5219
rect 34425 5179 34483 5185
rect 34701 5219 34759 5225
rect 34701 5185 34713 5219
rect 34747 5216 34759 5219
rect 34790 5216 34796 5228
rect 34747 5188 34796 5216
rect 34747 5185 34759 5188
rect 34701 5179 34759 5185
rect 34054 5108 34060 5160
rect 34112 5148 34118 5160
rect 34440 5148 34468 5179
rect 34790 5176 34796 5188
rect 34848 5176 34854 5228
rect 34885 5219 34943 5225
rect 34885 5185 34897 5219
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 35161 5219 35219 5225
rect 35161 5185 35173 5219
rect 35207 5216 35219 5219
rect 35342 5216 35348 5228
rect 35207 5188 35348 5216
rect 35207 5185 35219 5188
rect 35161 5179 35219 5185
rect 34900 5148 34928 5179
rect 35342 5176 35348 5188
rect 35400 5176 35406 5228
rect 34112 5120 34928 5148
rect 34112 5108 34118 5120
rect 33336 5052 33732 5080
rect 33336 5021 33364 5052
rect 33870 5040 33876 5092
rect 33928 5040 33934 5092
rect 33321 5015 33379 5021
rect 33321 5012 33333 5015
rect 32692 4984 33333 5012
rect 31573 4975 31631 4981
rect 33321 4981 33333 4984
rect 33367 4981 33379 5015
rect 33321 4975 33379 4981
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 5994 4768 6000 4820
rect 6052 4768 6058 4820
rect 8294 4768 8300 4820
rect 8352 4768 8358 4820
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 9030 4808 9036 4820
rect 8536 4780 9036 4808
rect 8536 4768 8542 4780
rect 9030 4768 9036 4780
rect 9088 4808 9094 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9088 4780 9413 4808
rect 9088 4768 9094 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 9674 4768 9680 4820
rect 9732 4768 9738 4820
rect 10873 4811 10931 4817
rect 10873 4777 10885 4811
rect 10919 4777 10931 4811
rect 10873 4771 10931 4777
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 4157 4743 4215 4749
rect 4157 4740 4169 4743
rect 4028 4712 4169 4740
rect 4028 4700 4034 4712
rect 4157 4709 4169 4712
rect 4203 4709 4215 4743
rect 4157 4703 4215 4709
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4120 4644 4997 4672
rect 4120 4632 4126 4644
rect 4985 4641 4997 4644
rect 5031 4672 5043 4675
rect 5350 4672 5356 4684
rect 5031 4644 5356 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5350 4632 5356 4644
rect 5408 4672 5414 4684
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 5408 4644 6561 4672
rect 5408 4632 5414 4644
rect 6549 4641 6561 4644
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 6822 4632 6828 4684
rect 6880 4632 6886 4684
rect 8312 4672 8340 4768
rect 10888 4740 10916 4771
rect 11146 4768 11152 4820
rect 11204 4768 11210 4820
rect 23293 4811 23351 4817
rect 23293 4777 23305 4811
rect 23339 4808 23351 4811
rect 23474 4808 23480 4820
rect 23339 4780 23480 4808
rect 23339 4777 23351 4780
rect 23293 4771 23351 4777
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 25222 4768 25228 4820
rect 25280 4808 25286 4820
rect 25777 4811 25835 4817
rect 25777 4808 25789 4811
rect 25280 4780 25789 4808
rect 25280 4768 25286 4780
rect 25777 4777 25789 4780
rect 25823 4777 25835 4811
rect 27614 4808 27620 4820
rect 25777 4771 25835 4777
rect 26344 4780 27620 4808
rect 9600 4712 10916 4740
rect 22741 4743 22799 4749
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8312 4644 9045 4672
rect 9033 4641 9045 4644
rect 9079 4672 9091 4675
rect 9214 4672 9220 4684
rect 9079 4644 9220 4672
rect 9079 4641 9091 4644
rect 9033 4635 9091 4641
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9600 4616 9628 4712
rect 22741 4709 22753 4743
rect 22787 4709 22799 4743
rect 22741 4703 22799 4709
rect 23569 4743 23627 4749
rect 23569 4709 23581 4743
rect 23615 4740 23627 4743
rect 26234 4740 26240 4752
rect 23615 4712 26240 4740
rect 23615 4709 23627 4712
rect 23569 4703 23627 4709
rect 12158 4632 12164 4684
rect 12216 4632 12222 4684
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 15838 4672 15844 4684
rect 13955 4644 15844 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 18506 4632 18512 4684
rect 18564 4672 18570 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 18564 4644 19257 4672
rect 18564 4632 18570 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 21269 4675 21327 4681
rect 21269 4641 21281 4675
rect 21315 4672 21327 4675
rect 21726 4672 21732 4684
rect 21315 4644 21732 4672
rect 21315 4641 21327 4644
rect 21269 4635 21327 4641
rect 21726 4632 21732 4644
rect 21784 4632 21790 4684
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 3881 4607 3939 4613
rect 3881 4604 3893 4607
rect 3844 4576 3893 4604
rect 3844 4564 3850 4576
rect 3881 4573 3893 4576
rect 3927 4573 3939 4607
rect 3881 4567 3939 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4203 4576 5273 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5592 4576 5825 4604
rect 5592 4564 5598 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6086 4604 6092 4616
rect 6043 4576 6092 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 4246 4496 4252 4548
rect 4304 4496 4310 4548
rect 6288 4536 6316 4567
rect 7926 4564 7932 4616
rect 7984 4564 7990 4616
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 9582 4604 9588 4616
rect 9539 4576 9588 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 6914 4536 6920 4548
rect 6288 4508 6920 4536
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 9140 4536 9168 4567
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11330 4604 11336 4616
rect 11011 4576 11336 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 10520 4536 10548 4567
rect 8628 4508 10548 4536
rect 10612 4536 10640 4567
rect 11330 4564 11336 4576
rect 11388 4604 11394 4616
rect 12176 4604 12204 4632
rect 11388 4576 12204 4604
rect 11388 4564 11394 4576
rect 12526 4564 12532 4616
rect 12584 4564 12590 4616
rect 22278 4564 22284 4616
rect 22336 4604 22342 4616
rect 22465 4607 22523 4613
rect 22465 4604 22477 4607
rect 22336 4576 22477 4604
rect 22336 4564 22342 4576
rect 22465 4573 22477 4576
rect 22511 4573 22523 4607
rect 22756 4604 22784 4703
rect 23584 4672 23612 4703
rect 26234 4700 26240 4712
rect 26292 4700 26298 4752
rect 23308 4644 23612 4672
rect 22925 4607 22983 4613
rect 22925 4604 22937 4607
rect 22756 4576 22937 4604
rect 22465 4567 22523 4573
rect 22925 4573 22937 4576
rect 22971 4573 22983 4607
rect 23308 4604 23336 4644
rect 23750 4632 23756 4684
rect 23808 4672 23814 4684
rect 26344 4672 26372 4780
rect 27614 4768 27620 4780
rect 27672 4768 27678 4820
rect 27709 4811 27767 4817
rect 27709 4777 27721 4811
rect 27755 4808 27767 4811
rect 28905 4811 28963 4817
rect 27755 4780 28856 4808
rect 27755 4777 27767 4780
rect 27709 4771 27767 4777
rect 27065 4743 27123 4749
rect 27065 4709 27077 4743
rect 27111 4740 27123 4743
rect 27798 4740 27804 4752
rect 27111 4712 27804 4740
rect 27111 4709 27123 4712
rect 27065 4703 27123 4709
rect 27798 4700 27804 4712
rect 27856 4700 27862 4752
rect 28828 4740 28856 4780
rect 28905 4777 28917 4811
rect 28951 4808 28963 4811
rect 29362 4808 29368 4820
rect 28951 4780 29368 4808
rect 28951 4777 28963 4780
rect 28905 4771 28963 4777
rect 29362 4768 29368 4780
rect 29420 4768 29426 4820
rect 33689 4811 33747 4817
rect 33689 4777 33701 4811
rect 33735 4808 33747 4811
rect 33870 4808 33876 4820
rect 33735 4780 33876 4808
rect 33735 4777 33747 4780
rect 33689 4771 33747 4777
rect 33870 4768 33876 4780
rect 33928 4768 33934 4820
rect 34054 4768 34060 4820
rect 34112 4768 34118 4820
rect 34146 4768 34152 4820
rect 34204 4768 34210 4820
rect 35342 4768 35348 4820
rect 35400 4768 35406 4820
rect 30834 4740 30840 4752
rect 28828 4712 30840 4740
rect 30834 4700 30840 4712
rect 30892 4700 30898 4752
rect 33888 4740 33916 4768
rect 34241 4743 34299 4749
rect 34241 4740 34253 4743
rect 33888 4712 34253 4740
rect 34241 4709 34253 4712
rect 34287 4709 34299 4743
rect 34241 4703 34299 4709
rect 23808 4644 26372 4672
rect 23808 4632 23814 4644
rect 26418 4632 26424 4684
rect 26476 4672 26482 4684
rect 27525 4675 27583 4681
rect 26476 4644 27200 4672
rect 26476 4632 26482 4644
rect 22925 4567 22983 4573
rect 23032 4576 23336 4604
rect 11422 4536 11428 4548
rect 10612 4508 11428 4536
rect 8628 4496 8634 4508
rect 11422 4496 11428 4508
rect 11480 4496 11486 4548
rect 13630 4496 13636 4548
rect 13688 4496 13694 4548
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 19521 4539 19579 4545
rect 19521 4536 19533 4539
rect 13780 4508 19533 4536
rect 13780 4496 13786 4508
rect 19521 4505 19533 4508
rect 19567 4505 19579 4539
rect 19521 4499 19579 4505
rect 19978 4496 19984 4548
rect 20036 4496 20042 4548
rect 22002 4496 22008 4548
rect 22060 4536 22066 4548
rect 22060 4508 22324 4536
rect 22060 4496 22066 4508
rect 842 4428 848 4480
rect 900 4468 906 4480
rect 1397 4471 1455 4477
rect 1397 4468 1409 4471
rect 900 4440 1409 4468
rect 900 4428 906 4440
rect 1397 4437 1409 4440
rect 1443 4437 1455 4471
rect 1397 4431 1455 4437
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 4614 4468 4620 4480
rect 4019 4440 4620 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 22296 4468 22324 4508
rect 22370 4496 22376 4548
rect 22428 4536 22434 4548
rect 22738 4536 22744 4548
rect 22428 4508 22744 4536
rect 22428 4496 22434 4508
rect 22738 4496 22744 4508
rect 22796 4536 22802 4548
rect 23032 4536 23060 4576
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 23440 4576 23888 4604
rect 23440 4564 23446 4576
rect 22796 4508 23060 4536
rect 22796 4496 22802 4508
rect 23106 4496 23112 4548
rect 23164 4496 23170 4548
rect 23860 4536 23888 4576
rect 23934 4564 23940 4616
rect 23992 4564 23998 4616
rect 24121 4607 24179 4613
rect 24121 4573 24133 4607
rect 24167 4604 24179 4607
rect 24854 4604 24860 4616
rect 24167 4576 24860 4604
rect 24167 4573 24179 4576
rect 24121 4567 24179 4573
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 25314 4564 25320 4616
rect 25372 4604 25378 4616
rect 26145 4607 26203 4613
rect 26145 4604 26157 4607
rect 25372 4576 26157 4604
rect 25372 4564 25378 4576
rect 26145 4573 26157 4576
rect 26191 4604 26203 4607
rect 26694 4604 26700 4616
rect 26191 4576 26700 4604
rect 26191 4573 26203 4576
rect 26145 4567 26203 4573
rect 26694 4564 26700 4576
rect 26752 4564 26758 4616
rect 26789 4607 26847 4613
rect 26789 4573 26801 4607
rect 26835 4604 26847 4607
rect 26878 4604 26884 4616
rect 26835 4576 26884 4604
rect 26835 4573 26847 4576
rect 26789 4567 26847 4573
rect 26878 4564 26884 4576
rect 26936 4564 26942 4616
rect 26970 4536 26976 4548
rect 23860 4508 26976 4536
rect 26970 4496 26976 4508
rect 27028 4496 27034 4548
rect 27065 4539 27123 4545
rect 27065 4505 27077 4539
rect 27111 4505 27123 4539
rect 27172 4536 27200 4644
rect 27525 4641 27537 4675
rect 27571 4672 27583 4675
rect 27890 4672 27896 4684
rect 27571 4644 27896 4672
rect 27571 4641 27583 4644
rect 27525 4635 27583 4641
rect 27890 4632 27896 4644
rect 27948 4632 27954 4684
rect 28626 4632 28632 4684
rect 28684 4632 28690 4684
rect 33502 4632 33508 4684
rect 33560 4672 33566 4684
rect 33597 4675 33655 4681
rect 33597 4672 33609 4675
rect 33560 4644 33609 4672
rect 33560 4632 33566 4644
rect 33597 4641 33609 4644
rect 33643 4672 33655 4675
rect 34425 4675 34483 4681
rect 34425 4672 34437 4675
rect 33643 4644 34437 4672
rect 33643 4641 33655 4644
rect 33597 4635 33655 4641
rect 34425 4641 34437 4644
rect 34471 4641 34483 4675
rect 34425 4635 34483 4641
rect 27430 4564 27436 4616
rect 27488 4564 27494 4616
rect 28166 4564 28172 4616
rect 28224 4604 28230 4616
rect 28537 4607 28595 4613
rect 28537 4604 28549 4607
rect 28224 4576 28549 4604
rect 28224 4564 28230 4576
rect 28537 4573 28549 4576
rect 28583 4573 28595 4607
rect 28537 4567 28595 4573
rect 33410 4564 33416 4616
rect 33468 4604 33474 4616
rect 33873 4607 33931 4613
rect 33873 4604 33885 4607
rect 33468 4576 33885 4604
rect 33468 4564 33474 4576
rect 33873 4573 33885 4576
rect 33919 4604 33931 4607
rect 34149 4607 34207 4613
rect 34149 4604 34161 4607
rect 33919 4576 34161 4604
rect 33919 4573 33931 4576
rect 33873 4567 33931 4573
rect 34149 4573 34161 4576
rect 34195 4573 34207 4607
rect 34149 4567 34207 4573
rect 34790 4564 34796 4616
rect 34848 4604 34854 4616
rect 35069 4607 35127 4613
rect 35069 4604 35081 4607
rect 34848 4576 35081 4604
rect 34848 4564 34854 4576
rect 35069 4573 35081 4576
rect 35115 4573 35127 4607
rect 35069 4567 35127 4573
rect 35161 4607 35219 4613
rect 35161 4573 35173 4607
rect 35207 4573 35219 4607
rect 35161 4567 35219 4573
rect 27522 4536 27528 4548
rect 27172 4508 27528 4536
rect 27065 4499 27123 4505
rect 22557 4471 22615 4477
rect 22557 4468 22569 4471
rect 22296 4440 22569 4468
rect 22557 4437 22569 4440
rect 22603 4468 22615 4471
rect 23750 4468 23756 4480
rect 22603 4440 23756 4468
rect 22603 4437 22615 4440
rect 22557 4431 22615 4437
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 23842 4428 23848 4480
rect 23900 4468 23906 4480
rect 24029 4471 24087 4477
rect 24029 4468 24041 4471
rect 23900 4440 24041 4468
rect 23900 4428 23906 4440
rect 24029 4437 24041 4440
rect 24075 4437 24087 4471
rect 24029 4431 24087 4437
rect 26234 4428 26240 4480
rect 26292 4428 26298 4480
rect 26602 4428 26608 4480
rect 26660 4468 26666 4480
rect 26881 4471 26939 4477
rect 26881 4468 26893 4471
rect 26660 4440 26893 4468
rect 26660 4428 26666 4440
rect 26881 4437 26893 4440
rect 26927 4437 26939 4471
rect 27080 4468 27108 4499
rect 27522 4496 27528 4508
rect 27580 4496 27586 4548
rect 27614 4496 27620 4548
rect 27672 4536 27678 4548
rect 28718 4536 28724 4548
rect 27672 4508 28724 4536
rect 27672 4496 27678 4508
rect 28718 4496 28724 4508
rect 28776 4496 28782 4548
rect 34054 4496 34060 4548
rect 34112 4536 34118 4548
rect 35176 4536 35204 4567
rect 34112 4508 35204 4536
rect 34112 4496 34118 4508
rect 27246 4468 27252 4480
rect 27080 4440 27252 4468
rect 26881 4431 26939 4437
rect 27246 4428 27252 4440
rect 27304 4468 27310 4480
rect 28074 4468 28080 4480
rect 27304 4440 28080 4468
rect 27304 4428 27310 4440
rect 28074 4428 28080 4440
rect 28132 4428 28138 4480
rect 34698 4428 34704 4480
rect 34756 4428 34762 4480
rect 1104 4378 38824 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 38824 4378
rect 1104 4304 38824 4326
rect 4154 4264 4160 4276
rect 3344 4236 4160 4264
rect 3344 4196 3372 4236
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 4304 4236 5365 4264
rect 4304 4224 4310 4236
rect 5353 4233 5365 4236
rect 5399 4264 5411 4267
rect 10410 4264 10416 4276
rect 5399 4236 10416 4264
rect 5399 4233 5411 4236
rect 5353 4227 5411 4233
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 10949 4267 11007 4273
rect 10949 4233 10961 4267
rect 10995 4264 11007 4267
rect 12342 4264 12348 4276
rect 10995 4236 12348 4264
rect 10995 4233 11007 4236
rect 10949 4227 11007 4233
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 12529 4267 12587 4273
rect 12529 4233 12541 4267
rect 12575 4264 12587 4267
rect 13630 4264 13636 4276
rect 12575 4236 13636 4264
rect 12575 4233 12587 4236
rect 12529 4227 12587 4233
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 22278 4224 22284 4276
rect 22336 4264 22342 4276
rect 22389 4267 22447 4273
rect 22389 4264 22401 4267
rect 22336 4236 22401 4264
rect 22336 4224 22342 4236
rect 22389 4233 22401 4236
rect 22435 4233 22447 4267
rect 22389 4227 22447 4233
rect 22557 4267 22615 4273
rect 22557 4233 22569 4267
rect 22603 4264 22615 4267
rect 23106 4264 23112 4276
rect 22603 4236 23112 4264
rect 22603 4233 22615 4236
rect 22557 4227 22615 4233
rect 23106 4224 23112 4236
rect 23164 4264 23170 4276
rect 24302 4264 24308 4276
rect 23164 4236 24308 4264
rect 23164 4224 23170 4236
rect 24302 4224 24308 4236
rect 24360 4224 24366 4276
rect 25406 4224 25412 4276
rect 25464 4264 25470 4276
rect 26145 4267 26203 4273
rect 25464 4236 25912 4264
rect 25464 4224 25470 4236
rect 4798 4196 4804 4208
rect 3252 4168 3372 4196
rect 4738 4168 4804 4196
rect 3252 4137 3280 4168
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 11149 4199 11207 4205
rect 11149 4165 11161 4199
rect 11195 4196 11207 4199
rect 11422 4196 11428 4208
rect 11195 4168 11428 4196
rect 11195 4165 11207 4168
rect 11149 4159 11207 4165
rect 11422 4156 11428 4168
rect 11480 4196 11486 4208
rect 12158 4196 12164 4208
rect 11480 4168 12164 4196
rect 11480 4156 11486 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 22002 4156 22008 4208
rect 22060 4196 22066 4208
rect 22189 4199 22247 4205
rect 22189 4196 22201 4199
rect 22060 4168 22201 4196
rect 22060 4156 22066 4168
rect 22189 4165 22201 4168
rect 22235 4165 22247 4199
rect 22189 4159 22247 4165
rect 23216 4168 23428 4196
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 5810 4128 5816 4140
rect 5767 4100 5816 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 5994 4128 6000 4140
rect 5951 4100 6000 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6362 4088 6368 4140
rect 6420 4088 6426 4140
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 7098 4128 7104 4140
rect 6687 4100 7104 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7616 4100 7665 4128
rect 7616 4088 7622 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7834 4088 7840 4140
rect 7892 4088 7898 4140
rect 8570 4088 8576 4140
rect 8628 4088 8634 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4128 8815 4131
rect 10321 4131 10379 4137
rect 8803 4100 9720 4128
rect 8803 4097 8815 4100
rect 8757 4091 8815 4097
rect 3510 4020 3516 4072
rect 3568 4020 3574 4072
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 6457 4063 6515 4069
rect 6457 4060 6469 4063
rect 5592 4032 6469 4060
rect 5592 4020 5598 4032
rect 6457 4029 6469 4032
rect 6503 4029 6515 4063
rect 6457 4023 6515 4029
rect 9692 4004 9720 4100
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 6825 3995 6883 4001
rect 6825 3961 6837 3995
rect 6871 3992 6883 3995
rect 9490 3992 9496 4004
rect 6871 3964 9496 3992
rect 6871 3961 6883 3964
rect 6825 3955 6883 3961
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 9674 3952 9680 4004
rect 9732 3992 9738 4004
rect 10336 3992 10364 4091
rect 10520 4060 10548 4091
rect 11514 4088 11520 4140
rect 11572 4088 11578 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 11882 4128 11888 4140
rect 11747 4100 11888 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 12400 4100 12449 4128
rect 12400 4088 12406 4100
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12618 4088 12624 4140
rect 12676 4088 12682 4140
rect 21726 4088 21732 4140
rect 21784 4128 21790 4140
rect 22097 4131 22155 4137
rect 22097 4128 22109 4131
rect 21784 4100 22109 4128
rect 21784 4088 21790 4100
rect 22097 4097 22109 4100
rect 22143 4097 22155 4131
rect 23216 4128 23244 4168
rect 22097 4091 22155 4097
rect 22848 4100 23244 4128
rect 23293 4131 23351 4137
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 10520 4032 11621 4060
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 21818 4020 21824 4072
rect 21876 4060 21882 4072
rect 22005 4063 22063 4069
rect 22005 4060 22017 4063
rect 21876 4032 22017 4060
rect 21876 4020 21882 4032
rect 22005 4029 22017 4032
rect 22051 4060 22063 4063
rect 22848 4060 22876 4100
rect 23293 4097 23305 4131
rect 23339 4097 23351 4131
rect 23400 4128 23428 4168
rect 23842 4156 23848 4208
rect 23900 4156 23906 4208
rect 23934 4156 23940 4208
rect 23992 4196 23998 4208
rect 25133 4199 25191 4205
rect 23992 4168 24624 4196
rect 23992 4156 23998 4168
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 23400 4100 23673 4128
rect 23293 4091 23351 4097
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 23661 4091 23719 4097
rect 23753 4131 23811 4137
rect 23753 4097 23765 4131
rect 23799 4128 23811 4131
rect 23799 4100 23980 4128
rect 23799 4097 23811 4100
rect 23753 4091 23811 4097
rect 22051 4032 22876 4060
rect 23308 4060 23336 4091
rect 23952 4060 23980 4100
rect 24026 4088 24032 4140
rect 24084 4088 24090 4140
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24394 4128 24400 4140
rect 24351 4100 24400 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 24394 4088 24400 4100
rect 24452 4088 24458 4140
rect 23308 4032 23796 4060
rect 23952 4032 24164 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 23768 4004 23796 4032
rect 24136 4004 24164 4032
rect 10781 3995 10839 4001
rect 10781 3992 10793 3995
rect 9732 3964 10793 3992
rect 9732 3952 9738 3964
rect 10781 3961 10793 3964
rect 10827 3961 10839 3995
rect 10781 3955 10839 3961
rect 23750 3952 23756 4004
rect 23808 3952 23814 4004
rect 24118 3952 24124 4004
rect 24176 3952 24182 4004
rect 24596 4001 24624 4168
rect 25133 4165 25145 4199
rect 25179 4196 25191 4199
rect 25774 4196 25780 4208
rect 25179 4168 25780 4196
rect 25179 4165 25191 4168
rect 25133 4159 25191 4165
rect 25774 4156 25780 4168
rect 25832 4156 25838 4208
rect 25884 4196 25912 4236
rect 26145 4233 26157 4267
rect 26191 4264 26203 4267
rect 26234 4264 26240 4276
rect 26191 4236 26240 4264
rect 26191 4233 26203 4236
rect 26145 4227 26203 4233
rect 26234 4224 26240 4236
rect 26292 4224 26298 4276
rect 26326 4224 26332 4276
rect 26384 4264 26390 4276
rect 27246 4264 27252 4276
rect 26384 4236 27252 4264
rect 26384 4224 26390 4236
rect 26436 4205 26464 4236
rect 27246 4224 27252 4236
rect 27304 4224 27310 4276
rect 27341 4267 27399 4273
rect 27341 4233 27353 4267
rect 27387 4264 27399 4267
rect 27387 4236 28120 4264
rect 27387 4233 27399 4236
rect 27341 4227 27399 4233
rect 26421 4199 26479 4205
rect 25884 4168 26280 4196
rect 24765 4131 24823 4137
rect 24765 4097 24777 4131
rect 24811 4097 24823 4131
rect 24765 4091 24823 4097
rect 24581 3995 24639 4001
rect 24581 3961 24593 3995
rect 24627 3992 24639 3995
rect 24670 3992 24676 4004
rect 24627 3964 24676 3992
rect 24627 3961 24639 3964
rect 24581 3955 24639 3961
rect 24670 3952 24676 3964
rect 24728 3952 24734 4004
rect 24780 3992 24808 4091
rect 25314 4088 25320 4140
rect 25372 4088 25378 4140
rect 25501 4131 25559 4137
rect 25501 4097 25513 4131
rect 25547 4128 25559 4131
rect 25682 4128 25688 4140
rect 25547 4100 25688 4128
rect 25547 4097 25559 4100
rect 25501 4091 25559 4097
rect 25682 4088 25688 4100
rect 25740 4088 25746 4140
rect 26145 4131 26203 4137
rect 26145 4097 26157 4131
rect 26191 4097 26203 4131
rect 26145 4091 26203 4097
rect 24854 4020 24860 4072
rect 24912 4020 24918 4072
rect 25038 4020 25044 4072
rect 25096 4020 25102 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 26160 4060 26188 4091
rect 25271 4032 26188 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25501 3995 25559 4001
rect 25501 3992 25513 3995
rect 24780 3964 25513 3992
rect 25501 3961 25513 3964
rect 25547 3961 25559 3995
rect 25501 3955 25559 3961
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 5534 3924 5540 3936
rect 5040 3896 5540 3924
rect 5040 3884 5046 3896
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5684 3896 5733 3924
rect 5684 3884 5690 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 6546 3884 6552 3936
rect 6604 3884 6610 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7340 3896 7849 3924
rect 7340 3884 7346 3896
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 7837 3887 7895 3893
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 9950 3924 9956 3936
rect 8803 3896 9956 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10502 3884 10508 3936
rect 10560 3884 10566 3936
rect 10962 3884 10968 3936
rect 11020 3884 11026 3936
rect 22370 3884 22376 3936
rect 22428 3884 22434 3936
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 23477 3927 23535 3933
rect 23477 3924 23489 3927
rect 22796 3896 23489 3924
rect 22796 3884 22802 3896
rect 23477 3893 23489 3896
rect 23523 3893 23535 3927
rect 26160 3924 26188 4032
rect 26252 3992 26280 4168
rect 26421 4165 26433 4199
rect 26467 4165 26479 4199
rect 26637 4199 26695 4205
rect 26637 4196 26649 4199
rect 26421 4159 26479 4165
rect 26620 4165 26649 4196
rect 26683 4196 26695 4199
rect 26878 4196 26884 4208
rect 26683 4168 26884 4196
rect 26683 4165 26695 4168
rect 26620 4159 26695 4165
rect 26329 4131 26387 4137
rect 26329 4097 26341 4131
rect 26375 4128 26387 4131
rect 26620 4128 26648 4159
rect 26878 4156 26884 4168
rect 26936 4156 26942 4208
rect 27798 4156 27804 4208
rect 27856 4156 27862 4208
rect 28092 4196 28120 4236
rect 28166 4224 28172 4276
rect 28224 4224 28230 4276
rect 28626 4224 28632 4276
rect 28684 4264 28690 4276
rect 28905 4267 28963 4273
rect 28905 4264 28917 4267
rect 28684 4236 28917 4264
rect 28684 4224 28690 4236
rect 28905 4233 28917 4236
rect 28951 4233 28963 4267
rect 28905 4227 28963 4233
rect 31570 4224 31576 4276
rect 31628 4264 31634 4276
rect 31665 4267 31723 4273
rect 31665 4264 31677 4267
rect 31628 4236 31677 4264
rect 31628 4224 31634 4236
rect 31665 4233 31677 4236
rect 31711 4233 31723 4267
rect 33410 4264 33416 4276
rect 31665 4227 31723 4233
rect 32416 4236 33416 4264
rect 30834 4196 30840 4208
rect 28092 4168 30840 4196
rect 30834 4156 30840 4168
rect 30892 4196 30898 4208
rect 32416 4196 32444 4236
rect 33410 4224 33416 4236
rect 33468 4224 33474 4276
rect 33502 4224 33508 4276
rect 33560 4224 33566 4276
rect 30892 4168 31524 4196
rect 30892 4156 30898 4168
rect 31496 4140 31524 4168
rect 31680 4168 32444 4196
rect 26375 4100 26648 4128
rect 27985 4131 28043 4137
rect 26375 4097 26387 4100
rect 26329 4091 26387 4097
rect 27985 4097 27997 4131
rect 28031 4097 28043 4131
rect 27985 4091 28043 4097
rect 27433 4063 27491 4069
rect 27433 4029 27445 4063
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 26789 3995 26847 4001
rect 26252 3964 26740 3992
rect 26602 3924 26608 3936
rect 26160 3896 26608 3924
rect 23477 3887 23535 3893
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 26712 3924 26740 3964
rect 26789 3961 26801 3995
rect 26835 3992 26847 3995
rect 27448 3992 27476 4023
rect 27522 4020 27528 4072
rect 27580 4020 27586 4072
rect 27706 3992 27712 4004
rect 26835 3964 27384 3992
rect 27448 3964 27712 3992
rect 26835 3961 26847 3964
rect 26789 3955 26847 3961
rect 26973 3927 27031 3933
rect 26973 3924 26985 3927
rect 26712 3896 26985 3924
rect 26973 3893 26985 3896
rect 27019 3893 27031 3927
rect 27356 3924 27384 3964
rect 27706 3952 27712 3964
rect 27764 3952 27770 4004
rect 27614 3924 27620 3936
rect 27356 3896 27620 3924
rect 26973 3887 27031 3893
rect 27614 3884 27620 3896
rect 27672 3924 27678 3936
rect 28000 3924 28028 4091
rect 29546 4088 29552 4140
rect 29604 4128 29610 4140
rect 29641 4131 29699 4137
rect 29641 4128 29653 4131
rect 29604 4100 29653 4128
rect 29604 4088 29610 4100
rect 29641 4097 29653 4100
rect 29687 4097 29699 4131
rect 29641 4091 29699 4097
rect 29822 4088 29828 4140
rect 29880 4088 29886 4140
rect 31021 4131 31079 4137
rect 31021 4097 31033 4131
rect 31067 4097 31079 4131
rect 31021 4091 31079 4097
rect 29086 4020 29092 4072
rect 29144 4020 29150 4072
rect 29178 4020 29184 4072
rect 29236 4060 29242 4072
rect 30745 4063 30803 4069
rect 30745 4060 30757 4063
rect 29236 4032 30757 4060
rect 29236 4020 29242 4032
rect 30745 4029 30757 4032
rect 30791 4060 30803 4063
rect 30926 4060 30932 4072
rect 30791 4032 30932 4060
rect 30791 4029 30803 4032
rect 30745 4023 30803 4029
rect 30926 4020 30932 4032
rect 30984 4020 30990 4072
rect 28994 3952 29000 4004
rect 29052 3992 29058 4004
rect 29733 3995 29791 4001
rect 29733 3992 29745 3995
rect 29052 3964 29745 3992
rect 29052 3952 29058 3964
rect 29733 3961 29745 3964
rect 29779 3961 29791 3995
rect 31036 3992 31064 4091
rect 31110 4088 31116 4140
rect 31168 4128 31174 4140
rect 31297 4131 31355 4137
rect 31297 4128 31309 4131
rect 31168 4100 31309 4128
rect 31168 4088 31174 4100
rect 31297 4097 31309 4100
rect 31343 4097 31355 4131
rect 31297 4091 31355 4097
rect 31478 4088 31484 4140
rect 31536 4088 31542 4140
rect 31570 4088 31576 4140
rect 31628 4088 31634 4140
rect 31205 4063 31263 4069
rect 31205 4029 31217 4063
rect 31251 4060 31263 4063
rect 31680 4060 31708 4168
rect 31757 4131 31815 4137
rect 31757 4097 31769 4131
rect 31803 4128 31815 4131
rect 32030 4128 32036 4140
rect 31803 4100 32036 4128
rect 31803 4097 31815 4100
rect 31757 4091 31815 4097
rect 32030 4088 32036 4100
rect 32088 4128 32094 4140
rect 32616 4134 32674 4137
rect 32416 4131 32674 4134
rect 32416 4128 32628 4131
rect 32088 4106 32628 4128
rect 32088 4100 32444 4106
rect 32600 4100 32628 4106
rect 32088 4088 32094 4100
rect 32616 4097 32628 4100
rect 32662 4128 32674 4131
rect 33045 4131 33103 4137
rect 33045 4128 33057 4131
rect 32662 4100 33057 4128
rect 32662 4097 32674 4100
rect 32616 4091 32674 4097
rect 33045 4097 33057 4100
rect 33091 4097 33103 4131
rect 33045 4091 33103 4097
rect 31251 4032 31708 4060
rect 31251 4029 31263 4032
rect 31205 4023 31263 4029
rect 32306 4020 32312 4072
rect 32364 4060 32370 4072
rect 32493 4063 32551 4069
rect 32493 4060 32505 4063
rect 32364 4032 32505 4060
rect 32364 4020 32370 4032
rect 32493 4029 32505 4032
rect 32539 4029 32551 4063
rect 32493 4023 32551 4029
rect 32953 4063 33011 4069
rect 32953 4029 32965 4063
rect 32999 4060 33011 4063
rect 33134 4060 33140 4072
rect 32999 4032 33140 4060
rect 32999 4029 33011 4032
rect 32953 4023 33011 4029
rect 31389 3995 31447 4001
rect 31389 3992 31401 3995
rect 31036 3964 31401 3992
rect 29733 3955 29791 3961
rect 31389 3961 31401 3964
rect 31435 3992 31447 3995
rect 32508 3992 32536 4023
rect 33134 4020 33140 4032
rect 33192 4020 33198 4072
rect 33321 3995 33379 4001
rect 33321 3992 33333 3995
rect 31435 3964 31754 3992
rect 32508 3964 33333 3992
rect 31435 3961 31447 3964
rect 31389 3955 31447 3961
rect 27672 3896 28028 3924
rect 27672 3884 27678 3896
rect 28166 3884 28172 3936
rect 28224 3924 28230 3936
rect 30650 3924 30656 3936
rect 28224 3896 30656 3924
rect 28224 3884 28230 3896
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 30837 3927 30895 3933
rect 30837 3893 30849 3927
rect 30883 3924 30895 3927
rect 31110 3924 31116 3936
rect 30883 3896 31116 3924
rect 30883 3893 30895 3896
rect 30837 3887 30895 3893
rect 31110 3884 31116 3896
rect 31168 3884 31174 3936
rect 31726 3924 31754 3964
rect 33321 3961 33333 3964
rect 33367 3961 33379 3995
rect 33321 3955 33379 3961
rect 34698 3924 34704 3936
rect 31726 3896 34704 3924
rect 34698 3884 34704 3896
rect 34756 3884 34762 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3568 3692 3801 3720
rect 3568 3680 3574 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 3789 3683 3847 3689
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 3936 3692 4077 3720
rect 3936 3680 3942 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 4614 3720 4620 3732
rect 4295 3692 4620 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 6086 3720 6092 3732
rect 4856 3692 6092 3720
rect 4856 3680 4862 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 7098 3680 7104 3732
rect 7156 3680 7162 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7892 3692 7941 3720
rect 7892 3680 7898 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 8478 3680 8484 3732
rect 8536 3680 8542 3732
rect 9950 3680 9956 3732
rect 10008 3680 10014 3732
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11514 3720 11520 3732
rect 10919 3692 11520 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 22833 3723 22891 3729
rect 22833 3689 22845 3723
rect 22879 3720 22891 3723
rect 23382 3720 23388 3732
rect 22879 3692 23388 3720
rect 22879 3689 22891 3692
rect 22833 3683 22891 3689
rect 23382 3680 23388 3692
rect 23440 3680 23446 3732
rect 23566 3680 23572 3732
rect 23624 3720 23630 3732
rect 23937 3723 23995 3729
rect 23937 3720 23949 3723
rect 23624 3692 23949 3720
rect 23624 3680 23630 3692
rect 842 3612 848 3664
rect 900 3652 906 3664
rect 1397 3655 1455 3661
rect 1397 3652 1409 3655
rect 900 3624 1409 3652
rect 900 3612 906 3624
rect 1397 3621 1409 3624
rect 1443 3621 1455 3655
rect 1397 3615 1455 3621
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 8297 3655 8355 3661
rect 8297 3652 8309 3655
rect 7616 3624 8309 3652
rect 7616 3612 7622 3624
rect 8297 3621 8309 3624
rect 8343 3621 8355 3655
rect 8297 3615 8355 3621
rect 9582 3612 9588 3664
rect 9640 3652 9646 3664
rect 10962 3652 10968 3664
rect 9640 3624 10968 3652
rect 9640 3612 9646 3624
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 5350 3584 5356 3596
rect 4212 3556 5356 3584
rect 4212 3544 4218 3556
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 5626 3544 5632 3596
rect 5684 3544 5690 3596
rect 8220 3556 9076 3584
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 3878 3516 3884 3528
rect 3835 3488 3884 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 4672 3488 5089 3516
rect 4672 3476 4678 3488
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4982 3448 4988 3460
rect 4479 3420 4988 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 5092 3448 5120 3479
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 8220 3525 8248 3556
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7156 3488 7757 3516
rect 7156 3476 7162 3488
rect 7745 3485 7757 3488
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8352 3488 8708 3516
rect 8352 3476 8358 3488
rect 8680 3460 8708 3488
rect 5626 3448 5632 3460
rect 5092 3420 5632 3448
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 6086 3408 6092 3460
rect 6144 3408 6150 3460
rect 7929 3451 7987 3457
rect 7929 3417 7941 3451
rect 7975 3448 7987 3451
rect 8570 3448 8576 3460
rect 7975 3420 8576 3448
rect 7975 3417 7987 3420
rect 7929 3411 7987 3417
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 8662 3408 8668 3460
rect 8720 3408 8726 3460
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 3970 3380 3976 3392
rect 3844 3352 3976 3380
rect 3844 3340 3850 3352
rect 3970 3340 3976 3352
rect 4028 3380 4034 3392
rect 4223 3383 4281 3389
rect 4223 3380 4235 3383
rect 4028 3352 4235 3380
rect 4028 3340 4034 3352
rect 4223 3349 4235 3352
rect 4269 3349 4281 3383
rect 4223 3343 4281 3349
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 5644 3380 5672 3408
rect 6362 3380 6368 3392
rect 5644 3352 6368 3380
rect 6362 3340 6368 3352
rect 6420 3340 6426 3392
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 8113 3383 8171 3389
rect 8113 3349 8125 3383
rect 8159 3380 8171 3383
rect 8294 3380 8300 3392
rect 8159 3352 8300 3380
rect 8159 3349 8171 3352
rect 8113 3343 8171 3349
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 8465 3383 8523 3389
rect 8465 3349 8477 3383
rect 8511 3380 8523 3383
rect 8772 3380 8800 3556
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8904 3488 8953 3516
rect 8904 3476 8910 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 9048 3516 9076 3556
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 10244 3593 10272 3624
rect 10962 3612 10968 3624
rect 11020 3612 11026 3664
rect 11238 3652 11244 3664
rect 11072 3624 11244 3652
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 9272 3556 10149 3584
rect 9272 3544 9278 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3553 10287 3587
rect 10229 3547 10287 3553
rect 9674 3516 9680 3528
rect 9048 3488 9680 3516
rect 8941 3479 8999 3485
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 11072 3525 11100 3624
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11793 3587 11851 3593
rect 11195 3556 11560 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11532 3525 11560 3556
rect 11793 3553 11805 3587
rect 11839 3584 11851 3587
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 11839 3556 12357 3584
rect 11839 3553 11851 3556
rect 11793 3547 11851 3553
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3584 21143 3587
rect 21131 3556 23152 3584
rect 21131 3553 21143 3556
rect 21085 3547 21143 3553
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10091 3488 11069 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3485 11575 3519
rect 11517 3479 11575 3485
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11747 3488 12081 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 11256 3448 11284 3479
rect 11882 3448 11888 3460
rect 11256 3420 11888 3448
rect 11882 3408 11888 3420
rect 11940 3408 11946 3460
rect 12084 3448 12112 3479
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12216 3488 13001 3516
rect 12216 3476 12222 3488
rect 12989 3485 13001 3488
rect 13035 3516 13047 3519
rect 13262 3516 13268 3528
rect 13035 3488 13268 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 12342 3448 12348 3460
rect 12084 3420 12348 3448
rect 12342 3408 12348 3420
rect 12400 3408 12406 3460
rect 21361 3451 21419 3457
rect 21361 3417 21373 3451
rect 21407 3417 21419 3451
rect 22646 3448 22652 3460
rect 22586 3420 22652 3448
rect 21361 3411 21419 3417
rect 8511 3352 8800 3380
rect 9585 3383 9643 3389
rect 8511 3349 8523 3352
rect 8465 3343 8523 3349
rect 9585 3349 9597 3383
rect 9631 3380 9643 3383
rect 9769 3383 9827 3389
rect 9769 3380 9781 3383
rect 9631 3352 9781 3380
rect 9631 3349 9643 3352
rect 9585 3343 9643 3349
rect 9769 3349 9781 3352
rect 9815 3349 9827 3383
rect 9769 3343 9827 3349
rect 11333 3383 11391 3389
rect 11333 3349 11345 3383
rect 11379 3380 11391 3383
rect 11790 3380 11796 3392
rect 11379 3352 11796 3380
rect 11379 3349 11391 3352
rect 11333 3343 11391 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 21376 3380 21404 3411
rect 22646 3408 22652 3420
rect 22704 3448 22710 3460
rect 23014 3448 23020 3460
rect 22704 3420 23020 3448
rect 22704 3408 22710 3420
rect 23014 3408 23020 3420
rect 23072 3408 23078 3460
rect 23124 3457 23152 3556
rect 23860 3525 23888 3692
rect 23937 3689 23949 3692
rect 23983 3689 23995 3723
rect 23937 3683 23995 3689
rect 24026 3680 24032 3732
rect 24084 3720 24090 3732
rect 25041 3723 25099 3729
rect 25041 3720 25053 3723
rect 24084 3692 25053 3720
rect 24084 3680 24090 3692
rect 25041 3689 25053 3692
rect 25087 3689 25099 3723
rect 25041 3683 25099 3689
rect 25406 3680 25412 3732
rect 25464 3680 25470 3732
rect 27890 3680 27896 3732
rect 27948 3680 27954 3732
rect 29181 3723 29239 3729
rect 29181 3689 29193 3723
rect 29227 3720 29239 3723
rect 29822 3720 29828 3732
rect 29227 3692 29828 3720
rect 29227 3689 29239 3692
rect 29181 3683 29239 3689
rect 29822 3680 29828 3692
rect 29880 3680 29886 3732
rect 30282 3720 30288 3732
rect 29932 3692 30288 3720
rect 24854 3612 24860 3664
rect 24912 3652 24918 3664
rect 25961 3655 26019 3661
rect 25961 3652 25973 3655
rect 24912 3624 25973 3652
rect 24912 3612 24918 3624
rect 25961 3621 25973 3624
rect 26007 3621 26019 3655
rect 25961 3615 26019 3621
rect 27617 3655 27675 3661
rect 27617 3621 27629 3655
rect 27663 3621 27675 3655
rect 27617 3615 27675 3621
rect 28629 3655 28687 3661
rect 28629 3621 28641 3655
rect 28675 3652 28687 3655
rect 29546 3652 29552 3664
rect 28675 3624 29552 3652
rect 28675 3621 28687 3624
rect 28629 3615 28687 3621
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 24573 3587 24631 3593
rect 24573 3584 24585 3587
rect 24360 3556 24585 3584
rect 24360 3544 24366 3556
rect 24573 3553 24585 3556
rect 24619 3553 24631 3587
rect 24573 3547 24631 3553
rect 24762 3544 24768 3596
rect 24820 3544 24826 3596
rect 25314 3584 25320 3596
rect 24877 3559 25320 3584
rect 24857 3556 25320 3559
rect 24857 3553 24915 3556
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 24486 3476 24492 3528
rect 24544 3516 24550 3528
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 24544 3488 24685 3516
rect 24544 3476 24550 3488
rect 24673 3485 24685 3488
rect 24719 3516 24731 3519
rect 24857 3519 24869 3553
rect 24903 3519 24915 3553
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 26878 3544 26884 3596
rect 26936 3584 26942 3596
rect 27632 3584 27660 3615
rect 29546 3612 29552 3624
rect 29604 3612 29610 3664
rect 29730 3612 29736 3664
rect 29788 3652 29794 3664
rect 29932 3652 29960 3692
rect 30282 3680 30288 3692
rect 30340 3680 30346 3732
rect 30650 3680 30656 3732
rect 30708 3720 30714 3732
rect 31018 3720 31024 3732
rect 30708 3692 31024 3720
rect 30708 3680 30714 3692
rect 29788 3624 29960 3652
rect 30009 3655 30067 3661
rect 29788 3612 29794 3624
rect 30009 3621 30021 3655
rect 30055 3652 30067 3655
rect 30742 3652 30748 3664
rect 30055 3624 30748 3652
rect 30055 3621 30067 3624
rect 30009 3615 30067 3621
rect 30742 3612 30748 3624
rect 30800 3612 30806 3664
rect 30558 3584 30564 3596
rect 26936 3556 27384 3584
rect 27632 3556 30564 3584
rect 26936 3544 26942 3556
rect 24719 3488 24809 3516
rect 24857 3513 24915 3519
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 24781 3482 24809 3488
rect 24964 3488 25237 3516
rect 24964 3482 24992 3488
rect 23109 3451 23167 3457
rect 23109 3417 23121 3451
rect 23155 3448 23167 3451
rect 23750 3448 23756 3460
rect 23155 3420 23756 3448
rect 23155 3417 23167 3420
rect 23109 3411 23167 3417
rect 23750 3408 23756 3420
rect 23808 3408 23814 3460
rect 24781 3454 24992 3482
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3485 25559 3519
rect 25501 3479 25559 3485
rect 25038 3408 25044 3460
rect 25096 3448 25102 3460
rect 25516 3448 25544 3479
rect 25682 3476 25688 3528
rect 25740 3516 25746 3528
rect 25777 3519 25835 3525
rect 25777 3516 25789 3519
rect 25740 3488 25789 3516
rect 25740 3476 25746 3488
rect 25777 3485 25789 3488
rect 25823 3516 25835 3519
rect 26053 3519 26111 3525
rect 26053 3516 26065 3519
rect 25823 3488 26065 3516
rect 25823 3485 25835 3488
rect 25777 3479 25835 3485
rect 26053 3485 26065 3488
rect 26099 3485 26111 3519
rect 26053 3479 26111 3485
rect 26234 3476 26240 3528
rect 26292 3476 26298 3528
rect 26418 3476 26424 3528
rect 26476 3516 26482 3528
rect 26476 3488 26740 3516
rect 26476 3476 26482 3488
rect 25096 3420 25544 3448
rect 25096 3408 25102 3420
rect 25590 3408 25596 3460
rect 25648 3408 25654 3460
rect 26712 3457 26740 3488
rect 26970 3476 26976 3528
rect 27028 3476 27034 3528
rect 27356 3525 27384 3556
rect 30558 3544 30564 3556
rect 30616 3544 30622 3596
rect 30852 3584 30880 3692
rect 31018 3680 31024 3692
rect 31076 3680 31082 3732
rect 31110 3680 31116 3732
rect 31168 3720 31174 3732
rect 31168 3692 31248 3720
rect 31168 3680 31174 3692
rect 31220 3652 31248 3692
rect 31294 3680 31300 3732
rect 31352 3720 31358 3732
rect 31665 3723 31723 3729
rect 31665 3720 31677 3723
rect 31352 3692 31677 3720
rect 31352 3680 31358 3692
rect 31665 3689 31677 3692
rect 31711 3689 31723 3723
rect 31665 3683 31723 3689
rect 32030 3680 32036 3732
rect 32088 3680 32094 3732
rect 32306 3680 32312 3732
rect 32364 3680 32370 3732
rect 31220 3624 32168 3652
rect 30852 3556 30972 3584
rect 27341 3519 27399 3525
rect 27341 3485 27353 3519
rect 27387 3485 27399 3519
rect 27341 3479 27399 3485
rect 27430 3476 27436 3528
rect 27488 3476 27494 3528
rect 27614 3476 27620 3528
rect 27672 3476 27678 3528
rect 27706 3476 27712 3528
rect 27764 3476 27770 3528
rect 27893 3519 27951 3525
rect 27893 3485 27905 3519
rect 27939 3485 27951 3519
rect 27893 3479 27951 3485
rect 26531 3451 26589 3457
rect 26531 3417 26543 3451
rect 26577 3448 26589 3451
rect 26697 3451 26755 3457
rect 26577 3420 26648 3448
rect 26577 3417 26589 3420
rect 26531 3411 26589 3417
rect 22186 3380 22192 3392
rect 21376 3352 22192 3380
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 24397 3383 24455 3389
rect 24397 3349 24409 3383
rect 24443 3380 24455 3383
rect 24762 3380 24768 3392
rect 24443 3352 24768 3380
rect 24443 3349 24455 3352
rect 24397 3343 24455 3349
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 26620 3380 26648 3420
rect 26697 3417 26709 3451
rect 26743 3448 26755 3451
rect 27062 3448 27068 3460
rect 26743 3420 27068 3448
rect 26743 3417 26755 3420
rect 26697 3411 26755 3417
rect 27062 3408 27068 3420
rect 27120 3448 27126 3460
rect 27632 3448 27660 3476
rect 27908 3448 27936 3479
rect 28534 3476 28540 3528
rect 28592 3476 28598 3528
rect 28718 3476 28724 3528
rect 28776 3516 28782 3528
rect 28997 3519 29055 3525
rect 28997 3516 29009 3519
rect 28776 3488 29009 3516
rect 28776 3476 28782 3488
rect 28997 3485 29009 3488
rect 29043 3485 29055 3519
rect 28997 3479 29055 3485
rect 27120 3420 27292 3448
rect 27632 3420 27936 3448
rect 28552 3448 28580 3476
rect 28813 3451 28871 3457
rect 28813 3448 28825 3451
rect 28552 3420 28825 3448
rect 27120 3408 27126 3420
rect 26786 3380 26792 3392
rect 26620 3352 26792 3380
rect 26786 3340 26792 3352
rect 26844 3380 26850 3392
rect 27154 3380 27160 3392
rect 26844 3352 27160 3380
rect 26844 3340 26850 3352
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 27264 3380 27292 3420
rect 28813 3417 28825 3420
rect 28859 3417 28871 3451
rect 29012 3448 29040 3479
rect 29730 3476 29736 3528
rect 29788 3476 29794 3528
rect 29825 3519 29883 3525
rect 29825 3485 29837 3519
rect 29871 3516 29883 3519
rect 30653 3519 30711 3525
rect 29871 3488 30236 3516
rect 29871 3485 29883 3488
rect 29825 3479 29883 3485
rect 30009 3451 30067 3457
rect 29012 3420 29776 3448
rect 28813 3411 28871 3417
rect 29178 3380 29184 3392
rect 27264 3352 29184 3380
rect 29178 3340 29184 3352
rect 29236 3340 29242 3392
rect 29748 3380 29776 3420
rect 30009 3417 30021 3451
rect 30055 3417 30067 3451
rect 30009 3411 30067 3417
rect 30024 3380 30052 3411
rect 30098 3408 30104 3460
rect 30156 3448 30162 3460
rect 30208 3448 30236 3488
rect 30653 3485 30665 3519
rect 30699 3485 30711 3519
rect 30653 3479 30711 3485
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3516 30803 3519
rect 30834 3516 30840 3528
rect 30791 3488 30840 3516
rect 30791 3485 30803 3488
rect 30745 3479 30803 3485
rect 30668 3448 30696 3479
rect 30834 3476 30840 3488
rect 30892 3476 30898 3528
rect 30944 3525 30972 3556
rect 30929 3519 30987 3525
rect 30929 3485 30941 3519
rect 30975 3485 30987 3519
rect 30929 3479 30987 3485
rect 31018 3476 31024 3528
rect 31076 3516 31082 3528
rect 31205 3519 31263 3525
rect 31205 3516 31217 3519
rect 31076 3488 31217 3516
rect 31076 3476 31082 3488
rect 31205 3485 31217 3488
rect 31251 3485 31263 3519
rect 31205 3479 31263 3485
rect 31386 3476 31392 3528
rect 31444 3476 31450 3528
rect 31478 3476 31484 3528
rect 31536 3516 31542 3528
rect 31573 3519 31631 3525
rect 31573 3516 31585 3519
rect 31536 3488 31585 3516
rect 31536 3476 31542 3488
rect 31573 3485 31585 3488
rect 31619 3485 31631 3519
rect 31573 3479 31631 3485
rect 31662 3476 31668 3528
rect 31720 3476 31726 3528
rect 32140 3525 32168 3624
rect 31757 3519 31815 3525
rect 31757 3485 31769 3519
rect 31803 3485 31815 3519
rect 31757 3479 31815 3485
rect 32125 3519 32183 3525
rect 32125 3485 32137 3519
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 31294 3448 31300 3460
rect 30156 3420 30236 3448
rect 30484 3420 31300 3448
rect 30156 3408 30162 3420
rect 30484 3389 30512 3420
rect 31294 3408 31300 3420
rect 31352 3408 31358 3460
rect 31772 3448 31800 3479
rect 32306 3476 32312 3528
rect 32364 3476 32370 3528
rect 38470 3476 38476 3528
rect 38528 3476 38534 3528
rect 31404 3420 31800 3448
rect 30301 3383 30359 3389
rect 30301 3380 30313 3383
rect 29748 3352 30313 3380
rect 30301 3349 30313 3352
rect 30347 3349 30359 3383
rect 30301 3343 30359 3349
rect 30469 3383 30527 3389
rect 30469 3349 30481 3383
rect 30515 3349 30527 3383
rect 30469 3343 30527 3349
rect 30742 3340 30748 3392
rect 30800 3380 30806 3392
rect 31404 3380 31432 3420
rect 30800 3352 31432 3380
rect 30800 3340 30806 3352
rect 1104 3290 38824 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 38824 3290
rect 1104 3216 38824 3238
rect 4522 3176 4528 3188
rect 3436 3148 4528 3176
rect 3436 3049 3464 3148
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5626 3136 5632 3188
rect 5684 3136 5690 3188
rect 5994 3136 6000 3188
rect 6052 3136 6058 3188
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 8294 3176 8300 3188
rect 7791 3148 8300 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8864 3148 9352 3176
rect 4154 3108 4160 3120
rect 3896 3080 4160 3108
rect 3896 3049 3924 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4798 3068 4804 3120
rect 4856 3068 4862 3120
rect 7190 3108 7196 3120
rect 6104 3080 7196 3108
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6104 3049 6132 3080
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 8754 3068 8760 3120
rect 8812 3108 8818 3120
rect 8864 3108 8892 3148
rect 8812 3080 8892 3108
rect 8812 3068 8818 3080
rect 9214 3068 9220 3120
rect 9272 3068 9278 3120
rect 9324 3108 9352 3148
rect 13262 3136 13268 3188
rect 13320 3136 13326 3188
rect 24213 3179 24271 3185
rect 22296 3148 23796 3176
rect 9766 3108 9772 3120
rect 9324 3080 9772 3108
rect 9766 3068 9772 3080
rect 9824 3108 9830 3120
rect 9824 3080 9890 3108
rect 9824 3068 9830 3080
rect 11790 3068 11796 3120
rect 11848 3068 11854 3120
rect 12526 3068 12532 3120
rect 12584 3068 12590 3120
rect 22296 3108 22324 3148
rect 23768 3120 23796 3148
rect 24213 3145 24225 3179
rect 24259 3176 24271 3179
rect 25590 3176 25596 3188
rect 24259 3148 25596 3176
rect 24259 3145 24271 3148
rect 24213 3139 24271 3145
rect 25590 3136 25596 3148
rect 25648 3136 25654 3188
rect 26513 3179 26571 3185
rect 26513 3145 26525 3179
rect 26559 3176 26571 3179
rect 26602 3176 26608 3188
rect 26559 3148 26608 3176
rect 26559 3145 26571 3148
rect 26513 3139 26571 3145
rect 26602 3136 26608 3148
rect 26660 3136 26666 3188
rect 27065 3179 27123 3185
rect 27065 3145 27077 3179
rect 27111 3176 27123 3179
rect 27706 3176 27712 3188
rect 27111 3148 27712 3176
rect 27111 3145 27123 3148
rect 27065 3139 27123 3145
rect 27706 3136 27712 3148
rect 27764 3136 27770 3188
rect 30098 3136 30104 3188
rect 30156 3136 30162 3188
rect 31021 3179 31079 3185
rect 31021 3145 31033 3179
rect 31067 3176 31079 3179
rect 31389 3179 31447 3185
rect 31067 3148 31248 3176
rect 31067 3145 31079 3148
rect 31021 3139 31079 3145
rect 22204 3080 22324 3108
rect 22465 3111 22523 3117
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5776 3012 5917 3040
rect 5776 3000 5782 3012
rect 5905 3009 5917 3012
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 7098 3040 7104 3052
rect 6779 3012 7104 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 900 2944 1409 2972
rect 900 2932 906 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2972 3847 2975
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 3835 2944 4169 2972
rect 3835 2941 3847 2944
rect 3789 2935 3847 2941
rect 4157 2941 4169 2944
rect 4203 2941 4215 2975
rect 5920 2972 5948 3003
rect 6564 2972 6592 3003
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 22204 3049 22232 3080
rect 22465 3077 22477 3111
rect 22511 3108 22523 3111
rect 22738 3108 22744 3120
rect 22511 3080 22744 3108
rect 22511 3077 22523 3080
rect 22465 3071 22523 3077
rect 22738 3068 22744 3080
rect 22796 3068 22802 3120
rect 23750 3068 23756 3120
rect 23808 3108 23814 3120
rect 30282 3108 30288 3120
rect 23808 3080 24532 3108
rect 23808 3068 23814 3080
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11379 3012 11529 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 5920 2944 6592 2972
rect 4157 2935 4215 2941
rect 3528 2836 3556 2935
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 8754 2972 8760 2984
rect 7984 2944 8760 2972
rect 7984 2932 7990 2944
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 9493 2975 9551 2981
rect 9493 2941 9505 2975
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6365 2907 6423 2913
rect 6365 2904 6377 2907
rect 5868 2876 6377 2904
rect 5868 2864 5874 2876
rect 6365 2873 6377 2876
rect 6411 2873 6423 2907
rect 6365 2867 6423 2873
rect 3970 2836 3976 2848
rect 3528 2808 3976 2836
rect 3970 2796 3976 2808
rect 4028 2836 4034 2848
rect 5828 2836 5856 2864
rect 4028 2808 5856 2836
rect 4028 2796 4034 2808
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 7156 2808 7205 2836
rect 7156 2796 7162 2808
rect 7193 2805 7205 2808
rect 7239 2805 7251 2839
rect 9508 2836 9536 2935
rect 9582 2932 9588 2984
rect 9640 2932 9646 2984
rect 10502 2932 10508 2984
rect 10560 2972 10566 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 10560 2944 11069 2972
rect 10560 2932 10566 2944
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 11054 2836 11060 2848
rect 9508 2808 11060 2836
rect 7193 2799 7251 2805
rect 11054 2796 11060 2808
rect 11112 2836 11118 2848
rect 11348 2836 11376 3003
rect 23014 2932 23020 2984
rect 23072 2972 23078 2984
rect 23584 2972 23612 3026
rect 24118 3000 24124 3052
rect 24176 3000 24182 3052
rect 24302 3000 24308 3052
rect 24360 3000 24366 3052
rect 24504 3049 24532 3080
rect 24489 3043 24547 3049
rect 24489 3009 24501 3043
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 24762 3000 24768 3052
rect 24820 3040 24826 3052
rect 24857 3043 24915 3049
rect 24857 3040 24869 3043
rect 24820 3012 24869 3040
rect 24820 3000 24826 3012
rect 24857 3009 24869 3012
rect 24903 3009 24915 3043
rect 24857 3003 24915 3009
rect 25608 2972 25636 3094
rect 26436 3080 27016 3108
rect 26436 3049 26464 3080
rect 26421 3043 26479 3049
rect 26421 3009 26433 3043
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 26605 3043 26663 3049
rect 26605 3009 26617 3043
rect 26651 3040 26663 3043
rect 26786 3040 26792 3052
rect 26651 3012 26792 3040
rect 26651 3009 26663 3012
rect 26605 3003 26663 3009
rect 26786 3000 26792 3012
rect 26844 3000 26850 3052
rect 26988 3049 27016 3080
rect 27264 3080 30288 3108
rect 26973 3043 27031 3049
rect 26973 3009 26985 3043
rect 27019 3040 27031 3043
rect 27062 3040 27068 3052
rect 27019 3012 27068 3040
rect 27019 3009 27031 3012
rect 26973 3003 27031 3009
rect 27062 3000 27068 3012
rect 27120 3000 27126 3052
rect 27154 3000 27160 3052
rect 27212 3049 27218 3052
rect 27212 3043 27227 3049
rect 27215 3040 27227 3043
rect 27264 3040 27292 3080
rect 30282 3068 30288 3080
rect 30340 3068 30346 3120
rect 31113 3111 31171 3117
rect 31113 3108 31125 3111
rect 30392 3080 31125 3108
rect 27215 3012 27292 3040
rect 28077 3043 28135 3049
rect 27215 3009 27227 3012
rect 27212 3003 27227 3009
rect 28077 3009 28089 3043
rect 28123 3040 28135 3043
rect 30009 3043 30067 3049
rect 30009 3040 30021 3043
rect 28123 3012 30021 3040
rect 28123 3009 28135 3012
rect 28077 3003 28135 3009
rect 30009 3009 30021 3012
rect 30055 3009 30067 3043
rect 30009 3003 30067 3009
rect 27212 3000 27218 3003
rect 28092 2972 28120 3003
rect 23072 2944 25636 2972
rect 26160 2944 28120 2972
rect 23072 2932 23078 2944
rect 11112 2808 11376 2836
rect 23937 2839 23995 2845
rect 11112 2796 11118 2808
rect 23937 2805 23949 2839
rect 23983 2836 23995 2839
rect 24394 2836 24400 2848
rect 23983 2808 24400 2836
rect 23983 2805 23995 2808
rect 23937 2799 23995 2805
rect 24394 2796 24400 2808
rect 24452 2836 24458 2848
rect 26160 2836 26188 2944
rect 28166 2932 28172 2984
rect 28224 2932 28230 2984
rect 28445 2975 28503 2981
rect 28445 2941 28457 2975
rect 28491 2972 28503 2975
rect 28534 2972 28540 2984
rect 28491 2944 28540 2972
rect 28491 2941 28503 2944
rect 28445 2935 28503 2941
rect 28534 2932 28540 2944
rect 28592 2932 28598 2984
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 30392 2972 30420 3080
rect 31113 3077 31125 3080
rect 31159 3077 31171 3111
rect 31220 3108 31248 3148
rect 31389 3145 31401 3179
rect 31435 3176 31447 3179
rect 32306 3176 32312 3188
rect 31435 3148 32312 3176
rect 31435 3145 31447 3148
rect 31389 3139 31447 3145
rect 32306 3136 32312 3148
rect 32364 3136 32370 3188
rect 31570 3108 31576 3120
rect 31220 3080 31576 3108
rect 31113 3071 31171 3077
rect 31570 3068 31576 3080
rect 31628 3068 31634 3120
rect 30742 3000 30748 3052
rect 30800 3000 30806 3052
rect 30837 3043 30895 3049
rect 30837 3009 30849 3043
rect 30883 3040 30895 3043
rect 30926 3040 30932 3052
rect 30883 3012 30932 3040
rect 30883 3009 30895 3012
rect 30837 3003 30895 3009
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 31294 3000 31300 3052
rect 31352 3000 31358 3052
rect 31389 3043 31447 3049
rect 31389 3009 31401 3043
rect 31435 3040 31447 3043
rect 31478 3040 31484 3052
rect 31435 3012 31484 3040
rect 31435 3009 31447 3012
rect 31389 3003 31447 3009
rect 31478 3000 31484 3012
rect 31536 3000 31542 3052
rect 29144 2944 30420 2972
rect 29144 2932 29150 2944
rect 30558 2932 30564 2984
rect 30616 2972 30622 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30616 2944 31033 2972
rect 30616 2932 30622 2944
rect 31021 2941 31033 2944
rect 31067 2972 31079 2975
rect 31662 2972 31668 2984
rect 31067 2944 31668 2972
rect 31067 2941 31079 2944
rect 31021 2935 31079 2941
rect 31662 2932 31668 2944
rect 31720 2932 31726 2984
rect 38470 2932 38476 2984
rect 38528 2932 38534 2984
rect 26283 2907 26341 2913
rect 26283 2873 26295 2907
rect 26329 2904 26341 2907
rect 26970 2904 26976 2916
rect 26329 2876 26976 2904
rect 26329 2873 26341 2876
rect 26283 2867 26341 2873
rect 26970 2864 26976 2876
rect 27028 2904 27034 2916
rect 31386 2904 31392 2916
rect 27028 2876 31392 2904
rect 27028 2864 27034 2876
rect 31386 2864 31392 2876
rect 31444 2864 31450 2916
rect 24452 2808 26188 2836
rect 24452 2796 24458 2808
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 34790 2836 34796 2848
rect 30340 2808 34796 2836
rect 30340 2796 30346 2808
rect 34790 2796 34796 2808
rect 34848 2796 34854 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8628 2604 8953 2632
rect 8628 2592 8634 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 14918 2592 14924 2644
rect 14976 2632 14982 2644
rect 15105 2635 15163 2641
rect 15105 2632 15117 2635
rect 14976 2604 15117 2632
rect 14976 2592 14982 2604
rect 15105 2601 15117 2604
rect 15151 2601 15163 2635
rect 15105 2595 15163 2601
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 5500 2468 6929 2496
rect 5500 2456 5506 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7282 2496 7288 2508
rect 7239 2468 7288 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8536 2468 8677 2496
rect 8536 2456 8542 2468
rect 8665 2465 8677 2468
rect 8711 2496 8723 2499
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 8711 2468 9505 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14844 2400 14933 2428
rect 7926 2320 7932 2372
rect 7984 2320 7990 2372
rect 14844 2304 14872 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 21358 2388 21364 2440
rect 21416 2388 21422 2440
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 23937 2431 23995 2437
rect 23937 2428 23949 2431
rect 23900 2400 23949 2428
rect 23900 2388 23906 2400
rect 23937 2397 23949 2400
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30377 2431 30435 2437
rect 30377 2428 30389 2431
rect 30340 2400 30389 2428
rect 30340 2388 30346 2400
rect 30377 2397 30389 2400
rect 30423 2397 30435 2431
rect 30377 2391 30435 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35492 2400 35541 2428
rect 35492 2388 35498 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 36136 2400 36185 2428
rect 36136 2388 36142 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 36173 2391 36231 2397
rect 14826 2252 14832 2304
rect 14884 2252 14890 2304
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 21324 2264 21557 2292
rect 21324 2252 21330 2264
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24544 2264 24593 2292
rect 24544 2252 24550 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 27062 2252 27068 2304
rect 27120 2292 27126 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 27120 2264 27169 2292
rect 27120 2252 27126 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27801 2295 27859 2301
rect 27801 2292 27813 2295
rect 27764 2264 27813 2292
rect 27764 2252 27770 2264
rect 27801 2261 27813 2264
rect 27847 2261 27859 2295
rect 27801 2255 27859 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29089 2295 29147 2301
rect 29089 2292 29101 2295
rect 29052 2264 29101 2292
rect 29052 2252 29058 2264
rect 29089 2261 29101 2264
rect 29135 2261 29147 2295
rect 29089 2255 29147 2261
rect 38470 2252 38476 2304
rect 38528 2252 38534 2304
rect 1104 2202 38824 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1308 37408 1360 37460
rect 3240 37408 3292 37460
rect 27712 37408 27764 37460
rect 29000 37408 29052 37460
rect 29644 37408 29696 37460
rect 34152 37408 34204 37460
rect 34796 37408 34848 37460
rect 35440 37408 35492 37460
rect 36084 37408 36136 37460
rect 36728 37408 36780 37460
rect 37924 37451 37976 37460
rect 37924 37417 37933 37451
rect 37933 37417 37967 37451
rect 37967 37417 37976 37451
rect 37924 37408 37976 37417
rect 38200 37451 38252 37460
rect 38200 37417 38209 37451
rect 38209 37417 38243 37451
rect 38243 37417 38252 37451
rect 38200 37408 38252 37417
rect 848 37272 900 37324
rect 5172 37204 5224 37256
rect 8116 37204 8168 37256
rect 24216 37247 24268 37256
rect 24216 37213 24225 37247
rect 24225 37213 24259 37247
rect 24259 37213 24268 37247
rect 24216 37204 24268 37213
rect 25504 37247 25556 37256
rect 25504 37213 25513 37247
rect 25513 37213 25547 37247
rect 25547 37213 25556 37247
rect 25504 37204 25556 37213
rect 20812 37179 20864 37188
rect 20812 37145 20821 37179
rect 20821 37145 20855 37179
rect 20855 37145 20864 37179
rect 20812 37136 20864 37145
rect 21180 37136 21232 37188
rect 6828 37068 6880 37120
rect 19616 37068 19668 37120
rect 23848 37068 23900 37120
rect 26976 37204 27028 37256
rect 27068 37204 27120 37256
rect 28356 37204 28408 37256
rect 30288 37204 30340 37256
rect 30932 37204 30984 37256
rect 31576 37204 31628 37256
rect 32220 37204 32272 37256
rect 32864 37204 32916 37256
rect 33508 37204 33560 37256
rect 25780 37068 25832 37120
rect 26424 37068 26476 37120
rect 38476 37111 38528 37120
rect 38476 37077 38485 37111
rect 38485 37077 38519 37111
rect 38519 37077 38528 37111
rect 38476 37068 38528 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 5724 36796 5776 36848
rect 19432 36839 19484 36848
rect 19432 36805 19441 36839
rect 19441 36805 19475 36839
rect 19475 36805 19484 36839
rect 19432 36796 19484 36805
rect 20076 36796 20128 36848
rect 20812 36864 20864 36916
rect 21732 36864 21784 36916
rect 24216 36907 24268 36916
rect 24216 36873 24225 36907
rect 24225 36873 24259 36907
rect 24259 36873 24268 36907
rect 24216 36864 24268 36873
rect 26976 36907 27028 36916
rect 26976 36873 26985 36907
rect 26985 36873 27019 36907
rect 27019 36873 27028 36907
rect 26976 36864 27028 36873
rect 30104 36864 30156 36916
rect 23940 36796 23992 36848
rect 27988 36796 28040 36848
rect 31852 36796 31904 36848
rect 8208 36728 8260 36780
rect 8392 36728 8444 36780
rect 5172 36660 5224 36712
rect 6552 36660 6604 36712
rect 7196 36660 7248 36712
rect 8944 36771 8996 36780
rect 8944 36737 8953 36771
rect 8953 36737 8987 36771
rect 8987 36737 8996 36771
rect 8944 36728 8996 36737
rect 19248 36660 19300 36712
rect 24400 36771 24452 36780
rect 24400 36737 24409 36771
rect 24409 36737 24443 36771
rect 24443 36737 24452 36771
rect 24400 36728 24452 36737
rect 27160 36771 27212 36780
rect 27160 36737 27169 36771
rect 27169 36737 27203 36771
rect 27203 36737 27212 36771
rect 27160 36728 27212 36737
rect 38292 36728 38344 36780
rect 38568 36728 38620 36780
rect 21364 36660 21416 36712
rect 6184 36567 6236 36576
rect 6184 36533 6193 36567
rect 6193 36533 6227 36567
rect 6227 36533 6236 36567
rect 6184 36524 6236 36533
rect 7288 36524 7340 36576
rect 8116 36524 8168 36576
rect 8668 36524 8720 36576
rect 19616 36567 19668 36576
rect 19616 36533 19625 36567
rect 19625 36533 19659 36567
rect 19659 36533 19668 36567
rect 19616 36524 19668 36533
rect 22652 36703 22704 36712
rect 22652 36669 22661 36703
rect 22661 36669 22695 36703
rect 22695 36669 22704 36703
rect 22652 36660 22704 36669
rect 24860 36703 24912 36712
rect 24860 36669 24869 36703
rect 24869 36669 24903 36703
rect 24903 36669 24912 36703
rect 24860 36660 24912 36669
rect 25136 36703 25188 36712
rect 25136 36669 25145 36703
rect 25145 36669 25179 36703
rect 25179 36669 25188 36703
rect 25136 36660 25188 36669
rect 27528 36660 27580 36712
rect 28356 36660 28408 36712
rect 29368 36660 29420 36712
rect 33140 36660 33192 36712
rect 24124 36567 24176 36576
rect 24124 36533 24133 36567
rect 24133 36533 24167 36567
rect 24167 36533 24176 36567
rect 24124 36524 24176 36533
rect 26608 36567 26660 36576
rect 26608 36533 26617 36567
rect 26617 36533 26651 36567
rect 26651 36533 26660 36567
rect 26608 36524 26660 36533
rect 29460 36567 29512 36576
rect 29460 36533 29469 36567
rect 29469 36533 29503 36567
rect 29503 36533 29512 36567
rect 29460 36524 29512 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 848 36252 900 36304
rect 3332 36184 3384 36236
rect 4436 36159 4488 36168
rect 4436 36125 4445 36159
rect 4445 36125 4479 36159
rect 4479 36125 4488 36159
rect 4436 36116 4488 36125
rect 5172 36363 5224 36372
rect 5172 36329 5181 36363
rect 5181 36329 5215 36363
rect 5215 36329 5224 36363
rect 5172 36320 5224 36329
rect 7196 36363 7248 36372
rect 7196 36329 7205 36363
rect 7205 36329 7239 36363
rect 7239 36329 7248 36363
rect 7196 36320 7248 36329
rect 7472 36363 7524 36372
rect 7472 36329 7481 36363
rect 7481 36329 7515 36363
rect 7515 36329 7524 36363
rect 7472 36320 7524 36329
rect 8116 36320 8168 36372
rect 8944 36363 8996 36372
rect 8944 36329 8953 36363
rect 8953 36329 8987 36363
rect 8987 36329 8996 36363
rect 8944 36320 8996 36329
rect 20076 36320 20128 36372
rect 5264 36252 5316 36304
rect 5632 36159 5684 36168
rect 5632 36125 5641 36159
rect 5641 36125 5675 36159
rect 5675 36125 5684 36159
rect 5632 36116 5684 36125
rect 6184 36116 6236 36168
rect 6644 36116 6696 36168
rect 6828 36159 6880 36168
rect 6828 36125 6837 36159
rect 6837 36125 6871 36159
rect 6871 36125 6880 36159
rect 6828 36116 6880 36125
rect 4712 35980 4764 36032
rect 5540 36048 5592 36100
rect 7196 36048 7248 36100
rect 8392 36184 8444 36236
rect 8668 36227 8720 36236
rect 8668 36193 8677 36227
rect 8677 36193 8711 36227
rect 8711 36193 8720 36227
rect 8668 36184 8720 36193
rect 8116 36116 8168 36168
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 20812 36116 20864 36168
rect 21272 36159 21324 36168
rect 21272 36125 21281 36159
rect 21281 36125 21315 36159
rect 21315 36125 21324 36159
rect 21272 36116 21324 36125
rect 21732 36363 21784 36372
rect 21732 36329 21741 36363
rect 21741 36329 21775 36363
rect 21775 36329 21784 36363
rect 21732 36320 21784 36329
rect 22652 36320 22704 36372
rect 24400 36363 24452 36372
rect 24400 36329 24409 36363
rect 24409 36329 24443 36363
rect 24443 36329 24452 36363
rect 24400 36320 24452 36329
rect 25136 36320 25188 36372
rect 27160 36320 27212 36372
rect 28356 36363 28408 36372
rect 28356 36329 28365 36363
rect 28365 36329 28399 36363
rect 28399 36329 28408 36363
rect 28356 36320 28408 36329
rect 29276 36320 29328 36372
rect 29368 36363 29420 36372
rect 29368 36329 29377 36363
rect 29377 36329 29411 36363
rect 29411 36329 29420 36363
rect 29368 36320 29420 36329
rect 19524 36091 19576 36100
rect 19524 36057 19533 36091
rect 19533 36057 19567 36091
rect 19567 36057 19576 36091
rect 19524 36048 19576 36057
rect 19984 36048 20036 36100
rect 22192 36116 22244 36168
rect 23664 36184 23716 36236
rect 22376 36116 22428 36168
rect 23756 36116 23808 36168
rect 24768 36184 24820 36236
rect 27620 36252 27672 36304
rect 25044 36184 25096 36236
rect 24124 36116 24176 36168
rect 24216 36116 24268 36168
rect 26608 36184 26660 36236
rect 26148 36159 26200 36168
rect 26148 36125 26160 36159
rect 26160 36125 26194 36159
rect 26194 36125 26200 36159
rect 26148 36116 26200 36125
rect 26976 36048 27028 36100
rect 7748 35980 7800 36032
rect 7840 36023 7892 36032
rect 7840 35989 7849 36023
rect 7849 35989 7883 36023
rect 7883 35989 7892 36023
rect 7840 35980 7892 35989
rect 20996 36023 21048 36032
rect 20996 35989 21005 36023
rect 21005 35989 21039 36023
rect 21039 35989 21048 36023
rect 20996 35980 21048 35989
rect 21456 36023 21508 36032
rect 21456 35989 21465 36023
rect 21465 35989 21499 36023
rect 21499 35989 21508 36023
rect 21456 35980 21508 35989
rect 22284 35980 22336 36032
rect 25228 36023 25280 36032
rect 25228 35989 25237 36023
rect 25237 35989 25271 36023
rect 25271 35989 25280 36023
rect 25228 35980 25280 35989
rect 27344 35980 27396 36032
rect 27620 36091 27672 36100
rect 27620 36057 27629 36091
rect 27629 36057 27663 36091
rect 27663 36057 27672 36091
rect 27620 36048 27672 36057
rect 27804 36091 27856 36100
rect 27804 36057 27813 36091
rect 27813 36057 27847 36091
rect 27847 36057 27856 36091
rect 27804 36048 27856 36057
rect 28172 36048 28224 36100
rect 29460 36116 29512 36168
rect 30104 36159 30156 36168
rect 30104 36125 30113 36159
rect 30113 36125 30147 36159
rect 30147 36125 30156 36159
rect 30104 36116 30156 36125
rect 31852 36116 31904 36168
rect 28816 35980 28868 36032
rect 29000 36091 29052 36100
rect 29000 36057 29009 36091
rect 29009 36057 29043 36091
rect 29043 36057 29052 36091
rect 29000 36048 29052 36057
rect 30748 36091 30800 36100
rect 30748 36057 30757 36091
rect 30757 36057 30791 36091
rect 30791 36057 30800 36091
rect 30748 36048 30800 36057
rect 38476 36091 38528 36100
rect 38476 36057 38485 36091
rect 38485 36057 38519 36091
rect 38519 36057 38528 36091
rect 38476 36048 38528 36057
rect 29184 36023 29236 36032
rect 29184 35989 29209 36023
rect 29209 35989 29236 36023
rect 29184 35980 29236 35989
rect 32220 36023 32272 36032
rect 32220 35989 32229 36023
rect 32229 35989 32263 36023
rect 32263 35989 32272 36023
rect 32220 35980 32272 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 4436 35776 4488 35828
rect 5448 35776 5500 35828
rect 5540 35819 5592 35828
rect 5540 35785 5549 35819
rect 5549 35785 5583 35819
rect 5583 35785 5592 35819
rect 5540 35776 5592 35785
rect 7288 35708 7340 35760
rect 5264 35683 5316 35692
rect 5264 35649 5273 35683
rect 5273 35649 5307 35683
rect 5307 35649 5316 35683
rect 5264 35640 5316 35649
rect 6552 35683 6604 35692
rect 6552 35649 6561 35683
rect 6561 35649 6595 35683
rect 6595 35649 6604 35683
rect 6552 35640 6604 35649
rect 8116 35776 8168 35828
rect 19524 35776 19576 35828
rect 23756 35819 23808 35828
rect 23756 35785 23765 35819
rect 23765 35785 23799 35819
rect 23799 35785 23808 35819
rect 23756 35776 23808 35785
rect 21824 35708 21876 35760
rect 8760 35640 8812 35692
rect 13084 35683 13136 35692
rect 13084 35649 13093 35683
rect 13093 35649 13127 35683
rect 13127 35649 13136 35683
rect 13084 35640 13136 35649
rect 19432 35640 19484 35692
rect 848 35572 900 35624
rect 4712 35572 4764 35624
rect 6092 35615 6144 35624
rect 6092 35581 6101 35615
rect 6101 35581 6135 35615
rect 6135 35581 6144 35615
rect 6092 35572 6144 35581
rect 7840 35572 7892 35624
rect 8024 35572 8076 35624
rect 11060 35572 11112 35624
rect 13636 35572 13688 35624
rect 10876 35504 10928 35556
rect 20076 35640 20128 35692
rect 21456 35640 21508 35692
rect 23664 35683 23716 35692
rect 23664 35649 23673 35683
rect 23673 35649 23707 35683
rect 23707 35649 23716 35683
rect 23664 35640 23716 35649
rect 23848 35683 23900 35692
rect 23848 35649 23857 35683
rect 23857 35649 23891 35683
rect 23891 35649 23900 35683
rect 24032 35751 24084 35760
rect 24032 35717 24041 35751
rect 24041 35717 24075 35751
rect 24075 35717 24084 35751
rect 24032 35708 24084 35717
rect 24768 35776 24820 35828
rect 23848 35640 23900 35649
rect 25228 35776 25280 35828
rect 29184 35776 29236 35828
rect 30748 35776 30800 35828
rect 20996 35572 21048 35624
rect 20444 35504 20496 35556
rect 3240 35436 3292 35488
rect 4620 35479 4672 35488
rect 4620 35445 4629 35479
rect 4629 35445 4663 35479
rect 4663 35445 4672 35479
rect 4620 35436 4672 35445
rect 8392 35479 8444 35488
rect 8392 35445 8401 35479
rect 8401 35445 8435 35479
rect 8435 35445 8444 35479
rect 8392 35436 8444 35445
rect 12440 35436 12492 35488
rect 20536 35479 20588 35488
rect 20536 35445 20545 35479
rect 20545 35445 20579 35479
rect 20579 35445 20588 35479
rect 20536 35436 20588 35445
rect 21272 35504 21324 35556
rect 21916 35504 21968 35556
rect 24768 35683 24820 35692
rect 24768 35649 24777 35683
rect 24777 35649 24811 35683
rect 24811 35649 24820 35683
rect 24768 35640 24820 35649
rect 25136 35683 25188 35692
rect 25136 35649 25145 35683
rect 25145 35649 25179 35683
rect 25179 35649 25188 35683
rect 25136 35640 25188 35649
rect 26148 35640 26200 35692
rect 26240 35504 26292 35556
rect 26608 35640 26660 35692
rect 27528 35708 27580 35760
rect 27988 35708 28040 35760
rect 29460 35708 29512 35760
rect 27620 35572 27672 35624
rect 30472 35708 30524 35760
rect 30104 35640 30156 35692
rect 30196 35504 30248 35556
rect 30840 35615 30892 35624
rect 30840 35581 30849 35615
rect 30849 35581 30883 35615
rect 30883 35581 30892 35615
rect 30840 35572 30892 35581
rect 31760 35572 31812 35624
rect 32220 35572 32272 35624
rect 22284 35436 22336 35488
rect 24216 35479 24268 35488
rect 24216 35445 24225 35479
rect 24225 35445 24259 35479
rect 24259 35445 24268 35479
rect 24216 35436 24268 35445
rect 24308 35436 24360 35488
rect 25136 35436 25188 35488
rect 27068 35436 27120 35488
rect 27436 35436 27488 35488
rect 29000 35436 29052 35488
rect 30472 35436 30524 35488
rect 32036 35436 32088 35488
rect 38476 35479 38528 35488
rect 38476 35445 38485 35479
rect 38485 35445 38519 35479
rect 38519 35445 38528 35479
rect 38476 35436 38528 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3976 35232 4028 35284
rect 5724 35232 5776 35284
rect 6092 35275 6144 35284
rect 6092 35241 6101 35275
rect 6101 35241 6135 35275
rect 6135 35241 6144 35275
rect 6092 35232 6144 35241
rect 7472 35232 7524 35284
rect 8024 35275 8076 35284
rect 8024 35241 8033 35275
rect 8033 35241 8067 35275
rect 8067 35241 8076 35275
rect 8024 35232 8076 35241
rect 10784 35232 10836 35284
rect 2872 35139 2924 35148
rect 2872 35105 2881 35139
rect 2881 35105 2915 35139
rect 2915 35105 2924 35139
rect 2872 35096 2924 35105
rect 3332 35139 3384 35148
rect 3332 35105 3341 35139
rect 3341 35105 3375 35139
rect 3375 35105 3384 35139
rect 3332 35096 3384 35105
rect 848 35028 900 35080
rect 3240 35071 3292 35080
rect 3240 35037 3249 35071
rect 3249 35037 3283 35071
rect 3283 35037 3292 35071
rect 3240 35028 3292 35037
rect 4620 35096 4672 35148
rect 8392 35164 8444 35216
rect 12716 35232 12768 35284
rect 13084 35232 13136 35284
rect 17040 35232 17092 35284
rect 20536 35232 20588 35284
rect 22192 35275 22244 35284
rect 22192 35241 22201 35275
rect 22201 35241 22235 35275
rect 22235 35241 22244 35275
rect 22192 35232 22244 35241
rect 24308 35232 24360 35284
rect 7748 35139 7800 35148
rect 7748 35105 7757 35139
rect 7757 35105 7791 35139
rect 7791 35105 7800 35139
rect 7748 35096 7800 35105
rect 11060 35096 11112 35148
rect 4344 35071 4396 35080
rect 4344 35037 4353 35071
rect 4353 35037 4387 35071
rect 4387 35037 4396 35071
rect 4344 35028 4396 35037
rect 5724 35028 5776 35080
rect 6644 35028 6696 35080
rect 7196 35071 7248 35080
rect 7196 35037 7205 35071
rect 7205 35037 7239 35071
rect 7239 35037 7248 35071
rect 7196 35028 7248 35037
rect 13544 35096 13596 35148
rect 12716 35028 12768 35080
rect 13452 35071 13504 35080
rect 13452 35037 13461 35071
rect 13461 35037 13495 35071
rect 13495 35037 13504 35071
rect 13452 35028 13504 35037
rect 13912 35028 13964 35080
rect 16304 35164 16356 35216
rect 24032 35207 24084 35216
rect 24032 35173 24041 35207
rect 24041 35173 24075 35207
rect 24075 35173 24084 35207
rect 24032 35164 24084 35173
rect 10968 34960 11020 35012
rect 15016 34960 15068 35012
rect 22192 35096 22244 35148
rect 24216 35096 24268 35148
rect 24952 35139 25004 35148
rect 24952 35105 24961 35139
rect 24961 35105 24995 35139
rect 24995 35105 25004 35139
rect 24952 35096 25004 35105
rect 15660 35071 15712 35080
rect 15660 35037 15669 35071
rect 15669 35037 15703 35071
rect 15703 35037 15712 35071
rect 15660 35028 15712 35037
rect 17500 35028 17552 35080
rect 18328 35071 18380 35080
rect 18328 35037 18337 35071
rect 18337 35037 18371 35071
rect 18371 35037 18380 35071
rect 18328 35028 18380 35037
rect 22376 35028 22428 35080
rect 23296 35028 23348 35080
rect 23664 35028 23716 35080
rect 15292 34960 15344 35012
rect 16120 34960 16172 35012
rect 17408 34960 17460 35012
rect 21364 34960 21416 35012
rect 23848 35028 23900 35080
rect 27252 35275 27304 35284
rect 27252 35241 27261 35275
rect 27261 35241 27295 35275
rect 27295 35241 27304 35275
rect 27252 35232 27304 35241
rect 27436 35275 27488 35284
rect 27436 35241 27445 35275
rect 27445 35241 27479 35275
rect 27479 35241 27488 35275
rect 27436 35232 27488 35241
rect 30840 35232 30892 35284
rect 31208 35232 31260 35284
rect 32404 35232 32456 35284
rect 26148 35164 26200 35216
rect 30196 35164 30248 35216
rect 26240 35096 26292 35148
rect 27160 35028 27212 35080
rect 26976 34960 27028 35012
rect 27344 34960 27396 35012
rect 27620 35028 27672 35080
rect 27804 35096 27856 35148
rect 30104 35096 30156 35148
rect 32128 35164 32180 35216
rect 29276 35028 29328 35080
rect 29736 35071 29788 35080
rect 29736 35037 29745 35071
rect 29745 35037 29779 35071
rect 29779 35037 29788 35071
rect 29736 35028 29788 35037
rect 30196 35071 30248 35080
rect 30196 35037 30205 35071
rect 30205 35037 30239 35071
rect 30239 35037 30248 35071
rect 30196 35028 30248 35037
rect 28172 34960 28224 35012
rect 28724 34960 28776 35012
rect 29920 34960 29972 35012
rect 30656 35028 30708 35080
rect 32036 35096 32088 35148
rect 33324 35096 33376 35148
rect 31208 35071 31260 35080
rect 31208 35037 31217 35071
rect 31217 35037 31251 35071
rect 31251 35037 31260 35071
rect 31208 35028 31260 35037
rect 31852 35028 31904 35080
rect 5264 34892 5316 34944
rect 7380 34935 7432 34944
rect 7380 34901 7389 34935
rect 7389 34901 7423 34935
rect 7423 34901 7432 34935
rect 7380 34892 7432 34901
rect 11704 34892 11756 34944
rect 13084 34892 13136 34944
rect 15476 34892 15528 34944
rect 16028 34892 16080 34944
rect 17500 34892 17552 34944
rect 17868 34892 17920 34944
rect 18880 34892 18932 34944
rect 22928 34935 22980 34944
rect 22928 34901 22937 34935
rect 22937 34901 22971 34935
rect 22971 34901 22980 34935
rect 22928 34892 22980 34901
rect 24584 34892 24636 34944
rect 25228 34892 25280 34944
rect 27436 34892 27488 34944
rect 30380 34935 30432 34944
rect 30380 34901 30389 34935
rect 30389 34901 30423 34935
rect 30423 34901 30432 34935
rect 30380 34892 30432 34901
rect 31024 34892 31076 34944
rect 31760 34960 31812 35012
rect 31668 34892 31720 34944
rect 31944 34892 31996 34944
rect 38476 34935 38528 34944
rect 38476 34901 38485 34935
rect 38485 34901 38519 34935
rect 38519 34901 38528 34935
rect 38476 34892 38528 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 2228 34484 2280 34536
rect 3884 34688 3936 34740
rect 10968 34731 11020 34740
rect 10968 34697 10977 34731
rect 10977 34697 11011 34731
rect 11011 34697 11020 34731
rect 10968 34688 11020 34697
rect 2872 34663 2924 34672
rect 2872 34629 2881 34663
rect 2881 34629 2915 34663
rect 2915 34629 2924 34663
rect 2872 34620 2924 34629
rect 4344 34620 4396 34672
rect 3976 34552 4028 34604
rect 6552 34552 6604 34604
rect 9772 34595 9824 34604
rect 9772 34561 9781 34595
rect 9781 34561 9815 34595
rect 9815 34561 9824 34595
rect 9772 34552 9824 34561
rect 6368 34484 6420 34536
rect 9220 34484 9272 34536
rect 9956 34527 10008 34536
rect 9956 34493 9965 34527
rect 9965 34493 9999 34527
rect 9999 34493 10008 34527
rect 10784 34595 10836 34604
rect 10784 34561 10793 34595
rect 10793 34561 10827 34595
rect 10827 34561 10836 34595
rect 10784 34552 10836 34561
rect 10876 34595 10928 34604
rect 10876 34561 10885 34595
rect 10885 34561 10919 34595
rect 10919 34561 10928 34595
rect 10876 34552 10928 34561
rect 11704 34620 11756 34672
rect 9956 34484 10008 34493
rect 12624 34688 12676 34740
rect 13912 34731 13964 34740
rect 13912 34697 13921 34731
rect 13921 34697 13955 34731
rect 13955 34697 13964 34731
rect 13912 34688 13964 34697
rect 12440 34663 12492 34672
rect 12440 34629 12449 34663
rect 12449 34629 12483 34663
rect 12483 34629 12492 34663
rect 12440 34620 12492 34629
rect 13728 34620 13780 34672
rect 14924 34620 14976 34672
rect 15476 34663 15528 34672
rect 15476 34629 15485 34663
rect 15485 34629 15519 34663
rect 15519 34629 15528 34663
rect 15476 34620 15528 34629
rect 15660 34688 15712 34740
rect 17408 34731 17460 34740
rect 17408 34697 17417 34731
rect 17417 34697 17451 34731
rect 17451 34697 17460 34731
rect 17408 34688 17460 34697
rect 17592 34688 17644 34740
rect 13544 34552 13596 34604
rect 14464 34552 14516 34604
rect 16120 34620 16172 34672
rect 19984 34688 20036 34740
rect 21732 34688 21784 34740
rect 21824 34731 21876 34740
rect 21824 34697 21833 34731
rect 21833 34697 21867 34731
rect 21867 34697 21876 34731
rect 21824 34688 21876 34697
rect 21916 34688 21968 34740
rect 22928 34688 22980 34740
rect 29736 34688 29788 34740
rect 16028 34595 16080 34604
rect 16028 34561 16037 34595
rect 16037 34561 16071 34595
rect 16071 34561 16080 34595
rect 16028 34552 16080 34561
rect 16304 34595 16356 34604
rect 16304 34561 16313 34595
rect 16313 34561 16347 34595
rect 16347 34561 16356 34595
rect 16304 34552 16356 34561
rect 12164 34527 12216 34536
rect 12164 34493 12173 34527
rect 12173 34493 12207 34527
rect 12207 34493 12216 34527
rect 12164 34484 12216 34493
rect 13084 34484 13136 34536
rect 15016 34484 15068 34536
rect 15752 34527 15804 34536
rect 15752 34493 15761 34527
rect 15761 34493 15795 34527
rect 15795 34493 15804 34527
rect 15752 34484 15804 34493
rect 17040 34595 17092 34604
rect 17040 34561 17049 34595
rect 17049 34561 17083 34595
rect 17083 34561 17092 34595
rect 17040 34552 17092 34561
rect 18880 34663 18932 34672
rect 18880 34629 18889 34663
rect 18889 34629 18923 34663
rect 18923 34629 18932 34663
rect 18880 34620 18932 34629
rect 23940 34620 23992 34672
rect 24584 34663 24636 34672
rect 24584 34629 24593 34663
rect 24593 34629 24627 34663
rect 24627 34629 24636 34663
rect 24584 34620 24636 34629
rect 24952 34620 25004 34672
rect 17868 34484 17920 34536
rect 19248 34484 19300 34536
rect 20352 34527 20404 34536
rect 20352 34493 20361 34527
rect 20361 34493 20395 34527
rect 20395 34493 20404 34527
rect 20352 34484 20404 34493
rect 4712 34348 4764 34400
rect 5080 34348 5132 34400
rect 5632 34348 5684 34400
rect 10232 34391 10284 34400
rect 10232 34357 10241 34391
rect 10241 34357 10275 34391
rect 10275 34357 10284 34391
rect 10232 34348 10284 34357
rect 10324 34391 10376 34400
rect 10324 34357 10333 34391
rect 10333 34357 10367 34391
rect 10367 34357 10376 34391
rect 10324 34348 10376 34357
rect 11612 34348 11664 34400
rect 16212 34348 16264 34400
rect 20352 34348 20404 34400
rect 21824 34416 21876 34468
rect 22100 34527 22152 34536
rect 22100 34493 22109 34527
rect 22109 34493 22143 34527
rect 22143 34493 22152 34527
rect 22100 34484 22152 34493
rect 22284 34595 22336 34604
rect 22284 34561 22293 34595
rect 22293 34561 22327 34595
rect 22327 34561 22336 34595
rect 22284 34552 22336 34561
rect 22468 34484 22520 34536
rect 22836 34595 22888 34604
rect 22836 34561 22845 34595
rect 22845 34561 22879 34595
rect 22879 34561 22888 34595
rect 22836 34552 22888 34561
rect 24860 34595 24912 34604
rect 24860 34561 24869 34595
rect 24869 34561 24903 34595
rect 24903 34561 24912 34595
rect 24860 34552 24912 34561
rect 25228 34595 25280 34604
rect 25228 34561 25237 34595
rect 25237 34561 25271 34595
rect 25271 34561 25280 34595
rect 25228 34552 25280 34561
rect 26148 34595 26200 34604
rect 26148 34561 26157 34595
rect 26157 34561 26191 34595
rect 26191 34561 26200 34595
rect 26148 34552 26200 34561
rect 28724 34595 28776 34604
rect 28724 34561 28733 34595
rect 28733 34561 28767 34595
rect 28767 34561 28776 34595
rect 28724 34552 28776 34561
rect 23848 34484 23900 34536
rect 25136 34527 25188 34536
rect 25136 34493 25145 34527
rect 25145 34493 25179 34527
rect 25179 34493 25188 34527
rect 25136 34484 25188 34493
rect 28448 34527 28500 34536
rect 28448 34493 28457 34527
rect 28457 34493 28491 34527
rect 28491 34493 28500 34527
rect 28448 34484 28500 34493
rect 28632 34527 28684 34536
rect 28632 34493 28641 34527
rect 28641 34493 28675 34527
rect 28675 34493 28684 34527
rect 28632 34484 28684 34493
rect 23020 34459 23072 34468
rect 23020 34425 23029 34459
rect 23029 34425 23063 34459
rect 23063 34425 23072 34459
rect 23020 34416 23072 34425
rect 27896 34416 27948 34468
rect 29184 34552 29236 34604
rect 29276 34552 29328 34604
rect 30196 34620 30248 34672
rect 29000 34484 29052 34536
rect 22100 34348 22152 34400
rect 22836 34348 22888 34400
rect 29000 34391 29052 34400
rect 29000 34357 29009 34391
rect 29009 34357 29043 34391
rect 29043 34357 29052 34391
rect 29000 34348 29052 34357
rect 30104 34595 30156 34604
rect 30104 34561 30113 34595
rect 30113 34561 30147 34595
rect 30147 34561 30156 34595
rect 30104 34552 30156 34561
rect 30288 34595 30340 34604
rect 30288 34561 30297 34595
rect 30297 34561 30331 34595
rect 30331 34561 30340 34595
rect 30288 34552 30340 34561
rect 31668 34731 31720 34740
rect 31668 34697 31677 34731
rect 31677 34697 31711 34731
rect 31711 34697 31720 34731
rect 31668 34688 31720 34697
rect 31760 34620 31812 34672
rect 30656 34552 30708 34604
rect 31024 34595 31076 34604
rect 31024 34561 31033 34595
rect 31033 34561 31067 34595
rect 31067 34561 31076 34595
rect 31024 34552 31076 34561
rect 29920 34484 29972 34536
rect 30472 34416 30524 34468
rect 30656 34416 30708 34468
rect 32036 34552 32088 34604
rect 32404 34595 32456 34604
rect 32404 34561 32413 34595
rect 32413 34561 32447 34595
rect 32447 34561 32456 34595
rect 32404 34552 32456 34561
rect 31944 34484 31996 34536
rect 32128 34527 32180 34536
rect 32128 34493 32137 34527
rect 32137 34493 32171 34527
rect 32171 34493 32180 34527
rect 32128 34484 32180 34493
rect 32772 34484 32824 34536
rect 33140 34484 33192 34536
rect 31208 34391 31260 34400
rect 31208 34357 31217 34391
rect 31217 34357 31251 34391
rect 31251 34357 31260 34391
rect 31208 34348 31260 34357
rect 38476 34391 38528 34400
rect 38476 34357 38485 34391
rect 38485 34357 38519 34391
rect 38519 34357 38528 34391
rect 38476 34348 38528 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5632 34187 5684 34196
rect 5632 34153 5641 34187
rect 5641 34153 5675 34187
rect 5675 34153 5684 34187
rect 5632 34144 5684 34153
rect 7380 34144 7432 34196
rect 13084 34187 13136 34196
rect 13084 34153 13093 34187
rect 13093 34153 13127 34187
rect 13127 34153 13136 34187
rect 13084 34144 13136 34153
rect 13452 34144 13504 34196
rect 13636 34144 13688 34196
rect 15292 34187 15344 34196
rect 15292 34153 15301 34187
rect 15301 34153 15335 34187
rect 15335 34153 15344 34187
rect 15292 34144 15344 34153
rect 18328 34144 18380 34196
rect 29184 34187 29236 34196
rect 29184 34153 29193 34187
rect 29193 34153 29227 34187
rect 29227 34153 29236 34187
rect 29184 34144 29236 34153
rect 30656 34144 30708 34196
rect 3240 33940 3292 33992
rect 5080 34051 5132 34060
rect 5080 34017 5089 34051
rect 5089 34017 5123 34051
rect 5123 34017 5132 34051
rect 5080 34008 5132 34017
rect 6092 34076 6144 34128
rect 3424 33983 3476 33992
rect 3424 33949 3433 33983
rect 3433 33949 3467 33983
rect 3467 33949 3476 33983
rect 3424 33940 3476 33949
rect 4528 33983 4580 33992
rect 4528 33949 4537 33983
rect 4537 33949 4571 33983
rect 4571 33949 4580 33983
rect 4528 33940 4580 33949
rect 5356 33940 5408 33992
rect 10324 34008 10376 34060
rect 11060 34008 11112 34060
rect 12164 34008 12216 34060
rect 6920 33983 6972 33992
rect 6920 33949 6929 33983
rect 6929 33949 6963 33983
rect 6963 33949 6972 33983
rect 6920 33940 6972 33949
rect 13544 33940 13596 33992
rect 15016 33983 15068 33992
rect 15016 33949 15025 33983
rect 15025 33949 15059 33983
rect 15059 33949 15068 33983
rect 15016 33940 15068 33949
rect 15752 34008 15804 34060
rect 16212 34051 16264 34060
rect 16212 34017 16221 34051
rect 16221 34017 16255 34051
rect 16255 34017 16264 34051
rect 16212 34008 16264 34017
rect 17408 34008 17460 34060
rect 19248 34051 19300 34060
rect 19248 34017 19257 34051
rect 19257 34017 19291 34051
rect 19291 34017 19300 34051
rect 19248 34008 19300 34017
rect 21732 34051 21784 34060
rect 21732 34017 21741 34051
rect 21741 34017 21775 34051
rect 21775 34017 21784 34051
rect 21732 34008 21784 34017
rect 22192 34008 22244 34060
rect 23204 34008 23256 34060
rect 24860 34008 24912 34060
rect 25504 34008 25556 34060
rect 27436 34051 27488 34060
rect 27436 34017 27445 34051
rect 27445 34017 27479 34051
rect 27479 34017 27488 34051
rect 27436 34008 27488 34017
rect 30380 34008 30432 34060
rect 17868 33940 17920 33992
rect 30472 33983 30524 33992
rect 30472 33949 30481 33983
rect 30481 33949 30515 33983
rect 30515 33949 30524 33983
rect 30472 33940 30524 33949
rect 31760 34008 31812 34060
rect 33140 34008 33192 34060
rect 6092 33872 6144 33924
rect 8760 33872 8812 33924
rect 11612 33915 11664 33924
rect 11612 33881 11621 33915
rect 11621 33881 11655 33915
rect 11655 33881 11664 33915
rect 11612 33872 11664 33881
rect 13084 33872 13136 33924
rect 13912 33872 13964 33924
rect 17592 33872 17644 33924
rect 19524 33915 19576 33924
rect 19524 33881 19533 33915
rect 19533 33881 19567 33915
rect 19567 33881 19576 33915
rect 19524 33872 19576 33881
rect 19984 33872 20036 33924
rect 22284 33872 22336 33924
rect 2504 33804 2556 33856
rect 5448 33847 5500 33856
rect 5448 33813 5457 33847
rect 5457 33813 5491 33847
rect 5491 33813 5500 33847
rect 5448 33804 5500 33813
rect 5724 33804 5776 33856
rect 7012 33804 7064 33856
rect 8024 33804 8076 33856
rect 9220 33847 9272 33856
rect 9220 33813 9229 33847
rect 9229 33813 9263 33847
rect 9263 33813 9272 33847
rect 9220 33804 9272 33813
rect 17040 33804 17092 33856
rect 20352 33804 20404 33856
rect 21180 33847 21232 33856
rect 21180 33813 21189 33847
rect 21189 33813 21223 33847
rect 21223 33813 21232 33847
rect 21180 33804 21232 33813
rect 21364 33804 21416 33856
rect 21916 33804 21968 33856
rect 27712 33915 27764 33924
rect 27712 33881 27721 33915
rect 27721 33881 27755 33915
rect 27755 33881 27764 33915
rect 27712 33872 27764 33881
rect 27988 33872 28040 33924
rect 29828 33872 29880 33924
rect 23664 33847 23716 33856
rect 23664 33813 23673 33847
rect 23673 33813 23707 33847
rect 23707 33813 23716 33847
rect 23664 33804 23716 33813
rect 25044 33804 25096 33856
rect 25228 33804 25280 33856
rect 28080 33804 28132 33856
rect 30380 33847 30432 33856
rect 30380 33813 30389 33847
rect 30389 33813 30423 33847
rect 30423 33813 30432 33847
rect 30380 33804 30432 33813
rect 30656 33847 30708 33856
rect 30656 33813 30665 33847
rect 30665 33813 30699 33847
rect 30699 33813 30708 33847
rect 30656 33804 30708 33813
rect 34796 33804 34848 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 3424 33600 3476 33652
rect 2504 33575 2556 33584
rect 2504 33541 2513 33575
rect 2513 33541 2547 33575
rect 2547 33541 2556 33575
rect 2504 33532 2556 33541
rect 3792 33532 3844 33584
rect 7104 33600 7156 33652
rect 10232 33600 10284 33652
rect 7012 33532 7064 33584
rect 9680 33532 9732 33584
rect 9772 33532 9824 33584
rect 10416 33532 10468 33584
rect 4620 33507 4672 33516
rect 4620 33473 4629 33507
rect 4629 33473 4663 33507
rect 4663 33473 4672 33507
rect 4620 33464 4672 33473
rect 4712 33507 4764 33516
rect 4712 33473 4721 33507
rect 4721 33473 4755 33507
rect 4755 33473 4764 33507
rect 4712 33464 4764 33473
rect 2228 33439 2280 33448
rect 2228 33405 2237 33439
rect 2237 33405 2271 33439
rect 2271 33405 2280 33439
rect 2228 33396 2280 33405
rect 4528 33439 4580 33448
rect 4528 33405 4537 33439
rect 4537 33405 4571 33439
rect 4571 33405 4580 33439
rect 4528 33396 4580 33405
rect 5632 33396 5684 33448
rect 7288 33507 7340 33516
rect 7288 33473 7297 33507
rect 7297 33473 7331 33507
rect 7331 33473 7340 33507
rect 7288 33464 7340 33473
rect 8116 33464 8168 33516
rect 11060 33575 11112 33584
rect 11060 33541 11069 33575
rect 11069 33541 11103 33575
rect 11103 33541 11112 33575
rect 11060 33532 11112 33541
rect 21180 33600 21232 33652
rect 22468 33600 22520 33652
rect 21824 33532 21876 33584
rect 23664 33600 23716 33652
rect 10968 33464 11020 33516
rect 7472 33396 7524 33448
rect 8852 33396 8904 33448
rect 9220 33396 9272 33448
rect 9496 33439 9548 33448
rect 9496 33405 9505 33439
rect 9505 33405 9539 33439
rect 9539 33405 9548 33439
rect 9496 33396 9548 33405
rect 15568 33507 15620 33516
rect 15568 33473 15577 33507
rect 15577 33473 15611 33507
rect 15611 33473 15620 33507
rect 15568 33464 15620 33473
rect 18696 33464 18748 33516
rect 21272 33464 21324 33516
rect 23204 33575 23256 33584
rect 23204 33541 23213 33575
rect 23213 33541 23247 33575
rect 23247 33541 23256 33575
rect 23204 33532 23256 33541
rect 16304 33396 16356 33448
rect 19340 33396 19392 33448
rect 22468 33464 22520 33516
rect 23020 33464 23072 33516
rect 23480 33507 23532 33516
rect 23480 33473 23489 33507
rect 23489 33473 23523 33507
rect 23523 33473 23532 33507
rect 23480 33464 23532 33473
rect 23940 33600 23992 33652
rect 27712 33600 27764 33652
rect 28448 33600 28500 33652
rect 29276 33643 29328 33652
rect 29276 33609 29285 33643
rect 29285 33609 29319 33643
rect 29319 33609 29328 33643
rect 29276 33600 29328 33609
rect 30380 33600 30432 33652
rect 24860 33507 24912 33516
rect 24860 33473 24869 33507
rect 24869 33473 24903 33507
rect 24903 33473 24912 33507
rect 24860 33464 24912 33473
rect 27160 33464 27212 33516
rect 27344 33464 27396 33516
rect 27896 33507 27948 33516
rect 27896 33473 27905 33507
rect 27905 33473 27939 33507
rect 27939 33473 27948 33507
rect 27896 33464 27948 33473
rect 29000 33532 29052 33584
rect 29736 33532 29788 33584
rect 34796 33532 34848 33584
rect 35532 33532 35584 33584
rect 28080 33464 28132 33516
rect 28264 33507 28316 33516
rect 28264 33473 28273 33507
rect 28273 33473 28307 33507
rect 28307 33473 28316 33507
rect 28264 33464 28316 33473
rect 28724 33464 28776 33516
rect 29184 33507 29236 33516
rect 29184 33473 29193 33507
rect 29193 33473 29227 33507
rect 29227 33473 29236 33507
rect 29184 33464 29236 33473
rect 33140 33464 33192 33516
rect 3240 33260 3292 33312
rect 4896 33303 4948 33312
rect 4896 33269 4905 33303
rect 4905 33269 4939 33303
rect 4939 33269 4948 33303
rect 4896 33260 4948 33269
rect 5724 33260 5776 33312
rect 6000 33260 6052 33312
rect 8576 33260 8628 33312
rect 22836 33328 22888 33380
rect 23480 33328 23532 33380
rect 15384 33303 15436 33312
rect 15384 33269 15393 33303
rect 15393 33269 15427 33303
rect 15427 33269 15436 33303
rect 15384 33260 15436 33269
rect 18696 33303 18748 33312
rect 18696 33269 18705 33303
rect 18705 33269 18739 33303
rect 18739 33269 18748 33303
rect 18696 33260 18748 33269
rect 22008 33260 22060 33312
rect 23296 33260 23348 33312
rect 29276 33396 29328 33448
rect 26240 33328 26292 33380
rect 29552 33328 29604 33380
rect 31024 33439 31076 33448
rect 31024 33405 31033 33439
rect 31033 33405 31067 33439
rect 31067 33405 31076 33439
rect 31024 33396 31076 33405
rect 26516 33260 26568 33312
rect 26608 33303 26660 33312
rect 26608 33269 26617 33303
rect 26617 33269 26651 33303
rect 26651 33269 26660 33303
rect 26608 33260 26660 33269
rect 27068 33303 27120 33312
rect 27068 33269 27077 33303
rect 27077 33269 27111 33303
rect 27111 33269 27120 33303
rect 27068 33260 27120 33269
rect 27988 33260 28040 33312
rect 28448 33260 28500 33312
rect 30748 33260 30800 33312
rect 33508 33439 33560 33448
rect 33508 33405 33517 33439
rect 33517 33405 33551 33439
rect 33551 33405 33560 33439
rect 33508 33396 33560 33405
rect 33600 33396 33652 33448
rect 34244 33396 34296 33448
rect 34520 33328 34572 33380
rect 38476 33371 38528 33380
rect 38476 33337 38485 33371
rect 38485 33337 38519 33371
rect 38519 33337 38528 33371
rect 38476 33328 38528 33337
rect 34796 33260 34848 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 3424 32895 3476 32904
rect 3424 32861 3433 32895
rect 3433 32861 3467 32895
rect 3467 32861 3476 32895
rect 3424 32852 3476 32861
rect 4896 33056 4948 33108
rect 9680 33099 9732 33108
rect 9680 33065 9689 33099
rect 9689 33065 9723 33099
rect 9723 33065 9732 33099
rect 9680 33056 9732 33065
rect 10784 33056 10836 33108
rect 10968 33099 11020 33108
rect 10968 33065 10977 33099
rect 10977 33065 11011 33099
rect 11011 33065 11020 33099
rect 10968 33056 11020 33065
rect 11796 33056 11848 33108
rect 17040 33099 17092 33108
rect 17040 33065 17049 33099
rect 17049 33065 17083 33099
rect 17083 33065 17092 33099
rect 17040 33056 17092 33065
rect 18144 33099 18196 33108
rect 18144 33065 18153 33099
rect 18153 33065 18187 33099
rect 18187 33065 18196 33099
rect 18144 33056 18196 33065
rect 19524 33056 19576 33108
rect 3884 32963 3936 32972
rect 3884 32929 3893 32963
rect 3893 32929 3927 32963
rect 3927 32929 3936 32963
rect 3884 32920 3936 32929
rect 6000 32963 6052 32972
rect 6000 32929 6009 32963
rect 6009 32929 6043 32963
rect 6043 32929 6052 32963
rect 6000 32920 6052 32929
rect 7288 32920 7340 32972
rect 8852 32920 8904 32972
rect 3700 32716 3752 32768
rect 3976 32716 4028 32768
rect 7012 32784 7064 32836
rect 8024 32852 8076 32904
rect 5632 32759 5684 32768
rect 5632 32725 5641 32759
rect 5641 32725 5675 32759
rect 5675 32725 5684 32759
rect 5632 32716 5684 32725
rect 7472 32759 7524 32768
rect 7472 32725 7481 32759
rect 7481 32725 7515 32759
rect 7515 32725 7524 32759
rect 7472 32716 7524 32725
rect 7564 32759 7616 32768
rect 7564 32725 7573 32759
rect 7573 32725 7607 32759
rect 7607 32725 7616 32759
rect 7564 32716 7616 32725
rect 8576 32895 8628 32904
rect 8576 32861 8585 32895
rect 8585 32861 8619 32895
rect 8619 32861 8628 32895
rect 8576 32852 8628 32861
rect 9956 32852 10008 32904
rect 11060 32988 11112 33040
rect 15568 32988 15620 33040
rect 15936 32988 15988 33040
rect 20444 32988 20496 33040
rect 22284 33056 22336 33108
rect 25504 33056 25556 33108
rect 26240 33099 26292 33108
rect 26240 33065 26249 33099
rect 26249 33065 26283 33099
rect 26283 33065 26292 33099
rect 26240 33056 26292 33065
rect 27896 33056 27948 33108
rect 28632 33056 28684 33108
rect 30656 33099 30708 33108
rect 30656 33065 30665 33099
rect 30665 33065 30699 33099
rect 30699 33065 30708 33099
rect 30656 33056 30708 33065
rect 31668 33056 31720 33108
rect 32772 33056 32824 33108
rect 33508 33056 33560 33108
rect 11060 32852 11112 32904
rect 18696 32920 18748 32972
rect 20352 32963 20404 32972
rect 20352 32929 20361 32963
rect 20361 32929 20395 32963
rect 20395 32929 20404 32963
rect 20352 32920 20404 32929
rect 14188 32852 14240 32904
rect 16304 32895 16356 32904
rect 16304 32861 16313 32895
rect 16313 32861 16347 32895
rect 16347 32861 16356 32895
rect 16304 32852 16356 32861
rect 17500 32895 17552 32904
rect 17500 32861 17509 32895
rect 17509 32861 17543 32895
rect 17543 32861 17552 32895
rect 17500 32852 17552 32861
rect 11336 32827 11388 32836
rect 11336 32793 11345 32827
rect 11345 32793 11379 32827
rect 11379 32793 11388 32827
rect 11336 32784 11388 32793
rect 12164 32784 12216 32836
rect 13084 32784 13136 32836
rect 13544 32784 13596 32836
rect 13636 32784 13688 32836
rect 14924 32784 14976 32836
rect 11152 32759 11204 32768
rect 11152 32725 11179 32759
rect 11179 32725 11204 32759
rect 11152 32716 11204 32725
rect 14648 32716 14700 32768
rect 16948 32716 17000 32768
rect 17684 32895 17736 32904
rect 17684 32861 17693 32895
rect 17693 32861 17727 32895
rect 17727 32861 17736 32895
rect 17684 32852 17736 32861
rect 18144 32852 18196 32904
rect 19340 32895 19392 32904
rect 19340 32861 19349 32895
rect 19349 32861 19383 32895
rect 19383 32861 19392 32895
rect 19340 32852 19392 32861
rect 23296 32988 23348 33040
rect 27436 32988 27488 33040
rect 26608 32920 26660 32972
rect 22192 32852 22244 32904
rect 27160 32852 27212 32904
rect 27252 32895 27304 32904
rect 27252 32861 27261 32895
rect 27261 32861 27295 32895
rect 27295 32861 27304 32895
rect 27252 32852 27304 32861
rect 28356 32988 28408 33040
rect 28540 32988 28592 33040
rect 35532 33056 35584 33108
rect 27804 32920 27856 32972
rect 28724 32895 28776 32904
rect 28724 32861 28733 32895
rect 28733 32861 28767 32895
rect 28767 32861 28776 32895
rect 28724 32852 28776 32861
rect 17776 32716 17828 32768
rect 23940 32784 23992 32836
rect 24216 32784 24268 32836
rect 25596 32784 25648 32836
rect 25964 32784 26016 32836
rect 18236 32716 18288 32768
rect 22008 32759 22060 32768
rect 22008 32725 22033 32759
rect 22033 32725 22060 32759
rect 22008 32716 22060 32725
rect 26700 32759 26752 32768
rect 26700 32725 26709 32759
rect 26709 32725 26743 32759
rect 26743 32725 26752 32759
rect 26700 32716 26752 32725
rect 28264 32784 28316 32836
rect 29552 32895 29604 32904
rect 29552 32861 29561 32895
rect 29561 32861 29595 32895
rect 29595 32861 29604 32895
rect 29552 32852 29604 32861
rect 30748 32895 30800 32904
rect 30748 32861 30757 32895
rect 30757 32861 30791 32895
rect 30791 32861 30800 32895
rect 30748 32852 30800 32861
rect 31024 32920 31076 32972
rect 31668 32852 31720 32904
rect 33324 32920 33376 32972
rect 34336 32988 34388 33040
rect 33876 32895 33928 32904
rect 33876 32861 33885 32895
rect 33885 32861 33919 32895
rect 33919 32861 33928 32895
rect 33876 32852 33928 32861
rect 34244 32895 34296 32904
rect 34244 32861 34253 32895
rect 34253 32861 34287 32895
rect 34287 32861 34296 32895
rect 34244 32852 34296 32861
rect 34796 32920 34848 32972
rect 35532 32920 35584 32972
rect 34612 32852 34664 32904
rect 30012 32784 30064 32836
rect 31024 32784 31076 32836
rect 32128 32784 32180 32836
rect 36176 32784 36228 32836
rect 27988 32716 28040 32768
rect 28172 32759 28224 32768
rect 28172 32725 28181 32759
rect 28181 32725 28215 32759
rect 28215 32725 28224 32759
rect 28172 32716 28224 32725
rect 33508 32759 33560 32768
rect 33508 32725 33517 32759
rect 33517 32725 33551 32759
rect 33551 32725 33560 32759
rect 33508 32716 33560 32725
rect 34520 32716 34572 32768
rect 36728 32716 36780 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 3976 32555 4028 32564
rect 3976 32521 4011 32555
rect 4011 32521 4028 32555
rect 3976 32512 4028 32521
rect 4528 32512 4580 32564
rect 4712 32512 4764 32564
rect 6920 32555 6972 32564
rect 6920 32521 6929 32555
rect 6929 32521 6963 32555
rect 6963 32521 6972 32555
rect 6920 32512 6972 32521
rect 7104 32555 7156 32564
rect 7104 32521 7113 32555
rect 7113 32521 7147 32555
rect 7147 32521 7156 32555
rect 7104 32512 7156 32521
rect 11796 32555 11848 32564
rect 11796 32521 11805 32555
rect 11805 32521 11839 32555
rect 11839 32521 11848 32555
rect 11796 32512 11848 32521
rect 12624 32512 12676 32564
rect 7472 32444 7524 32496
rect 9772 32444 9824 32496
rect 14188 32555 14240 32564
rect 14188 32521 14197 32555
rect 14197 32521 14231 32555
rect 14231 32521 14240 32555
rect 14188 32512 14240 32521
rect 13636 32444 13688 32496
rect 15660 32512 15712 32564
rect 16304 32512 16356 32564
rect 6644 32419 6696 32428
rect 6644 32385 6653 32419
rect 6653 32385 6687 32419
rect 6687 32385 6696 32419
rect 6644 32376 6696 32385
rect 6920 32376 6972 32428
rect 7564 32376 7616 32428
rect 9496 32376 9548 32428
rect 13544 32419 13596 32428
rect 13544 32385 13553 32419
rect 13553 32385 13587 32419
rect 13587 32385 13596 32419
rect 13544 32376 13596 32385
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 14648 32487 14700 32496
rect 14648 32453 14657 32487
rect 14657 32453 14691 32487
rect 14691 32453 14700 32487
rect 14648 32444 14700 32453
rect 14924 32444 14976 32496
rect 19340 32512 19392 32564
rect 23756 32512 23808 32564
rect 24308 32512 24360 32564
rect 24676 32512 24728 32564
rect 16948 32487 17000 32496
rect 16948 32453 16957 32487
rect 16957 32453 16991 32487
rect 16991 32453 17000 32487
rect 16948 32444 17000 32453
rect 18512 32487 18564 32496
rect 18512 32453 18521 32487
rect 18521 32453 18555 32487
rect 18555 32453 18564 32487
rect 18512 32444 18564 32453
rect 18880 32444 18932 32496
rect 21916 32444 21968 32496
rect 23664 32444 23716 32496
rect 4620 32308 4672 32360
rect 4804 32308 4856 32360
rect 3424 32240 3476 32292
rect 5632 32308 5684 32360
rect 10232 32308 10284 32360
rect 12532 32308 12584 32360
rect 15384 32308 15436 32360
rect 16396 32308 16448 32360
rect 18236 32376 18288 32428
rect 19156 32419 19208 32428
rect 19156 32385 19165 32419
rect 19165 32385 19199 32419
rect 19199 32385 19208 32419
rect 19156 32376 19208 32385
rect 22100 32419 22152 32428
rect 22100 32385 22109 32419
rect 22109 32385 22143 32419
rect 22143 32385 22152 32419
rect 22100 32376 22152 32385
rect 25136 32444 25188 32496
rect 25596 32555 25648 32564
rect 25596 32521 25605 32555
rect 25605 32521 25639 32555
rect 25639 32521 25648 32555
rect 25596 32512 25648 32521
rect 26700 32512 26752 32564
rect 27896 32512 27948 32564
rect 28724 32512 28776 32564
rect 32128 32555 32180 32564
rect 32128 32521 32137 32555
rect 32137 32521 32171 32555
rect 32171 32521 32180 32555
rect 32128 32512 32180 32521
rect 22376 32351 22428 32360
rect 22376 32317 22385 32351
rect 22385 32317 22419 32351
rect 22419 32317 22428 32351
rect 22376 32308 22428 32317
rect 23848 32351 23900 32360
rect 23848 32317 23857 32351
rect 23857 32317 23891 32351
rect 23891 32317 23900 32351
rect 24676 32419 24728 32428
rect 24676 32385 24685 32419
rect 24685 32385 24719 32419
rect 24719 32385 24728 32419
rect 24676 32376 24728 32385
rect 25044 32419 25096 32428
rect 25044 32385 25054 32419
rect 25054 32385 25088 32419
rect 25088 32385 25096 32419
rect 25044 32376 25096 32385
rect 25228 32419 25280 32428
rect 25228 32385 25237 32419
rect 25237 32385 25271 32419
rect 25271 32385 25280 32419
rect 25228 32376 25280 32385
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 23848 32308 23900 32317
rect 6276 32240 6328 32292
rect 5356 32172 5408 32224
rect 11336 32215 11388 32224
rect 11336 32181 11345 32215
rect 11345 32181 11379 32215
rect 11379 32181 11388 32215
rect 11336 32172 11388 32181
rect 17500 32172 17552 32224
rect 17960 32172 18012 32224
rect 18144 32172 18196 32224
rect 20720 32172 20772 32224
rect 25964 32376 26016 32428
rect 26424 32376 26476 32428
rect 27068 32376 27120 32428
rect 28080 32444 28132 32496
rect 29276 32444 29328 32496
rect 33876 32555 33928 32564
rect 33876 32521 33885 32555
rect 33885 32521 33919 32555
rect 33919 32521 33928 32555
rect 33876 32512 33928 32521
rect 34612 32555 34664 32564
rect 34612 32521 34621 32555
rect 34621 32521 34655 32555
rect 34655 32521 34664 32555
rect 34612 32512 34664 32521
rect 27804 32419 27856 32428
rect 27804 32385 27813 32419
rect 27813 32385 27847 32419
rect 27847 32385 27856 32419
rect 27804 32376 27856 32385
rect 28172 32376 28224 32428
rect 30012 32419 30064 32428
rect 30012 32385 30021 32419
rect 30021 32385 30055 32419
rect 30055 32385 30064 32419
rect 30012 32376 30064 32385
rect 30288 32376 30340 32428
rect 31392 32419 31444 32428
rect 31392 32385 31401 32419
rect 31401 32385 31435 32419
rect 31435 32385 31444 32419
rect 31392 32376 31444 32385
rect 31760 32419 31812 32428
rect 31760 32385 31769 32419
rect 31769 32385 31803 32419
rect 31803 32385 31812 32419
rect 31760 32376 31812 32385
rect 28080 32308 28132 32360
rect 26700 32240 26752 32292
rect 30564 32308 30616 32360
rect 24492 32172 24544 32224
rect 27344 32215 27396 32224
rect 27344 32181 27353 32215
rect 27353 32181 27387 32215
rect 27387 32181 27396 32215
rect 27344 32172 27396 32181
rect 33508 32419 33560 32428
rect 33508 32385 33517 32419
rect 33517 32385 33551 32419
rect 33551 32385 33560 32419
rect 33508 32376 33560 32385
rect 33600 32419 33652 32428
rect 33600 32385 33609 32419
rect 33609 32385 33643 32419
rect 33643 32385 33652 32419
rect 33600 32376 33652 32385
rect 33876 32376 33928 32428
rect 33140 32351 33192 32360
rect 33140 32317 33149 32351
rect 33149 32317 33183 32351
rect 33183 32317 33192 32351
rect 33140 32308 33192 32317
rect 33324 32240 33376 32292
rect 28264 32172 28316 32224
rect 30656 32172 30708 32224
rect 33416 32172 33468 32224
rect 36728 32376 36780 32428
rect 34612 32351 34664 32360
rect 34612 32317 34621 32351
rect 34621 32317 34655 32351
rect 34655 32317 34664 32351
rect 34612 32308 34664 32317
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2228 31968 2280 32020
rect 2504 31968 2556 32020
rect 6644 31968 6696 32020
rect 10232 32011 10284 32020
rect 10232 31977 10241 32011
rect 10241 31977 10275 32011
rect 10275 31977 10284 32011
rect 10232 31968 10284 31977
rect 10508 31968 10560 32020
rect 10876 31968 10928 32020
rect 2504 31832 2556 31884
rect 4620 31900 4672 31952
rect 6276 31943 6328 31952
rect 6276 31909 6285 31943
rect 6285 31909 6319 31943
rect 6319 31909 6328 31943
rect 6276 31900 6328 31909
rect 3792 31764 3844 31816
rect 6552 31875 6604 31884
rect 6552 31841 6561 31875
rect 6561 31841 6595 31875
rect 6595 31841 6604 31875
rect 6552 31832 6604 31841
rect 6920 31832 6972 31884
rect 7288 31832 7340 31884
rect 10508 31832 10560 31884
rect 4068 31696 4120 31748
rect 6736 31807 6788 31816
rect 6736 31773 6745 31807
rect 6745 31773 6779 31807
rect 6779 31773 6788 31807
rect 6736 31764 6788 31773
rect 7564 31764 7616 31816
rect 7748 31764 7800 31816
rect 10416 31807 10468 31816
rect 10416 31773 10425 31807
rect 10425 31773 10459 31807
rect 10459 31773 10468 31807
rect 10416 31764 10468 31773
rect 11152 31900 11204 31952
rect 12532 32011 12584 32020
rect 12532 31977 12541 32011
rect 12541 31977 12575 32011
rect 12575 31977 12584 32011
rect 12532 31968 12584 31977
rect 15384 31968 15436 32020
rect 11336 31832 11388 31884
rect 7196 31696 7248 31748
rect 7288 31739 7340 31748
rect 7288 31705 7297 31739
rect 7297 31705 7331 31739
rect 7331 31705 7340 31739
rect 7288 31696 7340 31705
rect 7656 31696 7708 31748
rect 10692 31696 10744 31748
rect 10968 31739 11020 31748
rect 10968 31705 10977 31739
rect 10977 31705 11011 31739
rect 11011 31705 11020 31739
rect 10968 31696 11020 31705
rect 5816 31671 5868 31680
rect 5816 31637 5825 31671
rect 5825 31637 5859 31671
rect 5859 31637 5868 31671
rect 5816 31628 5868 31637
rect 6736 31628 6788 31680
rect 7564 31671 7616 31680
rect 7564 31637 7573 31671
rect 7573 31637 7607 31671
rect 7607 31637 7616 31671
rect 7564 31628 7616 31637
rect 11796 31696 11848 31748
rect 12440 31807 12492 31816
rect 12440 31773 12449 31807
rect 12449 31773 12483 31807
rect 12483 31773 12492 31807
rect 12440 31764 12492 31773
rect 15292 31832 15344 31884
rect 15200 31764 15252 31816
rect 17040 31968 17092 32020
rect 18512 31968 18564 32020
rect 18880 31968 18932 32020
rect 25320 31968 25372 32020
rect 25596 31968 25648 32020
rect 17684 31900 17736 31952
rect 17776 31900 17828 31952
rect 17500 31832 17552 31884
rect 18236 31943 18288 31952
rect 18236 31909 18245 31943
rect 18245 31909 18279 31943
rect 18279 31909 18288 31943
rect 18236 31900 18288 31909
rect 11704 31671 11756 31680
rect 11704 31637 11713 31671
rect 11713 31637 11747 31671
rect 11747 31637 11756 31671
rect 11704 31628 11756 31637
rect 14372 31628 14424 31680
rect 15936 31739 15988 31748
rect 15936 31705 15961 31739
rect 15961 31705 15988 31739
rect 15936 31696 15988 31705
rect 16304 31696 16356 31748
rect 18144 31764 18196 31816
rect 18236 31764 18288 31816
rect 19156 31832 19208 31884
rect 20076 31832 20128 31884
rect 20720 31875 20772 31884
rect 20720 31841 20729 31875
rect 20729 31841 20763 31875
rect 20763 31841 20772 31875
rect 20720 31832 20772 31841
rect 24768 31900 24820 31952
rect 23664 31832 23716 31884
rect 26608 31832 26660 31884
rect 20996 31807 21048 31816
rect 20996 31773 21005 31807
rect 21005 31773 21039 31807
rect 21039 31773 21048 31807
rect 20996 31764 21048 31773
rect 23572 31764 23624 31816
rect 24952 31807 25004 31816
rect 24952 31773 24961 31807
rect 24961 31773 24995 31807
rect 24995 31773 25004 31807
rect 24952 31764 25004 31773
rect 25044 31764 25096 31816
rect 26700 31807 26752 31816
rect 26700 31773 26709 31807
rect 26709 31773 26743 31807
rect 26743 31773 26752 31807
rect 26700 31764 26752 31773
rect 27804 31968 27856 32020
rect 28080 31968 28132 32020
rect 31392 31968 31444 32020
rect 33232 31968 33284 32020
rect 33600 31968 33652 32020
rect 27620 31900 27672 31952
rect 27344 31832 27396 31884
rect 27988 31832 28040 31884
rect 27804 31807 27856 31816
rect 17684 31739 17736 31748
rect 17684 31705 17693 31739
rect 17693 31705 17727 31739
rect 17727 31705 17736 31739
rect 17684 31696 17736 31705
rect 19984 31696 20036 31748
rect 22008 31696 22060 31748
rect 22100 31696 22152 31748
rect 22560 31696 22612 31748
rect 16120 31671 16172 31680
rect 16120 31637 16129 31671
rect 16129 31637 16163 31671
rect 16163 31637 16172 31671
rect 16120 31628 16172 31637
rect 18604 31671 18656 31680
rect 18604 31637 18613 31671
rect 18613 31637 18647 31671
rect 18647 31637 18656 31671
rect 18604 31628 18656 31637
rect 22192 31628 22244 31680
rect 22836 31628 22888 31680
rect 24400 31671 24452 31680
rect 24400 31637 24409 31671
rect 24409 31637 24443 31671
rect 24443 31637 24452 31671
rect 24400 31628 24452 31637
rect 27804 31773 27813 31807
rect 27813 31773 27847 31807
rect 27847 31773 27856 31807
rect 27804 31764 27856 31773
rect 28264 31764 28316 31816
rect 30288 31832 30340 31884
rect 30656 31875 30708 31884
rect 30656 31841 30665 31875
rect 30665 31841 30699 31875
rect 30699 31841 30708 31875
rect 30656 31832 30708 31841
rect 28632 31807 28684 31816
rect 28632 31773 28641 31807
rect 28641 31773 28675 31807
rect 28675 31773 28684 31807
rect 28632 31764 28684 31773
rect 31852 31832 31904 31884
rect 32772 31764 32824 31816
rect 34704 31764 34756 31816
rect 36636 31764 36688 31816
rect 38476 31807 38528 31816
rect 38476 31773 38485 31807
rect 38485 31773 38519 31807
rect 38519 31773 38528 31807
rect 38476 31764 38528 31773
rect 28356 31628 28408 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 3792 31424 3844 31476
rect 6736 31467 6788 31476
rect 6736 31433 6745 31467
rect 6745 31433 6779 31467
rect 6779 31433 6788 31467
rect 6736 31424 6788 31433
rect 6828 31424 6880 31476
rect 7748 31467 7800 31476
rect 7748 31433 7757 31467
rect 7757 31433 7791 31467
rect 7791 31433 7800 31467
rect 7748 31424 7800 31433
rect 12440 31424 12492 31476
rect 14096 31424 14148 31476
rect 5724 31356 5776 31408
rect 7196 31356 7248 31408
rect 12624 31356 12676 31408
rect 13360 31356 13412 31408
rect 15200 31424 15252 31476
rect 15292 31467 15344 31476
rect 15292 31433 15301 31467
rect 15301 31433 15335 31467
rect 15335 31433 15344 31467
rect 15292 31424 15344 31433
rect 16212 31424 16264 31476
rect 17040 31467 17092 31476
rect 17040 31433 17049 31467
rect 17049 31433 17083 31467
rect 17083 31433 17092 31467
rect 17040 31424 17092 31433
rect 18236 31424 18288 31476
rect 18604 31467 18656 31476
rect 18604 31433 18613 31467
rect 18613 31433 18647 31467
rect 18647 31433 18656 31467
rect 18604 31424 18656 31433
rect 19984 31424 20036 31476
rect 22008 31424 22060 31476
rect 2228 31288 2280 31340
rect 5816 31331 5868 31340
rect 3608 31263 3660 31272
rect 3608 31229 3617 31263
rect 3617 31229 3651 31263
rect 3651 31229 3660 31263
rect 3608 31220 3660 31229
rect 5816 31297 5825 31331
rect 5825 31297 5859 31331
rect 5859 31297 5868 31331
rect 5816 31288 5868 31297
rect 6644 31331 6696 31340
rect 6644 31297 6653 31331
rect 6653 31297 6687 31331
rect 6687 31297 6696 31331
rect 6644 31288 6696 31297
rect 6828 31288 6880 31340
rect 7564 31288 7616 31340
rect 8116 31288 8168 31340
rect 7380 31263 7432 31272
rect 7380 31229 7389 31263
rect 7389 31229 7423 31263
rect 7423 31229 7432 31263
rect 7380 31220 7432 31229
rect 4620 31152 4672 31204
rect 7288 31152 7340 31204
rect 9496 31263 9548 31272
rect 9496 31229 9505 31263
rect 9505 31229 9539 31263
rect 9539 31229 9548 31263
rect 9496 31220 9548 31229
rect 10416 31220 10468 31272
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 12348 31288 12400 31340
rect 13084 31331 13136 31340
rect 13084 31297 13093 31331
rect 13093 31297 13127 31331
rect 13127 31297 13136 31331
rect 13084 31288 13136 31297
rect 16120 31356 16172 31408
rect 11152 31220 11204 31272
rect 11796 31263 11848 31272
rect 11796 31229 11805 31263
rect 11805 31229 11839 31263
rect 11839 31229 11848 31263
rect 11796 31220 11848 31229
rect 14372 31220 14424 31272
rect 16212 31331 16264 31340
rect 16212 31297 16221 31331
rect 16221 31297 16255 31331
rect 16255 31297 16264 31331
rect 16212 31288 16264 31297
rect 17684 31356 17736 31408
rect 20076 31356 20128 31408
rect 16948 31331 17000 31340
rect 16948 31297 16957 31331
rect 16957 31297 16991 31331
rect 16991 31297 17000 31331
rect 16948 31288 17000 31297
rect 4804 31084 4856 31136
rect 5448 31084 5500 31136
rect 10140 31084 10192 31136
rect 11244 31084 11296 31136
rect 13912 31084 13964 31136
rect 16120 31220 16172 31272
rect 16396 31220 16448 31272
rect 17960 31331 18012 31340
rect 17960 31297 17969 31331
rect 17969 31297 18003 31331
rect 18003 31297 18012 31331
rect 17960 31288 18012 31297
rect 18144 31288 18196 31340
rect 17592 31220 17644 31272
rect 20996 31288 21048 31340
rect 21824 31331 21876 31340
rect 21824 31297 21833 31331
rect 21833 31297 21867 31331
rect 21867 31297 21876 31331
rect 21824 31288 21876 31297
rect 21916 31288 21968 31340
rect 21640 31152 21692 31204
rect 22192 31331 22244 31340
rect 22192 31297 22201 31331
rect 22201 31297 22235 31331
rect 22235 31297 22244 31331
rect 22192 31288 22244 31297
rect 22284 31220 22336 31272
rect 22836 31399 22888 31408
rect 22836 31365 22845 31399
rect 22845 31365 22879 31399
rect 22879 31365 22888 31399
rect 22836 31356 22888 31365
rect 24952 31424 25004 31476
rect 25044 31467 25096 31476
rect 25044 31433 25053 31467
rect 25053 31433 25087 31467
rect 25087 31433 25096 31467
rect 25044 31424 25096 31433
rect 28264 31424 28316 31476
rect 36636 31467 36688 31476
rect 36636 31433 36645 31467
rect 36645 31433 36679 31467
rect 36679 31433 36688 31467
rect 36636 31424 36688 31433
rect 26240 31356 26292 31408
rect 22560 31331 22612 31340
rect 22560 31297 22569 31331
rect 22569 31297 22603 31331
rect 22603 31297 22612 31331
rect 22560 31288 22612 31297
rect 24492 31331 24544 31340
rect 24492 31297 24501 31331
rect 24501 31297 24535 31331
rect 24535 31297 24544 31331
rect 24492 31288 24544 31297
rect 26424 31220 26476 31272
rect 26792 31263 26844 31272
rect 26792 31229 26801 31263
rect 26801 31229 26835 31263
rect 26835 31229 26844 31263
rect 26792 31220 26844 31229
rect 27620 31399 27672 31408
rect 27620 31365 27629 31399
rect 27629 31365 27663 31399
rect 27663 31365 27672 31399
rect 27620 31356 27672 31365
rect 28356 31356 28408 31408
rect 34612 31356 34664 31408
rect 36176 31356 36228 31408
rect 27344 31331 27396 31340
rect 27344 31297 27353 31331
rect 27353 31297 27387 31331
rect 27387 31297 27396 31331
rect 27344 31288 27396 31297
rect 32772 31331 32824 31340
rect 32772 31297 32781 31331
rect 32781 31297 32815 31331
rect 32815 31297 32824 31331
rect 32772 31288 32824 31297
rect 33140 31288 33192 31340
rect 33508 31288 33560 31340
rect 28356 31220 28408 31272
rect 31760 31220 31812 31272
rect 34428 31220 34480 31272
rect 26976 31152 27028 31204
rect 15752 31084 15804 31136
rect 16672 31084 16724 31136
rect 17408 31127 17460 31136
rect 17408 31093 17417 31127
rect 17417 31093 17451 31127
rect 17451 31093 17460 31127
rect 17408 31084 17460 31093
rect 24860 31084 24912 31136
rect 29920 31127 29972 31136
rect 29920 31093 29929 31127
rect 29929 31093 29963 31127
rect 29963 31093 29972 31127
rect 29920 31084 29972 31093
rect 30472 31127 30524 31136
rect 30472 31093 30481 31127
rect 30481 31093 30515 31127
rect 30515 31093 30524 31127
rect 30472 31084 30524 31093
rect 32588 31127 32640 31136
rect 32588 31093 32597 31127
rect 32597 31093 32631 31127
rect 32631 31093 32640 31127
rect 32588 31084 32640 31093
rect 33140 31084 33192 31136
rect 33416 31084 33468 31136
rect 35348 31084 35400 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3608 30880 3660 30932
rect 6736 30923 6788 30932
rect 6736 30889 6745 30923
rect 6745 30889 6779 30923
rect 6779 30889 6788 30923
rect 6736 30880 6788 30889
rect 7380 30880 7432 30932
rect 11796 30880 11848 30932
rect 4804 30812 4856 30864
rect 4068 30719 4120 30728
rect 4068 30685 4077 30719
rect 4077 30685 4111 30719
rect 4111 30685 4120 30719
rect 4068 30676 4120 30685
rect 5356 30744 5408 30796
rect 9496 30744 9548 30796
rect 11152 30744 11204 30796
rect 4620 30719 4672 30728
rect 4620 30685 4629 30719
rect 4629 30685 4663 30719
rect 4663 30685 4672 30719
rect 4620 30676 4672 30685
rect 4804 30676 4856 30728
rect 7196 30719 7248 30728
rect 7196 30685 7205 30719
rect 7205 30685 7239 30719
rect 7239 30685 7248 30719
rect 7196 30676 7248 30685
rect 7380 30719 7432 30728
rect 7380 30685 7389 30719
rect 7389 30685 7423 30719
rect 7423 30685 7432 30719
rect 7380 30676 7432 30685
rect 7656 30719 7708 30728
rect 7656 30685 7665 30719
rect 7665 30685 7699 30719
rect 7699 30685 7708 30719
rect 7656 30676 7708 30685
rect 12624 30719 12676 30728
rect 12624 30685 12633 30719
rect 12633 30685 12667 30719
rect 12667 30685 12676 30719
rect 12624 30676 12676 30685
rect 14096 30880 14148 30932
rect 16028 30880 16080 30932
rect 16120 30923 16172 30932
rect 16120 30889 16129 30923
rect 16129 30889 16163 30923
rect 16163 30889 16172 30923
rect 16120 30880 16172 30889
rect 16304 30880 16356 30932
rect 16948 30880 17000 30932
rect 23572 30923 23624 30932
rect 23572 30889 23581 30923
rect 23581 30889 23615 30923
rect 23615 30889 23624 30923
rect 23572 30880 23624 30889
rect 26976 30923 27028 30932
rect 26976 30889 26985 30923
rect 26985 30889 27019 30923
rect 27019 30889 27028 30923
rect 26976 30880 27028 30889
rect 31760 30880 31812 30932
rect 33324 30880 33376 30932
rect 33876 30880 33928 30932
rect 34244 30880 34296 30932
rect 14648 30787 14700 30796
rect 13636 30719 13688 30728
rect 13636 30685 13645 30719
rect 13645 30685 13679 30719
rect 13679 30685 13688 30719
rect 13636 30676 13688 30685
rect 5724 30608 5776 30660
rect 10140 30651 10192 30660
rect 10140 30617 10149 30651
rect 10149 30617 10183 30651
rect 10183 30617 10192 30651
rect 10140 30608 10192 30617
rect 10232 30608 10284 30660
rect 9036 30540 9088 30592
rect 9772 30540 9824 30592
rect 11704 30583 11756 30592
rect 11704 30549 11713 30583
rect 11713 30549 11747 30583
rect 11747 30549 11756 30583
rect 11704 30540 11756 30549
rect 13912 30651 13964 30660
rect 13912 30617 13921 30651
rect 13921 30617 13955 30651
rect 13955 30617 13964 30651
rect 13912 30608 13964 30617
rect 14004 30608 14056 30660
rect 14648 30753 14657 30787
rect 14657 30753 14691 30787
rect 14691 30753 14700 30787
rect 14648 30744 14700 30753
rect 15200 30787 15252 30796
rect 15200 30753 15209 30787
rect 15209 30753 15243 30787
rect 15243 30753 15252 30787
rect 15200 30744 15252 30753
rect 16212 30812 16264 30864
rect 17224 30812 17276 30864
rect 17684 30812 17736 30864
rect 22100 30812 22152 30864
rect 14556 30719 14608 30728
rect 14556 30685 14565 30719
rect 14565 30685 14599 30719
rect 14599 30685 14608 30719
rect 14556 30676 14608 30685
rect 15016 30676 15068 30728
rect 15752 30719 15804 30728
rect 15752 30685 15761 30719
rect 15761 30685 15795 30719
rect 15795 30685 15804 30719
rect 15752 30676 15804 30685
rect 20996 30744 21048 30796
rect 18144 30719 18196 30728
rect 18144 30685 18153 30719
rect 18153 30685 18187 30719
rect 18187 30685 18196 30719
rect 18144 30676 18196 30685
rect 23756 30719 23808 30728
rect 23756 30685 23765 30719
rect 23765 30685 23799 30719
rect 23799 30685 23808 30719
rect 23756 30676 23808 30685
rect 23848 30719 23900 30728
rect 23848 30685 23857 30719
rect 23857 30685 23891 30719
rect 23891 30685 23900 30719
rect 23848 30676 23900 30685
rect 24860 30812 24912 30864
rect 15292 30651 15344 30660
rect 15292 30617 15326 30651
rect 15326 30617 15344 30651
rect 15292 30608 15344 30617
rect 14096 30540 14148 30592
rect 15752 30540 15804 30592
rect 16304 30651 16356 30660
rect 16304 30617 16313 30651
rect 16313 30617 16347 30651
rect 16347 30617 16356 30651
rect 16304 30608 16356 30617
rect 16396 30608 16448 30660
rect 16580 30608 16632 30660
rect 17316 30540 17368 30592
rect 17868 30651 17920 30660
rect 17868 30617 17877 30651
rect 17877 30617 17911 30651
rect 17911 30617 17920 30651
rect 17868 30608 17920 30617
rect 18788 30608 18840 30660
rect 21364 30651 21416 30660
rect 21364 30617 21398 30651
rect 21398 30617 21416 30651
rect 21364 30608 21416 30617
rect 22744 30651 22796 30660
rect 22744 30617 22753 30651
rect 22753 30617 22787 30651
rect 22787 30617 22796 30651
rect 22744 30608 22796 30617
rect 22284 30540 22336 30592
rect 22652 30540 22704 30592
rect 23480 30540 23532 30592
rect 24400 30744 24452 30796
rect 25228 30744 25280 30796
rect 32772 30812 32824 30864
rect 25412 30719 25464 30728
rect 25412 30685 25421 30719
rect 25421 30685 25455 30719
rect 25455 30685 25464 30719
rect 25412 30676 25464 30685
rect 25596 30719 25648 30728
rect 25596 30685 25605 30719
rect 25605 30685 25639 30719
rect 25639 30685 25648 30719
rect 25596 30676 25648 30685
rect 30288 30744 30340 30796
rect 25964 30719 26016 30728
rect 25964 30685 25973 30719
rect 25973 30685 26007 30719
rect 26007 30685 26016 30719
rect 25964 30676 26016 30685
rect 32312 30719 32364 30728
rect 32312 30685 32321 30719
rect 32321 30685 32355 30719
rect 32355 30685 32364 30719
rect 32312 30676 32364 30685
rect 24492 30608 24544 30660
rect 24584 30651 24636 30660
rect 24584 30617 24593 30651
rect 24593 30617 24627 30651
rect 24627 30617 24636 30651
rect 24584 30608 24636 30617
rect 25228 30608 25280 30660
rect 26056 30608 26108 30660
rect 29920 30651 29972 30660
rect 29920 30617 29929 30651
rect 29929 30617 29963 30651
rect 29963 30617 29972 30651
rect 29920 30608 29972 30617
rect 31852 30608 31904 30660
rect 32128 30651 32180 30660
rect 32128 30617 32137 30651
rect 32137 30617 32171 30651
rect 32171 30617 32180 30651
rect 32128 30608 32180 30617
rect 32864 30719 32916 30728
rect 32864 30685 32873 30719
rect 32873 30685 32907 30719
rect 32907 30685 32916 30719
rect 32864 30676 32916 30685
rect 33508 30787 33560 30796
rect 33508 30753 33517 30787
rect 33517 30753 33551 30787
rect 33551 30753 33560 30787
rect 33508 30744 33560 30753
rect 33968 30744 34020 30796
rect 34428 30744 34480 30796
rect 33140 30719 33192 30728
rect 33140 30685 33149 30719
rect 33149 30685 33183 30719
rect 33183 30685 33192 30719
rect 33140 30676 33192 30685
rect 33232 30676 33284 30728
rect 24860 30583 24912 30592
rect 24860 30549 24869 30583
rect 24869 30549 24903 30583
rect 24903 30549 24912 30583
rect 24860 30540 24912 30549
rect 33692 30719 33744 30728
rect 33692 30685 33701 30719
rect 33701 30685 33735 30719
rect 33735 30685 33744 30719
rect 34244 30719 34296 30728
rect 33692 30676 33744 30685
rect 34244 30685 34253 30719
rect 34253 30685 34287 30719
rect 34287 30685 34296 30719
rect 34244 30676 34296 30685
rect 35992 30744 36044 30796
rect 35348 30719 35400 30728
rect 35348 30685 35357 30719
rect 35357 30685 35391 30719
rect 35391 30685 35400 30719
rect 35348 30676 35400 30685
rect 38476 30719 38528 30728
rect 38476 30685 38485 30719
rect 38485 30685 38519 30719
rect 38519 30685 38528 30719
rect 38476 30676 38528 30685
rect 33968 30583 34020 30592
rect 33968 30549 33990 30583
rect 33990 30549 34020 30583
rect 33968 30540 34020 30549
rect 34520 30583 34572 30592
rect 34520 30549 34529 30583
rect 34529 30549 34563 30583
rect 34563 30549 34572 30583
rect 34520 30540 34572 30549
rect 35072 30583 35124 30592
rect 35072 30549 35081 30583
rect 35081 30549 35115 30583
rect 35115 30549 35124 30583
rect 35072 30540 35124 30549
rect 36084 30608 36136 30660
rect 37188 30540 37240 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 4068 30336 4120 30388
rect 7380 30336 7432 30388
rect 14648 30336 14700 30388
rect 16212 30336 16264 30388
rect 8024 30268 8076 30320
rect 9036 30311 9088 30320
rect 9036 30277 9045 30311
rect 9045 30277 9079 30311
rect 9079 30277 9088 30311
rect 9036 30268 9088 30277
rect 3792 30200 3844 30252
rect 5448 30200 5500 30252
rect 5816 30200 5868 30252
rect 6828 30243 6880 30252
rect 6828 30209 6837 30243
rect 6837 30209 6871 30243
rect 6871 30209 6880 30243
rect 6828 30200 6880 30209
rect 9496 30200 9548 30252
rect 11152 30268 11204 30320
rect 13360 30268 13412 30320
rect 13912 30268 13964 30320
rect 14556 30268 14608 30320
rect 10416 30200 10468 30252
rect 10876 30175 10928 30184
rect 10876 30141 10885 30175
rect 10885 30141 10919 30175
rect 10919 30141 10928 30175
rect 10876 30132 10928 30141
rect 11704 30200 11756 30252
rect 12348 30243 12400 30252
rect 12348 30209 12357 30243
rect 12357 30209 12391 30243
rect 12391 30209 12400 30243
rect 12348 30200 12400 30209
rect 14096 30200 14148 30252
rect 16028 30243 16080 30252
rect 16028 30209 16037 30243
rect 16037 30209 16071 30243
rect 16071 30209 16080 30243
rect 16028 30200 16080 30209
rect 848 30064 900 30116
rect 3884 30107 3936 30116
rect 3884 30073 3893 30107
rect 3893 30073 3927 30107
rect 3927 30073 3936 30107
rect 3884 30064 3936 30073
rect 7104 30064 7156 30116
rect 11244 30064 11296 30116
rect 9220 29996 9272 30048
rect 14648 30175 14700 30184
rect 14648 30141 14657 30175
rect 14657 30141 14691 30175
rect 14691 30141 14700 30175
rect 14648 30132 14700 30141
rect 14832 30132 14884 30184
rect 15292 30132 15344 30184
rect 17408 30336 17460 30388
rect 17868 30336 17920 30388
rect 19340 30200 19392 30252
rect 19432 30243 19484 30252
rect 19432 30209 19441 30243
rect 19441 30209 19475 30243
rect 19475 30209 19484 30243
rect 19432 30200 19484 30209
rect 21364 30336 21416 30388
rect 19984 30200 20036 30252
rect 20352 30243 20404 30252
rect 20352 30209 20361 30243
rect 20361 30209 20395 30243
rect 20395 30209 20404 30243
rect 20352 30200 20404 30209
rect 21088 30200 21140 30252
rect 16672 30175 16724 30184
rect 15016 30064 15068 30116
rect 16672 30141 16681 30175
rect 16681 30141 16715 30175
rect 16715 30141 16724 30175
rect 16672 30132 16724 30141
rect 22100 30311 22152 30320
rect 22100 30277 22109 30311
rect 22109 30277 22143 30311
rect 22143 30277 22152 30311
rect 22100 30268 22152 30277
rect 26240 30268 26292 30320
rect 29276 30268 29328 30320
rect 21732 30200 21784 30252
rect 21916 30200 21968 30252
rect 21640 30175 21692 30184
rect 21640 30141 21649 30175
rect 21649 30141 21683 30175
rect 21683 30141 21692 30175
rect 21640 30132 21692 30141
rect 22100 30132 22152 30184
rect 23480 30243 23532 30252
rect 23480 30209 23489 30243
rect 23489 30209 23523 30243
rect 23523 30209 23532 30243
rect 23480 30200 23532 30209
rect 23848 30243 23900 30252
rect 23848 30209 23857 30243
rect 23857 30209 23891 30243
rect 23891 30209 23900 30243
rect 23848 30200 23900 30209
rect 24032 30243 24084 30252
rect 24032 30209 24041 30243
rect 24041 30209 24075 30243
rect 24075 30209 24084 30243
rect 24032 30200 24084 30209
rect 24124 30243 24176 30252
rect 24124 30209 24133 30243
rect 24133 30209 24167 30243
rect 24167 30209 24176 30243
rect 24124 30200 24176 30209
rect 29644 30243 29696 30252
rect 29644 30209 29653 30243
rect 29653 30209 29687 30243
rect 29687 30209 29696 30243
rect 29644 30200 29696 30209
rect 30288 30268 30340 30320
rect 30472 30268 30524 30320
rect 31852 30336 31904 30388
rect 34244 30336 34296 30388
rect 30840 30268 30892 30320
rect 32128 30200 32180 30252
rect 32588 30200 32640 30252
rect 33324 30268 33376 30320
rect 34520 30311 34572 30320
rect 34520 30277 34529 30311
rect 34529 30277 34563 30311
rect 34563 30277 34572 30311
rect 34520 30268 34572 30277
rect 35072 30336 35124 30388
rect 32956 30243 33008 30252
rect 32956 30209 32965 30243
rect 32965 30209 32999 30243
rect 32999 30209 33008 30243
rect 32956 30200 33008 30209
rect 33876 30200 33928 30252
rect 34704 30200 34756 30252
rect 35348 30200 35400 30252
rect 35440 30200 35492 30252
rect 36636 30200 36688 30252
rect 23664 30175 23716 30184
rect 23664 30141 23673 30175
rect 23673 30141 23707 30175
rect 23707 30141 23716 30175
rect 23664 30132 23716 30141
rect 24860 30132 24912 30184
rect 26056 30132 26108 30184
rect 26976 30175 27028 30184
rect 26976 30141 26985 30175
rect 26985 30141 27019 30175
rect 27019 30141 27028 30175
rect 26976 30132 27028 30141
rect 34428 30132 34480 30184
rect 35992 30132 36044 30184
rect 37188 30132 37240 30184
rect 22560 30064 22612 30116
rect 24124 30064 24176 30116
rect 32312 30064 32364 30116
rect 34612 30064 34664 30116
rect 12624 29996 12676 30048
rect 17040 30039 17092 30048
rect 17040 30005 17049 30039
rect 17049 30005 17083 30039
rect 17083 30005 17092 30039
rect 17040 29996 17092 30005
rect 19156 29996 19208 30048
rect 20536 30039 20588 30048
rect 20536 30005 20545 30039
rect 20545 30005 20579 30039
rect 20579 30005 20588 30039
rect 20536 29996 20588 30005
rect 20812 29996 20864 30048
rect 24584 29996 24636 30048
rect 24952 29996 25004 30048
rect 25412 29996 25464 30048
rect 25964 30039 26016 30048
rect 25964 30005 25973 30039
rect 25973 30005 26007 30039
rect 26007 30005 26016 30039
rect 25964 29996 26016 30005
rect 27528 29996 27580 30048
rect 29920 30039 29972 30048
rect 29920 30005 29929 30039
rect 29929 30005 29963 30039
rect 29963 30005 29972 30039
rect 29920 29996 29972 30005
rect 37464 29996 37516 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 13360 29792 13412 29844
rect 14648 29792 14700 29844
rect 17224 29835 17276 29844
rect 17224 29801 17233 29835
rect 17233 29801 17267 29835
rect 17267 29801 17276 29835
rect 17224 29792 17276 29801
rect 17316 29835 17368 29844
rect 17316 29801 17325 29835
rect 17325 29801 17359 29835
rect 17359 29801 17368 29835
rect 17316 29792 17368 29801
rect 17408 29792 17460 29844
rect 19432 29792 19484 29844
rect 18328 29724 18380 29776
rect 22744 29792 22796 29844
rect 24032 29792 24084 29844
rect 26976 29792 27028 29844
rect 28908 29792 28960 29844
rect 30564 29792 30616 29844
rect 23664 29724 23716 29776
rect 24768 29724 24820 29776
rect 26056 29767 26108 29776
rect 26056 29733 26065 29767
rect 26065 29733 26099 29767
rect 26099 29733 26108 29767
rect 26056 29724 26108 29733
rect 28540 29767 28592 29776
rect 28540 29733 28549 29767
rect 28549 29733 28583 29767
rect 28583 29733 28592 29767
rect 28540 29724 28592 29733
rect 4712 29656 4764 29708
rect 5264 29656 5316 29708
rect 848 29588 900 29640
rect 3332 29588 3384 29640
rect 6184 29588 6236 29640
rect 9220 29699 9272 29708
rect 9220 29665 9229 29699
rect 9229 29665 9263 29699
rect 9263 29665 9272 29699
rect 9220 29656 9272 29665
rect 10416 29656 10468 29708
rect 15016 29699 15068 29708
rect 15016 29665 15025 29699
rect 15025 29665 15059 29699
rect 15059 29665 15068 29699
rect 15016 29656 15068 29665
rect 15752 29699 15804 29708
rect 15752 29665 15761 29699
rect 15761 29665 15795 29699
rect 15795 29665 15804 29699
rect 15752 29656 15804 29665
rect 23848 29656 23900 29708
rect 24584 29656 24636 29708
rect 7472 29588 7524 29640
rect 7656 29588 7708 29640
rect 8116 29588 8168 29640
rect 8944 29631 8996 29640
rect 8944 29597 8953 29631
rect 8953 29597 8987 29631
rect 8987 29597 8996 29631
rect 8944 29588 8996 29597
rect 11152 29588 11204 29640
rect 12624 29588 12676 29640
rect 15200 29588 15252 29640
rect 17224 29588 17276 29640
rect 3884 29520 3936 29572
rect 6368 29563 6420 29572
rect 6368 29529 6377 29563
rect 6377 29529 6411 29563
rect 6411 29529 6420 29563
rect 6368 29520 6420 29529
rect 6828 29520 6880 29572
rect 10232 29520 10284 29572
rect 11520 29520 11572 29572
rect 17500 29563 17552 29572
rect 3424 29495 3476 29504
rect 3424 29461 3433 29495
rect 3433 29461 3467 29495
rect 3467 29461 3476 29495
rect 3424 29452 3476 29461
rect 4252 29452 4304 29504
rect 7380 29495 7432 29504
rect 7380 29461 7389 29495
rect 7389 29461 7423 29495
rect 7423 29461 7432 29495
rect 7380 29452 7432 29461
rect 9404 29452 9456 29504
rect 10876 29452 10928 29504
rect 11428 29452 11480 29504
rect 15108 29452 15160 29504
rect 17500 29529 17527 29563
rect 17527 29529 17552 29563
rect 17500 29520 17552 29529
rect 18788 29631 18840 29640
rect 18788 29597 18797 29631
rect 18797 29597 18831 29631
rect 18831 29597 18840 29631
rect 18788 29588 18840 29597
rect 19248 29588 19300 29640
rect 19708 29563 19760 29572
rect 19708 29529 19717 29563
rect 19717 29529 19751 29563
rect 19751 29529 19760 29563
rect 19708 29520 19760 29529
rect 19892 29631 19944 29640
rect 19892 29597 19901 29631
rect 19901 29597 19935 29631
rect 19935 29597 19944 29631
rect 19892 29588 19944 29597
rect 20536 29588 20588 29640
rect 22560 29588 22612 29640
rect 20260 29520 20312 29572
rect 17868 29452 17920 29504
rect 20812 29452 20864 29504
rect 22468 29520 22520 29572
rect 23296 29563 23348 29572
rect 23296 29529 23305 29563
rect 23305 29529 23339 29563
rect 23339 29529 23348 29563
rect 23296 29520 23348 29529
rect 24124 29588 24176 29640
rect 25228 29631 25280 29640
rect 25228 29597 25237 29631
rect 25237 29597 25271 29631
rect 25271 29597 25280 29631
rect 25228 29588 25280 29597
rect 25964 29656 26016 29708
rect 27528 29699 27580 29708
rect 27528 29665 27537 29699
rect 27537 29665 27571 29699
rect 27571 29665 27580 29699
rect 27528 29656 27580 29665
rect 30288 29724 30340 29776
rect 28908 29699 28960 29708
rect 28908 29665 28917 29699
rect 28917 29665 28951 29699
rect 28951 29665 28960 29699
rect 28908 29656 28960 29665
rect 23112 29495 23164 29504
rect 23112 29461 23121 29495
rect 23121 29461 23155 29495
rect 23155 29461 23164 29495
rect 24032 29520 24084 29572
rect 24492 29520 24544 29572
rect 24768 29520 24820 29572
rect 25780 29631 25832 29640
rect 25780 29597 25789 29631
rect 25789 29597 25823 29631
rect 25823 29597 25832 29631
rect 25780 29588 25832 29597
rect 29736 29656 29788 29708
rect 32956 29792 33008 29844
rect 33508 29792 33560 29844
rect 34336 29835 34388 29844
rect 34336 29801 34345 29835
rect 34345 29801 34379 29835
rect 34379 29801 34388 29835
rect 34336 29792 34388 29801
rect 35440 29792 35492 29844
rect 37280 29724 37332 29776
rect 29828 29588 29880 29640
rect 35348 29656 35400 29708
rect 26240 29520 26292 29572
rect 32128 29588 32180 29640
rect 33048 29631 33100 29640
rect 33048 29597 33057 29631
rect 33057 29597 33091 29631
rect 33091 29597 33100 29631
rect 33048 29588 33100 29597
rect 33232 29631 33284 29640
rect 33232 29597 33241 29631
rect 33241 29597 33275 29631
rect 33275 29597 33284 29631
rect 33232 29588 33284 29597
rect 33692 29588 33744 29640
rect 33876 29588 33928 29640
rect 36084 29588 36136 29640
rect 36728 29631 36780 29640
rect 36728 29597 36737 29631
rect 36737 29597 36771 29631
rect 36771 29597 36780 29631
rect 36728 29588 36780 29597
rect 36820 29588 36872 29640
rect 23112 29452 23164 29461
rect 24400 29452 24452 29504
rect 24860 29452 24912 29504
rect 30380 29452 30432 29504
rect 30472 29495 30524 29504
rect 30472 29461 30481 29495
rect 30481 29461 30515 29495
rect 30515 29461 30524 29495
rect 30472 29452 30524 29461
rect 31116 29495 31168 29504
rect 31116 29461 31143 29495
rect 31143 29461 31168 29495
rect 31116 29452 31168 29461
rect 31852 29520 31904 29572
rect 34152 29452 34204 29504
rect 34336 29495 34388 29504
rect 34336 29461 34345 29495
rect 34345 29461 34379 29495
rect 34379 29461 34388 29495
rect 34336 29452 34388 29461
rect 36452 29495 36504 29504
rect 36452 29461 36461 29495
rect 36461 29461 36495 29495
rect 36495 29461 36504 29495
rect 36452 29452 36504 29461
rect 37188 29452 37240 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 3424 29180 3476 29232
rect 4068 29155 4120 29164
rect 4068 29121 4077 29155
rect 4077 29121 4111 29155
rect 4111 29121 4120 29155
rect 4068 29112 4120 29121
rect 4252 29155 4304 29164
rect 4252 29121 4261 29155
rect 4261 29121 4295 29155
rect 4295 29121 4304 29155
rect 4252 29112 4304 29121
rect 4804 29180 4856 29232
rect 8024 29248 8076 29300
rect 7380 29180 7432 29232
rect 10232 29248 10284 29300
rect 11520 29291 11572 29300
rect 11520 29257 11529 29291
rect 11529 29257 11563 29291
rect 11563 29257 11572 29291
rect 11520 29248 11572 29257
rect 12624 29291 12676 29300
rect 12624 29257 12633 29291
rect 12633 29257 12667 29291
rect 12667 29257 12676 29291
rect 12624 29248 12676 29257
rect 14832 29291 14884 29300
rect 14832 29257 14841 29291
rect 14841 29257 14875 29291
rect 14875 29257 14884 29291
rect 14832 29248 14884 29257
rect 19248 29248 19300 29300
rect 10876 29180 10928 29232
rect 5816 29112 5868 29164
rect 6828 29155 6880 29164
rect 6828 29121 6837 29155
rect 6837 29121 6871 29155
rect 6871 29121 6880 29155
rect 6828 29112 6880 29121
rect 848 29044 900 29096
rect 3332 29044 3384 29096
rect 3700 29087 3752 29096
rect 3700 29053 3709 29087
rect 3709 29053 3743 29087
rect 3743 29053 3752 29087
rect 3700 29044 3752 29053
rect 4712 29087 4764 29096
rect 4712 29053 4721 29087
rect 4721 29053 4755 29087
rect 4755 29053 4764 29087
rect 4712 29044 4764 29053
rect 4804 29044 4856 29096
rect 7104 29044 7156 29096
rect 9404 29155 9456 29164
rect 9404 29121 9413 29155
rect 9413 29121 9447 29155
rect 9447 29121 9456 29155
rect 9404 29112 9456 29121
rect 13360 29180 13412 29232
rect 18328 29223 18380 29232
rect 18328 29189 18337 29223
rect 18337 29189 18371 29223
rect 18371 29189 18380 29223
rect 18328 29180 18380 29189
rect 12900 29112 12952 29164
rect 19340 29180 19392 29232
rect 20260 29291 20312 29300
rect 20260 29257 20269 29291
rect 20269 29257 20303 29291
rect 20303 29257 20312 29291
rect 20260 29248 20312 29257
rect 20352 29291 20404 29300
rect 20352 29257 20361 29291
rect 20361 29257 20395 29291
rect 20395 29257 20404 29291
rect 20352 29248 20404 29257
rect 20720 29248 20772 29300
rect 21088 29291 21140 29300
rect 21088 29257 21097 29291
rect 21097 29257 21131 29291
rect 21131 29257 21140 29291
rect 21088 29248 21140 29257
rect 24308 29248 24360 29300
rect 24676 29248 24728 29300
rect 19156 29155 19208 29164
rect 19156 29121 19190 29155
rect 19190 29121 19208 29155
rect 8116 28976 8168 29028
rect 11244 29087 11296 29096
rect 11244 29053 11253 29087
rect 11253 29053 11287 29087
rect 11287 29053 11296 29087
rect 11244 29044 11296 29053
rect 2964 28908 3016 28960
rect 6184 28951 6236 28960
rect 6184 28917 6193 28951
rect 6193 28917 6227 28951
rect 6227 28917 6236 28951
rect 6184 28908 6236 28917
rect 10508 28951 10560 28960
rect 10508 28917 10517 28951
rect 10517 28917 10551 28951
rect 10551 28917 10560 28951
rect 10508 28908 10560 28917
rect 12624 29044 12676 29096
rect 14004 29044 14056 29096
rect 19156 29112 19208 29121
rect 19708 29112 19760 29164
rect 20812 29180 20864 29232
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 20904 29112 20956 29121
rect 21180 29155 21232 29164
rect 21180 29121 21189 29155
rect 21189 29121 21223 29155
rect 21223 29121 21232 29155
rect 21180 29112 21232 29121
rect 21916 29180 21968 29232
rect 23112 29180 23164 29232
rect 23480 29180 23532 29232
rect 24032 29180 24084 29232
rect 26424 29248 26476 29300
rect 26516 29291 26568 29300
rect 26516 29257 26525 29291
rect 26525 29257 26559 29291
rect 26559 29257 26568 29291
rect 26516 29248 26568 29257
rect 29828 29248 29880 29300
rect 30012 29248 30064 29300
rect 30840 29248 30892 29300
rect 28540 29180 28592 29232
rect 29276 29180 29328 29232
rect 30380 29180 30432 29232
rect 32864 29248 32916 29300
rect 33876 29291 33928 29300
rect 33876 29257 33885 29291
rect 33885 29257 33919 29291
rect 33919 29257 33928 29291
rect 33876 29248 33928 29257
rect 34336 29248 34388 29300
rect 36636 29248 36688 29300
rect 33140 29180 33192 29232
rect 21640 29112 21692 29164
rect 15200 28976 15252 29028
rect 18144 29019 18196 29028
rect 18144 28985 18153 29019
rect 18153 28985 18187 29019
rect 18187 28985 18196 29019
rect 18144 28976 18196 28985
rect 21180 28976 21232 29028
rect 21640 28976 21692 29028
rect 22100 29044 22152 29096
rect 22008 28976 22060 29028
rect 23572 29155 23624 29164
rect 23572 29121 23581 29155
rect 23581 29121 23615 29155
rect 23615 29121 23624 29155
rect 23572 29112 23624 29121
rect 26792 29112 26844 29164
rect 30196 29155 30248 29164
rect 30196 29121 30205 29155
rect 30205 29121 30239 29155
rect 30239 29121 30248 29155
rect 30196 29112 30248 29121
rect 32772 29155 32824 29164
rect 32772 29121 32781 29155
rect 32781 29121 32815 29155
rect 32815 29121 32824 29155
rect 33600 29180 33652 29232
rect 34152 29180 34204 29232
rect 35992 29180 36044 29232
rect 32772 29112 32824 29121
rect 22468 29019 22520 29028
rect 22468 28985 22477 29019
rect 22477 28985 22511 29019
rect 22511 28985 22520 29019
rect 22468 28976 22520 28985
rect 25228 29044 25280 29096
rect 25596 29087 25648 29096
rect 25596 29053 25605 29087
rect 25605 29053 25639 29087
rect 25639 29053 25648 29087
rect 25596 29044 25648 29053
rect 26332 29087 26384 29096
rect 26332 29053 26341 29087
rect 26341 29053 26375 29087
rect 26375 29053 26384 29087
rect 26332 29044 26384 29053
rect 24124 28976 24176 29028
rect 25780 28976 25832 29028
rect 27620 29044 27672 29096
rect 31484 29044 31536 29096
rect 33048 29044 33100 29096
rect 34428 29112 34480 29164
rect 34612 29155 34664 29164
rect 34612 29121 34621 29155
rect 34621 29121 34655 29155
rect 34655 29121 34664 29155
rect 34612 29112 34664 29121
rect 36636 29155 36688 29164
rect 36636 29121 36645 29155
rect 36645 29121 36679 29155
rect 36679 29121 36688 29155
rect 36636 29112 36688 29121
rect 37188 29112 37240 29164
rect 34060 29087 34112 29096
rect 34060 29053 34069 29087
rect 34069 29053 34103 29087
rect 34103 29053 34112 29087
rect 34060 29044 34112 29053
rect 35440 29087 35492 29096
rect 35440 29053 35449 29087
rect 35449 29053 35483 29087
rect 35483 29053 35492 29087
rect 35440 29044 35492 29053
rect 26240 28908 26292 28960
rect 31852 28908 31904 28960
rect 33140 28908 33192 28960
rect 34060 28908 34112 28960
rect 34336 28976 34388 29028
rect 34796 28908 34848 28960
rect 36820 28951 36872 28960
rect 36820 28917 36829 28951
rect 36829 28917 36863 28951
rect 36863 28917 36872 28951
rect 36820 28908 36872 28917
rect 37004 28951 37056 28960
rect 37004 28917 37013 28951
rect 37013 28917 37047 28951
rect 37047 28917 37056 28951
rect 37004 28908 37056 28917
rect 37648 28908 37700 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3700 28704 3752 28756
rect 4068 28636 4120 28688
rect 7472 28704 7524 28756
rect 2964 28543 3016 28552
rect 2964 28509 2973 28543
rect 2973 28509 3007 28543
rect 3007 28509 3016 28543
rect 2964 28500 3016 28509
rect 3332 28543 3384 28552
rect 3332 28509 3341 28543
rect 3341 28509 3375 28543
rect 3375 28509 3384 28543
rect 3332 28500 3384 28509
rect 3608 28500 3660 28552
rect 3792 28543 3844 28552
rect 3792 28509 3801 28543
rect 3801 28509 3835 28543
rect 3835 28509 3844 28543
rect 3792 28500 3844 28509
rect 4068 28543 4120 28552
rect 4068 28509 4077 28543
rect 4077 28509 4111 28543
rect 4111 28509 4120 28543
rect 4068 28500 4120 28509
rect 4804 28611 4856 28620
rect 4804 28577 4813 28611
rect 4813 28577 4847 28611
rect 4847 28577 4856 28611
rect 4804 28568 4856 28577
rect 7012 28636 7064 28688
rect 8208 28704 8260 28756
rect 11244 28704 11296 28756
rect 12900 28747 12952 28756
rect 12900 28713 12909 28747
rect 12909 28713 12943 28747
rect 12943 28713 12952 28747
rect 12900 28704 12952 28713
rect 21916 28704 21968 28756
rect 25780 28704 25832 28756
rect 30012 28704 30064 28756
rect 6736 28568 6788 28620
rect 7380 28568 7432 28620
rect 8944 28568 8996 28620
rect 11428 28611 11480 28620
rect 11428 28577 11437 28611
rect 11437 28577 11471 28611
rect 11471 28577 11480 28611
rect 11428 28568 11480 28577
rect 13544 28568 13596 28620
rect 24676 28679 24728 28688
rect 24676 28645 24685 28679
rect 24685 28645 24719 28679
rect 24719 28645 24728 28679
rect 24676 28636 24728 28645
rect 15200 28611 15252 28620
rect 15200 28577 15209 28611
rect 15209 28577 15243 28611
rect 15243 28577 15252 28611
rect 15200 28568 15252 28577
rect 16028 28611 16080 28620
rect 16028 28577 16037 28611
rect 16037 28577 16071 28611
rect 16071 28577 16080 28611
rect 16028 28568 16080 28577
rect 16304 28568 16356 28620
rect 23572 28568 23624 28620
rect 23940 28611 23992 28620
rect 23940 28577 23949 28611
rect 23949 28577 23983 28611
rect 23983 28577 23992 28611
rect 23940 28568 23992 28577
rect 24216 28568 24268 28620
rect 4712 28543 4764 28552
rect 4712 28509 4721 28543
rect 4721 28509 4755 28543
rect 4755 28509 4764 28543
rect 4712 28500 4764 28509
rect 6920 28500 6972 28552
rect 8116 28500 8168 28552
rect 11152 28543 11204 28552
rect 11152 28509 11161 28543
rect 11161 28509 11195 28543
rect 11195 28509 11204 28543
rect 11152 28500 11204 28509
rect 13360 28500 13412 28552
rect 16948 28500 17000 28552
rect 21548 28500 21600 28552
rect 22376 28543 22428 28552
rect 22376 28509 22385 28543
rect 22385 28509 22419 28543
rect 22419 28509 22428 28543
rect 22376 28500 22428 28509
rect 5172 28432 5224 28484
rect 5816 28432 5868 28484
rect 5448 28364 5500 28416
rect 7472 28432 7524 28484
rect 8208 28475 8260 28484
rect 8208 28441 8217 28475
rect 8217 28441 8251 28475
rect 8251 28441 8260 28475
rect 8208 28432 8260 28441
rect 9588 28475 9640 28484
rect 9588 28441 9597 28475
rect 9597 28441 9631 28475
rect 9631 28441 9640 28475
rect 9588 28432 9640 28441
rect 10232 28432 10284 28484
rect 13452 28475 13504 28484
rect 13452 28441 13461 28475
rect 13461 28441 13495 28475
rect 13495 28441 13504 28475
rect 13452 28432 13504 28441
rect 6644 28407 6696 28416
rect 6644 28373 6653 28407
rect 6653 28373 6687 28407
rect 6687 28373 6696 28407
rect 6644 28364 6696 28373
rect 12992 28407 13044 28416
rect 12992 28373 13001 28407
rect 13001 28373 13035 28407
rect 13035 28373 13044 28407
rect 12992 28364 13044 28373
rect 13912 28364 13964 28416
rect 14188 28407 14240 28416
rect 14188 28373 14197 28407
rect 14197 28373 14231 28407
rect 14231 28373 14240 28407
rect 17592 28432 17644 28484
rect 17960 28432 18012 28484
rect 19064 28475 19116 28484
rect 19064 28441 19073 28475
rect 19073 28441 19107 28475
rect 19107 28441 19116 28475
rect 19064 28432 19116 28441
rect 22652 28543 22704 28552
rect 22652 28509 22661 28543
rect 22661 28509 22695 28543
rect 22695 28509 22704 28543
rect 22652 28500 22704 28509
rect 26516 28568 26568 28620
rect 30196 28636 30248 28688
rect 30472 28704 30524 28756
rect 31484 28704 31536 28756
rect 31668 28704 31720 28756
rect 34612 28704 34664 28756
rect 34888 28704 34940 28756
rect 26424 28500 26476 28552
rect 22928 28432 22980 28484
rect 24216 28432 24268 28484
rect 25596 28432 25648 28484
rect 28448 28543 28500 28552
rect 28448 28509 28457 28543
rect 28457 28509 28491 28543
rect 28491 28509 28500 28543
rect 28448 28500 28500 28509
rect 29000 28543 29052 28552
rect 29000 28509 29009 28543
rect 29009 28509 29043 28543
rect 29043 28509 29052 28543
rect 29000 28500 29052 28509
rect 29184 28500 29236 28552
rect 29736 28543 29788 28552
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 30012 28543 30064 28552
rect 30012 28509 30021 28543
rect 30021 28509 30055 28543
rect 30055 28509 30064 28543
rect 30012 28500 30064 28509
rect 30196 28543 30248 28552
rect 30196 28509 30205 28543
rect 30205 28509 30239 28543
rect 30239 28509 30248 28543
rect 31116 28568 31168 28620
rect 30196 28500 30248 28509
rect 14188 28364 14240 28373
rect 15476 28364 15528 28416
rect 15752 28407 15804 28416
rect 15752 28373 15761 28407
rect 15761 28373 15795 28407
rect 15795 28373 15804 28407
rect 15752 28364 15804 28373
rect 15844 28407 15896 28416
rect 15844 28373 15853 28407
rect 15853 28373 15887 28407
rect 15887 28373 15896 28407
rect 15844 28364 15896 28373
rect 22836 28364 22888 28416
rect 30748 28432 30800 28484
rect 27620 28364 27672 28416
rect 28264 28364 28316 28416
rect 29736 28364 29788 28416
rect 29828 28364 29880 28416
rect 31116 28475 31168 28484
rect 31116 28441 31125 28475
rect 31125 28441 31159 28475
rect 31159 28441 31168 28475
rect 33968 28636 34020 28688
rect 34060 28636 34112 28688
rect 35532 28636 35584 28688
rect 33508 28611 33560 28620
rect 33508 28577 33517 28611
rect 33517 28577 33551 28611
rect 33551 28577 33560 28611
rect 33508 28568 33560 28577
rect 34336 28568 34388 28620
rect 33140 28500 33192 28552
rect 31116 28432 31168 28441
rect 32772 28432 32824 28484
rect 33784 28543 33836 28552
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 33784 28500 33836 28509
rect 33968 28500 34020 28552
rect 34152 28500 34204 28552
rect 33048 28407 33100 28416
rect 33048 28373 33057 28407
rect 33057 28373 33091 28407
rect 33091 28373 33100 28407
rect 33048 28364 33100 28373
rect 33600 28432 33652 28484
rect 34336 28432 34388 28484
rect 34888 28568 34940 28620
rect 35348 28500 35400 28552
rect 35532 28543 35584 28552
rect 35532 28509 35541 28543
rect 35541 28509 35575 28543
rect 35575 28509 35584 28543
rect 35532 28500 35584 28509
rect 35992 28747 36044 28756
rect 35992 28713 36001 28747
rect 36001 28713 36035 28747
rect 36035 28713 36044 28747
rect 35992 28704 36044 28713
rect 36452 28611 36504 28620
rect 36452 28577 36461 28611
rect 36461 28577 36495 28611
rect 36495 28577 36504 28611
rect 36452 28568 36504 28577
rect 36820 28611 36872 28620
rect 36820 28577 36829 28611
rect 36829 28577 36863 28611
rect 36863 28577 36872 28611
rect 36820 28568 36872 28577
rect 36176 28543 36228 28552
rect 36176 28509 36185 28543
rect 36185 28509 36219 28543
rect 36219 28509 36228 28543
rect 36176 28500 36228 28509
rect 36360 28543 36412 28552
rect 36360 28509 36369 28543
rect 36369 28509 36403 28543
rect 36403 28509 36412 28543
rect 36360 28500 36412 28509
rect 37004 28543 37056 28552
rect 37004 28509 37013 28543
rect 37013 28509 37047 28543
rect 37047 28509 37056 28543
rect 37004 28500 37056 28509
rect 37464 28543 37516 28552
rect 37464 28509 37473 28543
rect 37473 28509 37507 28543
rect 37507 28509 37516 28543
rect 37464 28500 37516 28509
rect 37740 28543 37792 28552
rect 37740 28509 37749 28543
rect 37749 28509 37783 28543
rect 37783 28509 37792 28543
rect 37740 28500 37792 28509
rect 37924 28543 37976 28552
rect 37924 28509 37933 28543
rect 37933 28509 37967 28543
rect 37967 28509 37976 28543
rect 37924 28500 37976 28509
rect 33692 28364 33744 28416
rect 34796 28364 34848 28416
rect 37556 28432 37608 28484
rect 35348 28364 35400 28416
rect 35532 28364 35584 28416
rect 36176 28364 36228 28416
rect 38016 28364 38068 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 2780 28092 2832 28144
rect 3608 28092 3660 28144
rect 3976 28024 4028 28076
rect 1400 27956 1452 28008
rect 3424 27956 3476 28008
rect 4068 27956 4120 28008
rect 3148 27888 3200 27940
rect 4620 28024 4672 28076
rect 4712 28067 4764 28076
rect 4712 28033 4721 28067
rect 4721 28033 4755 28067
rect 4755 28033 4764 28067
rect 4712 28024 4764 28033
rect 5264 28092 5316 28144
rect 6644 28160 6696 28212
rect 7012 28135 7064 28144
rect 7012 28101 7021 28135
rect 7021 28101 7055 28135
rect 7055 28101 7064 28135
rect 7012 28092 7064 28101
rect 6736 28067 6788 28076
rect 6736 28033 6745 28067
rect 6745 28033 6779 28067
rect 6779 28033 6788 28067
rect 6736 28024 6788 28033
rect 7564 28160 7616 28212
rect 8852 28160 8904 28212
rect 9588 28160 9640 28212
rect 15292 28160 15344 28212
rect 15752 28160 15804 28212
rect 17592 28203 17644 28212
rect 17592 28169 17601 28203
rect 17601 28169 17635 28203
rect 17635 28169 17644 28203
rect 17592 28160 17644 28169
rect 10232 28092 10284 28144
rect 10416 28067 10468 28076
rect 10416 28033 10425 28067
rect 10425 28033 10459 28067
rect 10459 28033 10468 28067
rect 10416 28024 10468 28033
rect 10508 28024 10560 28076
rect 11152 28024 11204 28076
rect 12624 28092 12676 28144
rect 13636 28092 13688 28144
rect 15200 28092 15252 28144
rect 16488 28092 16540 28144
rect 19064 28160 19116 28212
rect 20904 28160 20956 28212
rect 21824 28160 21876 28212
rect 23940 28203 23992 28212
rect 23940 28169 23949 28203
rect 23949 28169 23983 28203
rect 23983 28169 23992 28203
rect 23940 28160 23992 28169
rect 28448 28160 28500 28212
rect 29736 28203 29788 28212
rect 29736 28169 29745 28203
rect 29745 28169 29779 28203
rect 29779 28169 29788 28203
rect 29736 28160 29788 28169
rect 30748 28160 30800 28212
rect 19340 28092 19392 28144
rect 20720 28092 20772 28144
rect 22008 28135 22060 28144
rect 22008 28101 22017 28135
rect 22017 28101 22051 28135
rect 22051 28101 22060 28135
rect 22008 28092 22060 28101
rect 24216 28092 24268 28144
rect 6920 27999 6972 28008
rect 6920 27965 6929 27999
rect 6929 27965 6963 27999
rect 6963 27965 6972 27999
rect 6920 27956 6972 27965
rect 7380 27956 7432 28008
rect 8208 27956 8260 28008
rect 12992 27956 13044 28008
rect 13820 27956 13872 28008
rect 2872 27820 2924 27872
rect 3792 27820 3844 27872
rect 5448 27863 5500 27872
rect 5448 27829 5457 27863
rect 5457 27829 5491 27863
rect 5491 27829 5500 27863
rect 5448 27820 5500 27829
rect 6184 27888 6236 27940
rect 6920 27820 6972 27872
rect 13912 27820 13964 27872
rect 15476 27999 15528 28008
rect 15476 27965 15485 27999
rect 15485 27965 15519 27999
rect 15519 27965 15528 27999
rect 15476 27956 15528 27965
rect 15936 28024 15988 28076
rect 17960 28024 18012 28076
rect 18880 28024 18932 28076
rect 19524 28067 19576 28076
rect 19524 28033 19533 28067
rect 19533 28033 19567 28067
rect 19567 28033 19576 28067
rect 19524 28024 19576 28033
rect 16028 27956 16080 28008
rect 18052 27999 18104 28008
rect 18052 27965 18061 27999
rect 18061 27965 18095 27999
rect 18095 27965 18104 27999
rect 18052 27956 18104 27965
rect 18144 27999 18196 28008
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 16856 27820 16908 27872
rect 19616 27820 19668 27872
rect 21272 28024 21324 28076
rect 22192 28067 22244 28076
rect 22192 28033 22201 28067
rect 22201 28033 22235 28067
rect 22235 28033 22244 28067
rect 22192 28024 22244 28033
rect 22560 28067 22612 28076
rect 22560 28033 22569 28067
rect 22569 28033 22603 28067
rect 22603 28033 22612 28067
rect 22560 28024 22612 28033
rect 22836 28067 22888 28076
rect 22836 28033 22870 28067
rect 22870 28033 22888 28067
rect 22836 28024 22888 28033
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 24400 28024 24452 28033
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 24860 28024 24912 28076
rect 24952 28067 25004 28076
rect 24952 28033 24961 28067
rect 24961 28033 24995 28067
rect 24995 28033 25004 28067
rect 24952 28024 25004 28033
rect 25228 28067 25280 28076
rect 25228 28033 25237 28067
rect 25237 28033 25271 28067
rect 25271 28033 25280 28067
rect 25228 28024 25280 28033
rect 26240 28092 26292 28144
rect 28264 28135 28316 28144
rect 28264 28101 28273 28135
rect 28273 28101 28307 28135
rect 28307 28101 28316 28135
rect 28264 28092 28316 28101
rect 29276 28092 29328 28144
rect 25688 28024 25740 28076
rect 27620 28024 27672 28076
rect 20720 27956 20772 28008
rect 21088 27999 21140 28008
rect 21088 27965 21097 27999
rect 21097 27965 21131 27999
rect 21131 27965 21140 27999
rect 21088 27956 21140 27965
rect 21180 27999 21232 28008
rect 21180 27965 21189 27999
rect 21189 27965 21223 27999
rect 21223 27965 21232 27999
rect 21180 27956 21232 27965
rect 24768 27999 24820 28008
rect 24768 27965 24777 27999
rect 24777 27965 24811 27999
rect 24811 27965 24820 27999
rect 24768 27956 24820 27965
rect 26240 27956 26292 28008
rect 26976 27999 27028 28008
rect 26976 27965 26985 27999
rect 26985 27965 27019 27999
rect 27019 27965 27028 27999
rect 26976 27956 27028 27965
rect 29920 28092 29972 28144
rect 31484 28092 31536 28144
rect 30748 28024 30800 28076
rect 31852 28160 31904 28212
rect 34796 28160 34848 28212
rect 36360 28160 36412 28212
rect 37740 28160 37792 28212
rect 32956 28092 33008 28144
rect 33692 28092 33744 28144
rect 34336 28067 34388 28076
rect 34336 28033 34345 28067
rect 34345 28033 34379 28067
rect 34379 28033 34388 28067
rect 34336 28024 34388 28033
rect 37556 28135 37608 28144
rect 37556 28101 37565 28135
rect 37565 28101 37599 28135
rect 37599 28101 37608 28135
rect 37556 28092 37608 28101
rect 37648 28135 37700 28144
rect 37648 28101 37657 28135
rect 37657 28101 37691 28135
rect 37691 28101 37700 28135
rect 37648 28092 37700 28101
rect 37280 28067 37332 28076
rect 37280 28033 37289 28067
rect 37289 28033 37323 28067
rect 37323 28033 37332 28067
rect 37280 28024 37332 28033
rect 30840 27956 30892 28008
rect 31116 27956 31168 28008
rect 26332 27888 26384 27940
rect 32772 27956 32824 28008
rect 33968 27999 34020 28008
rect 33968 27965 33977 27999
rect 33977 27965 34011 27999
rect 34011 27965 34020 27999
rect 33968 27956 34020 27965
rect 35440 27956 35492 28008
rect 20076 27863 20128 27872
rect 20076 27829 20085 27863
rect 20085 27829 20119 27863
rect 20119 27829 20128 27863
rect 20076 27820 20128 27829
rect 21548 27820 21600 27872
rect 27528 27820 27580 27872
rect 31484 27820 31536 27872
rect 32680 27820 32732 27872
rect 35256 27888 35308 27940
rect 37740 28067 37792 28076
rect 37740 28033 37754 28067
rect 37754 28033 37788 28067
rect 37788 28033 37792 28067
rect 37740 28024 37792 28033
rect 38016 28067 38068 28076
rect 38016 28033 38025 28067
rect 38025 28033 38059 28067
rect 38059 28033 38068 28067
rect 38016 28024 38068 28033
rect 38016 27888 38068 27940
rect 34520 27863 34572 27872
rect 34520 27829 34529 27863
rect 34529 27829 34563 27863
rect 34563 27829 34572 27863
rect 34520 27820 34572 27829
rect 38200 27863 38252 27872
rect 38200 27829 38209 27863
rect 38209 27829 38243 27863
rect 38243 27829 38252 27863
rect 38200 27820 38252 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3424 27659 3476 27668
rect 3424 27625 3433 27659
rect 3433 27625 3467 27659
rect 3467 27625 3476 27659
rect 3424 27616 3476 27625
rect 3608 27659 3660 27668
rect 3608 27625 3617 27659
rect 3617 27625 3651 27659
rect 3651 27625 3660 27659
rect 3608 27616 3660 27625
rect 3976 27659 4028 27668
rect 3976 27625 3985 27659
rect 3985 27625 4019 27659
rect 4019 27625 4028 27659
rect 3976 27616 4028 27625
rect 7564 27616 7616 27668
rect 7288 27548 7340 27600
rect 13912 27616 13964 27668
rect 14372 27659 14424 27668
rect 14372 27625 14381 27659
rect 14381 27625 14415 27659
rect 14415 27625 14424 27659
rect 14372 27616 14424 27625
rect 14556 27548 14608 27600
rect 15108 27591 15160 27600
rect 15108 27557 15117 27591
rect 15117 27557 15151 27591
rect 15151 27557 15160 27591
rect 16396 27616 16448 27668
rect 16856 27616 16908 27668
rect 17776 27616 17828 27668
rect 15108 27548 15160 27557
rect 17592 27548 17644 27600
rect 3332 27480 3384 27532
rect 13544 27523 13596 27532
rect 13544 27489 13553 27523
rect 13553 27489 13587 27523
rect 13587 27489 13596 27523
rect 13544 27480 13596 27489
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 2780 27412 2832 27464
rect 3056 27412 3108 27464
rect 3148 27412 3200 27464
rect 1676 27387 1728 27396
rect 1676 27353 1685 27387
rect 1685 27353 1719 27387
rect 1719 27353 1728 27387
rect 1676 27344 1728 27353
rect 3608 27412 3660 27464
rect 3332 27276 3384 27328
rect 4620 27412 4672 27464
rect 7012 27412 7064 27464
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 10232 27412 10284 27464
rect 15292 27480 15344 27532
rect 5264 27344 5316 27396
rect 12624 27344 12676 27396
rect 13636 27344 13688 27396
rect 5448 27319 5500 27328
rect 5448 27285 5457 27319
rect 5457 27285 5491 27319
rect 5491 27285 5500 27319
rect 5448 27276 5500 27285
rect 6368 27276 6420 27328
rect 13084 27276 13136 27328
rect 13452 27319 13504 27328
rect 13452 27285 13461 27319
rect 13461 27285 13495 27319
rect 13495 27285 13504 27319
rect 13452 27276 13504 27285
rect 14832 27319 14884 27328
rect 14832 27285 14841 27319
rect 14841 27285 14875 27319
rect 14875 27285 14884 27319
rect 14832 27276 14884 27285
rect 15200 27455 15252 27464
rect 15200 27421 15209 27455
rect 15209 27421 15243 27455
rect 15243 27421 15252 27455
rect 15660 27480 15712 27532
rect 15936 27480 15988 27532
rect 16948 27480 17000 27532
rect 18788 27616 18840 27668
rect 19524 27616 19576 27668
rect 19340 27548 19392 27600
rect 19432 27548 19484 27600
rect 19064 27480 19116 27532
rect 15200 27412 15252 27421
rect 16396 27344 16448 27396
rect 17684 27412 17736 27464
rect 17960 27344 18012 27396
rect 18972 27412 19024 27464
rect 19340 27455 19392 27464
rect 19340 27421 19349 27455
rect 19349 27421 19383 27455
rect 19383 27421 19392 27455
rect 19340 27412 19392 27421
rect 19524 27455 19576 27464
rect 19524 27421 19533 27455
rect 19533 27421 19567 27455
rect 19567 27421 19576 27455
rect 19524 27412 19576 27421
rect 21180 27548 21232 27600
rect 22836 27616 22888 27668
rect 27528 27616 27580 27668
rect 27712 27616 27764 27668
rect 28724 27616 28776 27668
rect 29828 27616 29880 27668
rect 31392 27616 31444 27668
rect 31760 27659 31812 27668
rect 31760 27625 31769 27659
rect 31769 27625 31803 27659
rect 31803 27625 31812 27659
rect 31760 27616 31812 27625
rect 33968 27616 34020 27668
rect 18696 27387 18748 27396
rect 18696 27353 18705 27387
rect 18705 27353 18739 27387
rect 18739 27353 18748 27387
rect 18696 27344 18748 27353
rect 18880 27387 18932 27396
rect 18880 27353 18889 27387
rect 18889 27353 18923 27387
rect 18923 27353 18932 27387
rect 18880 27344 18932 27353
rect 19432 27344 19484 27396
rect 16304 27276 16356 27328
rect 17868 27319 17920 27328
rect 17868 27285 17877 27319
rect 17877 27285 17911 27319
rect 17911 27285 17920 27319
rect 17868 27276 17920 27285
rect 18144 27319 18196 27328
rect 18144 27285 18153 27319
rect 18153 27285 18187 27319
rect 18187 27285 18196 27319
rect 18144 27276 18196 27285
rect 18420 27276 18472 27328
rect 20444 27412 20496 27464
rect 21548 27523 21600 27532
rect 21548 27489 21557 27523
rect 21557 27489 21591 27523
rect 21591 27489 21600 27523
rect 21548 27480 21600 27489
rect 21456 27455 21508 27464
rect 21456 27421 21465 27455
rect 21465 27421 21499 27455
rect 21499 27421 21508 27455
rect 21456 27412 21508 27421
rect 19708 27344 19760 27396
rect 19800 27276 19852 27328
rect 21088 27344 21140 27396
rect 21548 27344 21600 27396
rect 20628 27319 20680 27328
rect 20628 27285 20637 27319
rect 20637 27285 20671 27319
rect 20671 27285 20680 27319
rect 20628 27276 20680 27285
rect 21364 27276 21416 27328
rect 21824 27455 21876 27464
rect 21824 27421 21833 27455
rect 21833 27421 21867 27455
rect 21867 27421 21876 27455
rect 21824 27412 21876 27421
rect 22928 27412 22980 27464
rect 24768 27548 24820 27600
rect 26240 27548 26292 27600
rect 29000 27548 29052 27600
rect 24584 27480 24636 27532
rect 24032 27412 24084 27464
rect 25688 27480 25740 27532
rect 26976 27480 27028 27532
rect 27620 27523 27672 27532
rect 27620 27489 27629 27523
rect 27629 27489 27663 27523
rect 27663 27489 27672 27523
rect 27620 27480 27672 27489
rect 30840 27523 30892 27532
rect 30840 27489 30849 27523
rect 30849 27489 30883 27523
rect 30883 27489 30892 27523
rect 30840 27480 30892 27489
rect 31116 27523 31168 27532
rect 31116 27489 31125 27523
rect 31125 27489 31159 27523
rect 31159 27489 31168 27523
rect 31116 27480 31168 27489
rect 24308 27344 24360 27396
rect 22744 27276 22796 27328
rect 23296 27276 23348 27328
rect 24860 27344 24912 27396
rect 25872 27412 25924 27464
rect 30748 27455 30800 27464
rect 30748 27421 30757 27455
rect 30757 27421 30791 27455
rect 30791 27421 30800 27455
rect 30748 27412 30800 27421
rect 31484 27455 31536 27464
rect 31484 27421 31493 27455
rect 31493 27421 31527 27455
rect 31527 27421 31536 27455
rect 31484 27412 31536 27421
rect 32128 27591 32180 27600
rect 32128 27557 32137 27591
rect 32137 27557 32171 27591
rect 32171 27557 32180 27591
rect 32128 27548 32180 27557
rect 33140 27548 33192 27600
rect 35348 27548 35400 27600
rect 37740 27616 37792 27668
rect 37924 27616 37976 27668
rect 37556 27548 37608 27600
rect 31852 27523 31904 27532
rect 31852 27489 31861 27523
rect 31861 27489 31895 27523
rect 31895 27489 31904 27523
rect 31852 27480 31904 27489
rect 32772 27523 32824 27532
rect 32772 27489 32781 27523
rect 32781 27489 32815 27523
rect 32815 27489 32824 27523
rect 32772 27480 32824 27489
rect 33048 27455 33100 27464
rect 33048 27421 33057 27455
rect 33057 27421 33091 27455
rect 33091 27421 33100 27455
rect 33048 27412 33100 27421
rect 26884 27344 26936 27396
rect 28264 27344 28316 27396
rect 32404 27344 32456 27396
rect 35256 27412 35308 27464
rect 26424 27276 26476 27328
rect 27988 27319 28040 27328
rect 27988 27285 27997 27319
rect 27997 27285 28031 27319
rect 28031 27285 28040 27319
rect 27988 27276 28040 27285
rect 28172 27319 28224 27328
rect 28172 27285 28181 27319
rect 28181 27285 28215 27319
rect 28215 27285 28224 27319
rect 28172 27276 28224 27285
rect 28816 27319 28868 27328
rect 28816 27285 28843 27319
rect 28843 27285 28868 27319
rect 28816 27276 28868 27285
rect 29644 27276 29696 27328
rect 32956 27276 33008 27328
rect 34796 27276 34848 27328
rect 35348 27276 35400 27328
rect 37372 27412 37424 27464
rect 37464 27319 37516 27328
rect 37464 27285 37473 27319
rect 37473 27285 37507 27319
rect 37507 27285 37516 27319
rect 37464 27276 37516 27285
rect 37556 27276 37608 27328
rect 37924 27455 37976 27464
rect 37924 27421 37933 27455
rect 37933 27421 37967 27455
rect 37967 27421 37976 27455
rect 37924 27412 37976 27421
rect 38016 27455 38068 27464
rect 38016 27421 38025 27455
rect 38025 27421 38059 27455
rect 38059 27421 38068 27455
rect 38016 27412 38068 27421
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 3424 27072 3476 27124
rect 3976 27072 4028 27124
rect 6276 27004 6328 27056
rect 13452 27072 13504 27124
rect 17776 27072 17828 27124
rect 18420 27072 18472 27124
rect 19524 27072 19576 27124
rect 21364 27115 21416 27124
rect 21364 27081 21373 27115
rect 21373 27081 21407 27115
rect 21407 27081 21416 27115
rect 21364 27072 21416 27081
rect 21824 27072 21876 27124
rect 13268 27004 13320 27056
rect 3332 26979 3384 26988
rect 3332 26945 3341 26979
rect 3341 26945 3375 26979
rect 3375 26945 3384 26979
rect 3332 26936 3384 26945
rect 1676 26868 1728 26920
rect 3148 26868 3200 26920
rect 3976 26868 4028 26920
rect 5264 26911 5316 26920
rect 5264 26877 5273 26911
rect 5273 26877 5307 26911
rect 5307 26877 5316 26911
rect 6092 26936 6144 26988
rect 6368 26936 6420 26988
rect 13176 26936 13228 26988
rect 14004 26979 14056 26988
rect 14004 26945 14013 26979
rect 14013 26945 14047 26979
rect 14047 26945 14056 26979
rect 14004 26936 14056 26945
rect 5264 26868 5316 26877
rect 8300 26868 8352 26920
rect 5816 26732 5868 26784
rect 9404 26732 9456 26784
rect 9680 26911 9732 26920
rect 9680 26877 9689 26911
rect 9689 26877 9723 26911
rect 9723 26877 9732 26911
rect 9680 26868 9732 26877
rect 11152 26911 11204 26920
rect 11152 26877 11161 26911
rect 11161 26877 11195 26911
rect 11195 26877 11204 26911
rect 11152 26868 11204 26877
rect 13728 26868 13780 26920
rect 13452 26800 13504 26852
rect 14372 26936 14424 26988
rect 15292 26979 15344 26988
rect 15292 26945 15301 26979
rect 15301 26945 15335 26979
rect 15335 26945 15344 26979
rect 15292 26936 15344 26945
rect 15476 26979 15528 26988
rect 15476 26945 15485 26979
rect 15485 26945 15519 26979
rect 15519 26945 15528 26979
rect 15476 26936 15528 26945
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 17868 27004 17920 27056
rect 19340 27004 19392 27056
rect 22376 27004 22428 27056
rect 25872 27004 25924 27056
rect 17960 26936 18012 26988
rect 18052 26936 18104 26988
rect 14832 26868 14884 26920
rect 16212 26868 16264 26920
rect 19616 26979 19668 26988
rect 19616 26945 19625 26979
rect 19625 26945 19659 26979
rect 19659 26945 19668 26979
rect 19616 26936 19668 26945
rect 19800 26979 19852 26988
rect 19800 26945 19809 26979
rect 19809 26945 19843 26979
rect 19843 26945 19852 26979
rect 19800 26936 19852 26945
rect 19708 26868 19760 26920
rect 20076 26979 20128 26988
rect 20076 26945 20085 26979
rect 20085 26945 20119 26979
rect 20119 26945 20128 26979
rect 20076 26936 20128 26945
rect 21456 26979 21508 26988
rect 21456 26945 21465 26979
rect 21465 26945 21499 26979
rect 21499 26945 21508 26979
rect 21456 26936 21508 26945
rect 21548 26936 21600 26988
rect 21824 26979 21876 26988
rect 21824 26945 21833 26979
rect 21833 26945 21867 26979
rect 21867 26945 21876 26979
rect 21824 26936 21876 26945
rect 22744 26936 22796 26988
rect 23296 26979 23348 26988
rect 23296 26945 23305 26979
rect 23305 26945 23339 26979
rect 23339 26945 23348 26979
rect 23296 26936 23348 26945
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 25596 26936 25648 26988
rect 26056 26979 26108 26988
rect 26056 26945 26065 26979
rect 26065 26945 26099 26979
rect 26099 26945 26108 26979
rect 26056 26936 26108 26945
rect 20628 26868 20680 26920
rect 22192 26868 22244 26920
rect 23572 26911 23624 26920
rect 23572 26877 23581 26911
rect 23581 26877 23615 26911
rect 23615 26877 23624 26911
rect 23572 26868 23624 26877
rect 24584 26868 24636 26920
rect 26424 26979 26476 26988
rect 26424 26945 26433 26979
rect 26433 26945 26467 26979
rect 26467 26945 26476 26979
rect 26424 26936 26476 26945
rect 33784 27072 33836 27124
rect 34888 27072 34940 27124
rect 26700 27004 26752 27056
rect 27988 27004 28040 27056
rect 29644 27004 29696 27056
rect 31208 27004 31260 27056
rect 28080 26936 28132 26988
rect 31024 26979 31076 26988
rect 20996 26800 21048 26852
rect 26516 26868 26568 26920
rect 10232 26732 10284 26784
rect 11520 26775 11572 26784
rect 11520 26741 11529 26775
rect 11529 26741 11563 26775
rect 11563 26741 11572 26775
rect 11520 26732 11572 26741
rect 14096 26732 14148 26784
rect 14464 26732 14516 26784
rect 19524 26732 19576 26784
rect 20168 26732 20220 26784
rect 24860 26732 24912 26784
rect 26700 26800 26752 26852
rect 27896 26800 27948 26852
rect 28264 26732 28316 26784
rect 31024 26945 31033 26979
rect 31033 26945 31067 26979
rect 31067 26945 31076 26979
rect 32128 27004 32180 27056
rect 32956 27004 33008 27056
rect 35256 27004 35308 27056
rect 31024 26936 31076 26945
rect 32680 26979 32732 26988
rect 32680 26945 32689 26979
rect 32689 26945 32723 26979
rect 32723 26945 32732 26979
rect 32680 26936 32732 26945
rect 35440 26979 35492 26988
rect 35440 26945 35449 26979
rect 35449 26945 35483 26979
rect 35483 26945 35492 26979
rect 35440 26936 35492 26945
rect 37924 27072 37976 27124
rect 38384 27115 38436 27124
rect 38384 27081 38393 27115
rect 38393 27081 38427 27115
rect 38427 27081 38436 27115
rect 38384 27072 38436 27081
rect 36544 26979 36596 26988
rect 36544 26945 36553 26979
rect 36553 26945 36587 26979
rect 36587 26945 36596 26979
rect 36544 26936 36596 26945
rect 36728 26979 36780 26988
rect 36728 26945 36737 26979
rect 36737 26945 36771 26979
rect 36771 26945 36780 26979
rect 36728 26936 36780 26945
rect 31760 26868 31812 26920
rect 34520 26868 34572 26920
rect 35624 26911 35676 26920
rect 35624 26877 35633 26911
rect 35633 26877 35667 26911
rect 35667 26877 35676 26911
rect 35624 26868 35676 26877
rect 36176 26868 36228 26920
rect 37648 26979 37700 26988
rect 37648 26945 37657 26979
rect 37657 26945 37691 26979
rect 37691 26945 37700 26979
rect 37648 26936 37700 26945
rect 37372 26911 37424 26920
rect 37372 26877 37381 26911
rect 37381 26877 37415 26911
rect 37415 26877 37424 26911
rect 37372 26868 37424 26877
rect 37464 26868 37516 26920
rect 38016 26868 38068 26920
rect 37556 26800 37608 26852
rect 38200 26979 38252 26988
rect 38200 26945 38209 26979
rect 38209 26945 38243 26979
rect 38243 26945 38252 26979
rect 38200 26936 38252 26945
rect 30748 26732 30800 26784
rect 33600 26732 33652 26784
rect 37464 26775 37516 26784
rect 37464 26741 37473 26775
rect 37473 26741 37507 26775
rect 37507 26741 37516 26775
rect 37464 26732 37516 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3148 26528 3200 26580
rect 3976 26571 4028 26580
rect 3976 26537 3985 26571
rect 3985 26537 4019 26571
rect 4019 26537 4028 26571
rect 3976 26528 4028 26537
rect 5264 26528 5316 26580
rect 2780 26367 2832 26376
rect 2780 26333 2789 26367
rect 2789 26333 2823 26367
rect 2823 26333 2832 26367
rect 2780 26324 2832 26333
rect 3332 26324 3384 26376
rect 3424 26367 3476 26376
rect 3424 26333 3433 26367
rect 3433 26333 3467 26367
rect 3467 26333 3476 26367
rect 3424 26324 3476 26333
rect 5264 26392 5316 26444
rect 8300 26571 8352 26580
rect 8300 26537 8309 26571
rect 8309 26537 8343 26571
rect 8343 26537 8352 26571
rect 8300 26528 8352 26537
rect 9680 26528 9732 26580
rect 13176 26571 13228 26580
rect 13176 26537 13185 26571
rect 13185 26537 13219 26571
rect 13219 26537 13228 26571
rect 13176 26528 13228 26537
rect 13268 26528 13320 26580
rect 19708 26528 19760 26580
rect 20352 26571 20404 26580
rect 20352 26537 20361 26571
rect 20361 26537 20395 26571
rect 20395 26537 20404 26571
rect 20352 26528 20404 26537
rect 20444 26528 20496 26580
rect 23572 26528 23624 26580
rect 26516 26528 26568 26580
rect 28172 26528 28224 26580
rect 29644 26528 29696 26580
rect 35348 26528 35400 26580
rect 35624 26528 35676 26580
rect 36544 26571 36596 26580
rect 36544 26537 36553 26571
rect 36553 26537 36587 26571
rect 36587 26537 36596 26571
rect 36544 26528 36596 26537
rect 37740 26528 37792 26580
rect 8116 26392 8168 26444
rect 10232 26435 10284 26444
rect 10232 26401 10241 26435
rect 10241 26401 10275 26435
rect 10275 26401 10284 26435
rect 10232 26392 10284 26401
rect 2688 26256 2740 26308
rect 8484 26367 8536 26376
rect 8484 26333 8493 26367
rect 8493 26333 8527 26367
rect 8527 26333 8536 26367
rect 8484 26324 8536 26333
rect 8576 26324 8628 26376
rect 6276 26256 6328 26308
rect 5632 26188 5684 26240
rect 6368 26231 6420 26240
rect 6368 26197 6377 26231
rect 6377 26197 6411 26231
rect 6411 26197 6420 26231
rect 6368 26188 6420 26197
rect 7012 26256 7064 26308
rect 9496 26324 9548 26376
rect 9772 26324 9824 26376
rect 10048 26367 10100 26376
rect 10048 26333 10057 26367
rect 10057 26333 10091 26367
rect 10091 26333 10100 26367
rect 10048 26324 10100 26333
rect 15384 26460 15436 26512
rect 15476 26460 15528 26512
rect 14096 26435 14148 26444
rect 14096 26401 14105 26435
rect 14105 26401 14139 26435
rect 14139 26401 14148 26435
rect 14096 26392 14148 26401
rect 15568 26392 15620 26444
rect 15752 26392 15804 26444
rect 18880 26460 18932 26512
rect 19064 26460 19116 26512
rect 16488 26392 16540 26444
rect 10508 26299 10560 26308
rect 10508 26265 10517 26299
rect 10517 26265 10551 26299
rect 10551 26265 10560 26299
rect 10508 26256 10560 26265
rect 11796 26256 11848 26308
rect 12624 26256 12676 26308
rect 13452 26324 13504 26376
rect 13728 26324 13780 26376
rect 14464 26367 14516 26376
rect 14464 26333 14473 26367
rect 14473 26333 14507 26367
rect 14507 26333 14516 26367
rect 14464 26324 14516 26333
rect 9588 26188 9640 26240
rect 11980 26231 12032 26240
rect 11980 26197 11989 26231
rect 11989 26197 12023 26231
rect 12023 26197 12032 26231
rect 11980 26188 12032 26197
rect 13084 26188 13136 26240
rect 13636 26188 13688 26240
rect 15200 26256 15252 26308
rect 15660 26324 15712 26376
rect 17316 26367 17368 26376
rect 17316 26333 17325 26367
rect 17325 26333 17359 26367
rect 17359 26333 17368 26367
rect 17316 26324 17368 26333
rect 17500 26367 17552 26376
rect 17500 26333 17513 26367
rect 17513 26333 17552 26367
rect 17500 26324 17552 26333
rect 17960 26367 18012 26376
rect 17960 26333 17969 26367
rect 17969 26333 18003 26367
rect 18003 26333 18012 26367
rect 17960 26324 18012 26333
rect 18144 26367 18196 26376
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 18420 26324 18472 26376
rect 18788 26367 18840 26376
rect 18788 26333 18797 26367
rect 18797 26333 18831 26367
rect 18831 26333 18840 26367
rect 18788 26324 18840 26333
rect 18972 26324 19024 26376
rect 14004 26188 14056 26240
rect 14464 26188 14516 26240
rect 14740 26231 14792 26240
rect 14740 26197 14749 26231
rect 14749 26197 14783 26231
rect 14783 26197 14792 26231
rect 14740 26188 14792 26197
rect 15292 26231 15344 26240
rect 15292 26197 15301 26231
rect 15301 26197 15335 26231
rect 15335 26197 15344 26231
rect 15292 26188 15344 26197
rect 16212 26188 16264 26240
rect 16488 26231 16540 26240
rect 16488 26197 16497 26231
rect 16497 26197 16531 26231
rect 16531 26197 16540 26231
rect 16488 26188 16540 26197
rect 17500 26188 17552 26240
rect 19064 26256 19116 26308
rect 19984 26392 20036 26444
rect 19616 26324 19668 26376
rect 21640 26460 21692 26512
rect 24584 26460 24636 26512
rect 24124 26324 24176 26376
rect 24768 26367 24820 26376
rect 24768 26333 24777 26367
rect 24777 26333 24811 26367
rect 24811 26333 24820 26367
rect 24768 26324 24820 26333
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 27804 26460 27856 26512
rect 28816 26460 28868 26512
rect 27620 26392 27672 26444
rect 27896 26435 27948 26444
rect 27896 26401 27905 26435
rect 27905 26401 27939 26435
rect 27939 26401 27948 26435
rect 27896 26392 27948 26401
rect 18604 26188 18656 26240
rect 18696 26231 18748 26240
rect 18696 26197 18705 26231
rect 18705 26197 18739 26231
rect 18739 26197 18748 26231
rect 18696 26188 18748 26197
rect 20628 26188 20680 26240
rect 20812 26188 20864 26240
rect 24032 26299 24084 26308
rect 24032 26265 24041 26299
rect 24041 26265 24075 26299
rect 24075 26265 24084 26299
rect 24032 26256 24084 26265
rect 28264 26367 28316 26376
rect 28264 26333 28273 26367
rect 28273 26333 28307 26367
rect 28307 26333 28316 26367
rect 28264 26324 28316 26333
rect 29092 26367 29144 26376
rect 29092 26333 29101 26367
rect 29101 26333 29135 26367
rect 29135 26333 29144 26367
rect 29092 26324 29144 26333
rect 29828 26392 29880 26444
rect 31208 26460 31260 26512
rect 37372 26460 37424 26512
rect 38016 26460 38068 26512
rect 30104 26392 30156 26444
rect 37464 26392 37516 26444
rect 25596 26256 25648 26308
rect 28540 26299 28592 26308
rect 28540 26265 28549 26299
rect 28549 26265 28583 26299
rect 28583 26265 28592 26299
rect 28540 26256 28592 26265
rect 30104 26299 30156 26308
rect 30104 26265 30113 26299
rect 30113 26265 30147 26299
rect 30147 26265 30156 26299
rect 30104 26256 30156 26265
rect 31024 26367 31076 26376
rect 31024 26333 31033 26367
rect 31033 26333 31067 26367
rect 31067 26333 31076 26367
rect 31024 26324 31076 26333
rect 31208 26367 31260 26376
rect 31208 26333 31217 26367
rect 31217 26333 31251 26367
rect 31251 26333 31260 26367
rect 31208 26324 31260 26333
rect 33784 26324 33836 26376
rect 31668 26256 31720 26308
rect 32680 26256 32732 26308
rect 35992 26324 36044 26376
rect 36084 26367 36136 26376
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 36176 26367 36228 26376
rect 36176 26333 36185 26367
rect 36185 26333 36219 26367
rect 36219 26333 36228 26367
rect 36176 26324 36228 26333
rect 36728 26324 36780 26376
rect 37372 26324 37424 26376
rect 37648 26256 37700 26308
rect 24308 26188 24360 26240
rect 29184 26231 29236 26240
rect 29184 26197 29193 26231
rect 29193 26197 29227 26231
rect 29227 26197 29236 26231
rect 29184 26188 29236 26197
rect 30932 26188 30984 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 8484 25984 8536 26036
rect 5632 25959 5684 25968
rect 5632 25925 5641 25959
rect 5641 25925 5675 25959
rect 5675 25925 5684 25959
rect 5632 25916 5684 25925
rect 3240 25891 3292 25900
rect 3240 25857 3249 25891
rect 3249 25857 3283 25891
rect 3283 25857 3292 25891
rect 3240 25848 3292 25857
rect 3332 25848 3384 25900
rect 5816 25891 5868 25900
rect 5816 25857 5825 25891
rect 5825 25857 5859 25891
rect 5859 25857 5868 25891
rect 5816 25848 5868 25857
rect 6092 25891 6144 25900
rect 6092 25857 6101 25891
rect 6101 25857 6135 25891
rect 6135 25857 6144 25891
rect 6092 25848 6144 25857
rect 6000 25780 6052 25832
rect 6368 25780 6420 25832
rect 6828 25712 6880 25764
rect 8576 25916 8628 25968
rect 9496 25984 9548 26036
rect 9588 26027 9640 26036
rect 9588 25993 9597 26027
rect 9597 25993 9631 26027
rect 9631 25993 9640 26027
rect 9588 25984 9640 25993
rect 11520 25984 11572 26036
rect 13176 25984 13228 26036
rect 10140 25916 10192 25968
rect 8852 25891 8904 25900
rect 8852 25857 8861 25891
rect 8861 25857 8895 25891
rect 8895 25857 8904 25891
rect 8852 25848 8904 25857
rect 8392 25780 8444 25832
rect 11980 25848 12032 25900
rect 10140 25823 10192 25832
rect 4068 25644 4120 25696
rect 7104 25644 7156 25696
rect 8116 25712 8168 25764
rect 10140 25789 10149 25823
rect 10149 25789 10183 25823
rect 10183 25789 10192 25823
rect 10140 25780 10192 25789
rect 10508 25780 10560 25832
rect 9772 25755 9824 25764
rect 9772 25721 9781 25755
rect 9781 25721 9815 25755
rect 9815 25721 9824 25755
rect 9772 25712 9824 25721
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 15844 25984 15896 26036
rect 17960 25984 18012 26036
rect 19156 25984 19208 26036
rect 14096 25891 14148 25900
rect 14096 25857 14105 25891
rect 14105 25857 14139 25891
rect 14139 25857 14148 25891
rect 14096 25848 14148 25857
rect 14280 25848 14332 25900
rect 14372 25891 14424 25900
rect 14372 25857 14381 25891
rect 14381 25857 14415 25891
rect 14415 25857 14424 25891
rect 14372 25848 14424 25857
rect 14924 25891 14976 25900
rect 14924 25857 14933 25891
rect 14933 25857 14967 25891
rect 14967 25857 14976 25891
rect 14924 25848 14976 25857
rect 13084 25823 13136 25832
rect 13084 25789 13093 25823
rect 13093 25789 13127 25823
rect 13127 25789 13136 25823
rect 13084 25780 13136 25789
rect 13820 25780 13872 25832
rect 14464 25780 14516 25832
rect 15200 25823 15252 25832
rect 15200 25789 15209 25823
rect 15209 25789 15243 25823
rect 15243 25789 15252 25823
rect 15200 25780 15252 25789
rect 15660 25848 15712 25900
rect 17316 25916 17368 25968
rect 16212 25891 16264 25900
rect 16212 25857 16221 25891
rect 16221 25857 16255 25891
rect 16255 25857 16264 25891
rect 16212 25848 16264 25857
rect 17868 25916 17920 25968
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 18144 25848 18196 25900
rect 18512 25891 18564 25900
rect 18512 25857 18521 25891
rect 18521 25857 18555 25891
rect 18555 25857 18564 25891
rect 18512 25848 18564 25857
rect 18696 25891 18748 25900
rect 18696 25857 18705 25891
rect 18705 25857 18739 25891
rect 18739 25857 18748 25891
rect 18696 25848 18748 25857
rect 18880 25891 18932 25900
rect 18880 25857 18889 25891
rect 18889 25857 18923 25891
rect 18923 25857 18932 25891
rect 18880 25848 18932 25857
rect 19064 25891 19116 25900
rect 19064 25857 19073 25891
rect 19073 25857 19107 25891
rect 19107 25857 19116 25891
rect 19064 25848 19116 25857
rect 18328 25780 18380 25832
rect 13636 25712 13688 25764
rect 18604 25712 18656 25764
rect 19524 25891 19576 25900
rect 19524 25857 19533 25891
rect 19533 25857 19567 25891
rect 19567 25857 19576 25891
rect 19524 25848 19576 25857
rect 20812 25984 20864 26036
rect 20352 25848 20404 25900
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 20812 25848 20864 25900
rect 21272 25959 21324 25968
rect 21272 25925 21281 25959
rect 21281 25925 21315 25959
rect 21315 25925 21324 25959
rect 21272 25916 21324 25925
rect 24032 25984 24084 26036
rect 21640 25916 21692 25968
rect 19248 25780 19300 25832
rect 20904 25712 20956 25764
rect 10048 25644 10100 25696
rect 11152 25644 11204 25696
rect 13268 25644 13320 25696
rect 13544 25644 13596 25696
rect 17684 25644 17736 25696
rect 18236 25644 18288 25696
rect 18972 25644 19024 25696
rect 19892 25644 19944 25696
rect 22284 25891 22336 25900
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 22284 25848 22336 25857
rect 22560 25848 22612 25900
rect 23112 25891 23164 25900
rect 23112 25857 23146 25891
rect 23146 25857 23164 25891
rect 23112 25848 23164 25857
rect 26056 25984 26108 26036
rect 24308 25916 24360 25968
rect 29184 25984 29236 26036
rect 29828 26027 29880 26036
rect 29828 25993 29837 26027
rect 29837 25993 29871 26027
rect 29871 25993 29880 26027
rect 29828 25984 29880 25993
rect 30288 25984 30340 26036
rect 31668 25984 31720 26036
rect 29644 25916 29696 25968
rect 32404 25959 32456 25968
rect 32404 25925 32413 25959
rect 32413 25925 32447 25959
rect 32447 25925 32456 25959
rect 32404 25916 32456 25925
rect 25228 25891 25280 25900
rect 25228 25857 25237 25891
rect 25237 25857 25271 25891
rect 25271 25857 25280 25891
rect 25228 25848 25280 25857
rect 26332 25848 26384 25900
rect 27804 25891 27856 25900
rect 27804 25857 27813 25891
rect 27813 25857 27847 25891
rect 27847 25857 27856 25891
rect 27804 25848 27856 25857
rect 27896 25891 27948 25900
rect 27896 25857 27905 25891
rect 27905 25857 27939 25891
rect 27939 25857 27948 25891
rect 27896 25848 27948 25857
rect 29828 25848 29880 25900
rect 31116 25848 31168 25900
rect 31576 25848 31628 25900
rect 32312 25891 32364 25900
rect 32312 25857 32321 25891
rect 32321 25857 32355 25891
rect 32355 25857 32364 25891
rect 32312 25848 32364 25857
rect 22192 25823 22244 25832
rect 22192 25789 22201 25823
rect 22201 25789 22235 25823
rect 22235 25789 22244 25823
rect 22192 25780 22244 25789
rect 25872 25780 25924 25832
rect 27712 25780 27764 25832
rect 28080 25823 28132 25832
rect 28080 25789 28089 25823
rect 28089 25789 28123 25823
rect 28123 25789 28132 25823
rect 28080 25780 28132 25789
rect 21364 25687 21416 25696
rect 21364 25653 21373 25687
rect 21373 25653 21407 25687
rect 21407 25653 21416 25687
rect 21364 25644 21416 25653
rect 22100 25687 22152 25696
rect 22100 25653 22109 25687
rect 22109 25653 22143 25687
rect 22143 25653 22152 25687
rect 22100 25644 22152 25653
rect 22652 25644 22704 25696
rect 22836 25644 22888 25696
rect 26884 25712 26936 25764
rect 27528 25712 27580 25764
rect 24308 25687 24360 25696
rect 24308 25653 24317 25687
rect 24317 25653 24351 25687
rect 24351 25653 24360 25687
rect 24308 25644 24360 25653
rect 29092 25644 29144 25696
rect 32956 25891 33008 25900
rect 32956 25857 32965 25891
rect 32965 25857 32999 25891
rect 32999 25857 33008 25891
rect 32956 25848 33008 25857
rect 33140 25823 33192 25832
rect 33140 25789 33149 25823
rect 33149 25789 33183 25823
rect 33183 25789 33192 25823
rect 33140 25780 33192 25789
rect 33600 25891 33652 25900
rect 33600 25857 33609 25891
rect 33609 25857 33643 25891
rect 33643 25857 33652 25891
rect 33600 25848 33652 25857
rect 34336 25891 34388 25900
rect 34336 25857 34345 25891
rect 34345 25857 34379 25891
rect 34379 25857 34388 25891
rect 34336 25848 34388 25857
rect 35992 25984 36044 26036
rect 36084 25984 36136 26036
rect 34796 25916 34848 25968
rect 35440 25891 35492 25900
rect 35440 25857 35449 25891
rect 35449 25857 35483 25891
rect 35483 25857 35492 25891
rect 35440 25848 35492 25857
rect 37464 25916 37516 25968
rect 37832 25891 37884 25900
rect 37832 25857 37841 25891
rect 37841 25857 37875 25891
rect 37875 25857 37884 25891
rect 37832 25848 37884 25857
rect 37556 25780 37608 25832
rect 35992 25712 36044 25764
rect 33140 25644 33192 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3332 25440 3384 25492
rect 3148 25372 3200 25424
rect 6092 25483 6144 25492
rect 6092 25449 6101 25483
rect 6101 25449 6135 25483
rect 6135 25449 6144 25483
rect 6092 25440 6144 25449
rect 7012 25440 7064 25492
rect 8116 25440 8168 25492
rect 9220 25440 9272 25492
rect 11152 25440 11204 25492
rect 13176 25440 13228 25492
rect 6000 25372 6052 25424
rect 8852 25372 8904 25424
rect 14096 25440 14148 25492
rect 14832 25440 14884 25492
rect 15384 25440 15436 25492
rect 15568 25483 15620 25492
rect 15568 25449 15577 25483
rect 15577 25449 15611 25483
rect 15611 25449 15620 25483
rect 15568 25440 15620 25449
rect 15660 25483 15712 25492
rect 15660 25449 15669 25483
rect 15669 25449 15703 25483
rect 15703 25449 15712 25483
rect 15660 25440 15712 25449
rect 18512 25440 18564 25492
rect 20076 25483 20128 25492
rect 20076 25449 20085 25483
rect 20085 25449 20119 25483
rect 20119 25449 20128 25483
rect 20076 25440 20128 25449
rect 21456 25440 21508 25492
rect 21824 25440 21876 25492
rect 23112 25440 23164 25492
rect 25688 25440 25740 25492
rect 26976 25440 27028 25492
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 2688 25304 2740 25356
rect 4068 25347 4120 25356
rect 4068 25313 4077 25347
rect 4077 25313 4111 25347
rect 4111 25313 4120 25347
rect 4068 25304 4120 25313
rect 3056 25236 3108 25288
rect 1768 25168 1820 25220
rect 2964 25168 3016 25220
rect 5632 25279 5684 25288
rect 5632 25245 5641 25279
rect 5641 25245 5675 25279
rect 5675 25245 5684 25279
rect 5632 25236 5684 25245
rect 3148 25143 3200 25152
rect 3148 25109 3157 25143
rect 3157 25109 3191 25143
rect 3191 25109 3200 25143
rect 3148 25100 3200 25109
rect 6828 25236 6880 25288
rect 7104 25279 7156 25288
rect 7104 25245 7113 25279
rect 7113 25245 7147 25279
rect 7147 25245 7156 25279
rect 7104 25236 7156 25245
rect 8392 25304 8444 25356
rect 14924 25372 14976 25424
rect 18144 25372 18196 25424
rect 6184 25168 6236 25220
rect 6368 25168 6420 25220
rect 9220 25236 9272 25288
rect 9496 25236 9548 25288
rect 12072 25236 12124 25288
rect 12808 25236 12860 25288
rect 12992 25279 13044 25288
rect 12992 25245 13001 25279
rect 13001 25245 13035 25279
rect 13035 25245 13044 25279
rect 12992 25236 13044 25245
rect 13268 25279 13320 25288
rect 13268 25245 13303 25279
rect 13303 25245 13320 25279
rect 13268 25236 13320 25245
rect 15292 25304 15344 25356
rect 15568 25304 15620 25356
rect 9036 25168 9088 25220
rect 11152 25168 11204 25220
rect 4712 25100 4764 25152
rect 5724 25143 5776 25152
rect 5724 25109 5733 25143
rect 5733 25109 5767 25143
rect 5767 25109 5776 25143
rect 5724 25100 5776 25109
rect 5908 25143 5960 25152
rect 5908 25109 5917 25143
rect 5917 25109 5951 25143
rect 5951 25109 5960 25143
rect 5908 25100 5960 25109
rect 8484 25143 8536 25152
rect 8484 25109 8493 25143
rect 8493 25109 8527 25143
rect 8527 25109 8536 25143
rect 8484 25100 8536 25109
rect 10324 25143 10376 25152
rect 10324 25109 10333 25143
rect 10333 25109 10367 25143
rect 10367 25109 10376 25143
rect 10324 25100 10376 25109
rect 11060 25143 11112 25152
rect 11060 25109 11069 25143
rect 11069 25109 11103 25143
rect 11103 25109 11112 25143
rect 12624 25143 12676 25152
rect 11060 25100 11112 25109
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 14372 25168 14424 25220
rect 14740 25100 14792 25152
rect 15384 25279 15436 25288
rect 15384 25245 15393 25279
rect 15393 25245 15427 25279
rect 15427 25245 15436 25279
rect 15384 25236 15436 25245
rect 15752 25236 15804 25288
rect 18328 25347 18380 25356
rect 18328 25313 18337 25347
rect 18337 25313 18371 25347
rect 18371 25313 18380 25347
rect 18328 25304 18380 25313
rect 16304 25279 16356 25288
rect 16304 25245 16313 25279
rect 16313 25245 16347 25279
rect 16347 25245 16356 25279
rect 16304 25236 16356 25245
rect 17960 25236 18012 25288
rect 18144 25279 18196 25288
rect 18144 25245 18153 25279
rect 18153 25245 18187 25279
rect 18187 25245 18196 25279
rect 18144 25236 18196 25245
rect 18236 25236 18288 25288
rect 15476 25168 15528 25220
rect 16396 25168 16448 25220
rect 21364 25372 21416 25424
rect 27528 25372 27580 25424
rect 21640 25304 21692 25356
rect 22744 25304 22796 25356
rect 18604 25279 18656 25288
rect 18604 25245 18613 25279
rect 18613 25245 18647 25279
rect 18647 25245 18656 25279
rect 18604 25236 18656 25245
rect 19892 25279 19944 25288
rect 19892 25245 19901 25279
rect 19901 25245 19935 25279
rect 19935 25245 19944 25279
rect 19892 25236 19944 25245
rect 20536 25236 20588 25288
rect 20812 25236 20864 25288
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 20720 25168 20772 25220
rect 21364 25233 21416 25285
rect 22008 25279 22060 25288
rect 22008 25245 22017 25279
rect 22017 25245 22051 25279
rect 22051 25245 22060 25279
rect 22008 25236 22060 25245
rect 22284 25236 22336 25288
rect 22652 25279 22704 25288
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 22836 25279 22888 25288
rect 22836 25245 22845 25279
rect 22845 25245 22879 25279
rect 22879 25245 22888 25279
rect 22836 25236 22888 25245
rect 27896 25304 27948 25356
rect 24308 25236 24360 25288
rect 27988 25279 28040 25288
rect 27988 25245 27997 25279
rect 27997 25245 28031 25279
rect 28031 25245 28040 25279
rect 27988 25236 28040 25245
rect 28172 25279 28224 25288
rect 28172 25245 28181 25279
rect 28181 25245 28215 25279
rect 28215 25245 28224 25279
rect 28172 25236 28224 25245
rect 30288 25304 30340 25356
rect 15752 25100 15804 25152
rect 18788 25100 18840 25152
rect 18880 25100 18932 25152
rect 21180 25100 21232 25152
rect 21272 25100 21324 25152
rect 21640 25143 21692 25152
rect 21640 25109 21643 25143
rect 21643 25109 21677 25143
rect 21677 25109 21692 25143
rect 21640 25100 21692 25109
rect 24768 25143 24820 25152
rect 24768 25109 24777 25143
rect 24777 25109 24811 25143
rect 24811 25109 24820 25143
rect 24768 25100 24820 25109
rect 25044 25100 25096 25152
rect 26332 25168 26384 25220
rect 25320 25100 25372 25152
rect 25872 25143 25924 25152
rect 25872 25109 25881 25143
rect 25881 25109 25915 25143
rect 25915 25109 25924 25143
rect 25872 25100 25924 25109
rect 26884 25168 26936 25220
rect 30932 25279 30984 25288
rect 30932 25245 30941 25279
rect 30941 25245 30975 25279
rect 30975 25245 30984 25279
rect 30932 25236 30984 25245
rect 31208 25279 31260 25288
rect 31208 25245 31217 25279
rect 31217 25245 31251 25279
rect 31251 25245 31260 25279
rect 31208 25236 31260 25245
rect 32312 25440 32364 25492
rect 33140 25440 33192 25492
rect 34336 25440 34388 25492
rect 36728 25483 36780 25492
rect 36728 25449 36737 25483
rect 36737 25449 36771 25483
rect 36771 25449 36780 25483
rect 36728 25440 36780 25449
rect 31576 25347 31628 25356
rect 31576 25313 31585 25347
rect 31585 25313 31619 25347
rect 31619 25313 31628 25347
rect 31576 25304 31628 25313
rect 35992 25372 36044 25424
rect 37464 25440 37516 25492
rect 37832 25483 37884 25492
rect 37832 25449 37841 25483
rect 37841 25449 37875 25483
rect 37875 25449 37884 25483
rect 37832 25440 37884 25449
rect 32220 25279 32272 25288
rect 32220 25245 32229 25279
rect 32229 25245 32263 25279
rect 32263 25245 32272 25279
rect 32220 25236 32272 25245
rect 29092 25168 29144 25220
rect 30748 25211 30800 25220
rect 30748 25177 30757 25211
rect 30757 25177 30791 25211
rect 30791 25177 30800 25211
rect 30748 25168 30800 25177
rect 31116 25168 31168 25220
rect 32128 25168 32180 25220
rect 32680 25279 32732 25288
rect 32680 25245 32689 25279
rect 32689 25245 32723 25279
rect 32723 25245 32732 25279
rect 32680 25236 32732 25245
rect 32588 25168 32640 25220
rect 33416 25279 33468 25288
rect 33416 25245 33425 25279
rect 33425 25245 33459 25279
rect 33459 25245 33468 25279
rect 33416 25236 33468 25245
rect 33600 25279 33652 25288
rect 33600 25245 33609 25279
rect 33609 25245 33643 25279
rect 33643 25245 33652 25279
rect 33600 25236 33652 25245
rect 37096 25304 37148 25356
rect 34704 25211 34756 25220
rect 34704 25177 34713 25211
rect 34713 25177 34747 25211
rect 34747 25177 34756 25211
rect 34704 25168 34756 25177
rect 34888 25211 34940 25220
rect 34888 25177 34897 25211
rect 34897 25177 34931 25211
rect 34931 25177 34940 25211
rect 34888 25168 34940 25177
rect 27436 25100 27488 25152
rect 29828 25143 29880 25152
rect 29828 25109 29837 25143
rect 29837 25109 29871 25143
rect 29871 25109 29880 25143
rect 29828 25100 29880 25109
rect 32956 25100 33008 25152
rect 36912 25236 36964 25288
rect 37740 25236 37792 25288
rect 37924 25279 37976 25288
rect 37924 25245 37933 25279
rect 37933 25245 37967 25279
rect 37967 25245 37976 25279
rect 37924 25236 37976 25245
rect 37004 25143 37056 25152
rect 37004 25109 37031 25143
rect 37031 25109 37056 25143
rect 37004 25100 37056 25109
rect 37096 25100 37148 25152
rect 37832 25100 37884 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 6092 24896 6144 24948
rect 1308 24624 1360 24676
rect 1768 24735 1820 24744
rect 1768 24701 1777 24735
rect 1777 24701 1811 24735
rect 1811 24701 1820 24735
rect 1768 24692 1820 24701
rect 2044 24735 2096 24744
rect 2044 24701 2053 24735
rect 2053 24701 2087 24735
rect 2087 24701 2096 24735
rect 2044 24692 2096 24701
rect 2872 24760 2924 24812
rect 4712 24828 4764 24880
rect 6276 24828 6328 24880
rect 8024 24896 8076 24948
rect 9588 24896 9640 24948
rect 12992 24896 13044 24948
rect 15200 24896 15252 24948
rect 6368 24760 6420 24812
rect 8116 24828 8168 24880
rect 9036 24871 9088 24880
rect 9036 24837 9045 24871
rect 9045 24837 9079 24871
rect 9079 24837 9088 24871
rect 9036 24828 9088 24837
rect 3148 24692 3200 24744
rect 3884 24692 3936 24744
rect 5724 24692 5776 24744
rect 7012 24692 7064 24744
rect 7656 24760 7708 24812
rect 8208 24803 8260 24812
rect 8208 24769 8217 24803
rect 8217 24769 8251 24803
rect 8251 24769 8260 24803
rect 8208 24760 8260 24769
rect 8484 24803 8536 24812
rect 8484 24769 8493 24803
rect 8493 24769 8527 24803
rect 8527 24769 8536 24803
rect 8484 24760 8536 24769
rect 8760 24803 8812 24812
rect 8760 24769 8769 24803
rect 8769 24769 8803 24803
rect 8803 24769 8812 24803
rect 8760 24760 8812 24769
rect 7288 24735 7340 24744
rect 7288 24701 7297 24735
rect 7297 24701 7331 24735
rect 7331 24701 7340 24735
rect 7288 24692 7340 24701
rect 7840 24692 7892 24744
rect 9128 24803 9180 24812
rect 9128 24769 9137 24803
rect 9137 24769 9171 24803
rect 9171 24769 9180 24803
rect 9128 24760 9180 24769
rect 9680 24760 9732 24812
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 10324 24692 10376 24744
rect 10784 24803 10836 24812
rect 10784 24769 10793 24803
rect 10793 24769 10827 24803
rect 10827 24769 10836 24803
rect 10784 24760 10836 24769
rect 12072 24803 12124 24812
rect 12072 24769 12081 24803
rect 12081 24769 12115 24803
rect 12115 24769 12124 24803
rect 12072 24760 12124 24769
rect 12716 24760 12768 24812
rect 13084 24760 13136 24812
rect 13452 24760 13504 24812
rect 13912 24803 13964 24812
rect 13912 24769 13921 24803
rect 13921 24769 13955 24803
rect 13955 24769 13964 24803
rect 13912 24760 13964 24769
rect 14832 24828 14884 24880
rect 15844 24896 15896 24948
rect 16304 24896 16356 24948
rect 18144 24896 18196 24948
rect 19064 24896 19116 24948
rect 9864 24624 9916 24676
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 18788 24871 18840 24880
rect 18788 24837 18797 24871
rect 18797 24837 18831 24871
rect 18831 24837 18840 24871
rect 18788 24828 18840 24837
rect 19984 24896 20036 24948
rect 20260 24896 20312 24948
rect 21824 24896 21876 24948
rect 22192 24896 22244 24948
rect 30748 24896 30800 24948
rect 31208 24896 31260 24948
rect 32588 24939 32640 24948
rect 32588 24905 32597 24939
rect 32597 24905 32631 24939
rect 32631 24905 32640 24939
rect 32588 24896 32640 24905
rect 32680 24939 32732 24948
rect 32680 24905 32689 24939
rect 32689 24905 32723 24939
rect 32723 24905 32732 24939
rect 32680 24896 32732 24905
rect 33416 24896 33468 24948
rect 20444 24828 20496 24880
rect 15660 24760 15712 24812
rect 15752 24803 15804 24812
rect 15752 24769 15761 24803
rect 15761 24769 15795 24803
rect 15795 24769 15804 24803
rect 15752 24760 15804 24769
rect 15844 24803 15896 24812
rect 15844 24769 15853 24803
rect 15853 24769 15887 24803
rect 15887 24769 15896 24803
rect 15844 24760 15896 24769
rect 15384 24692 15436 24744
rect 16212 24760 16264 24812
rect 17776 24760 17828 24812
rect 18696 24760 18748 24812
rect 18420 24692 18472 24744
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 19984 24760 20036 24812
rect 20536 24760 20588 24812
rect 22008 24828 22060 24880
rect 24768 24871 24820 24880
rect 24768 24837 24777 24871
rect 24777 24837 24811 24871
rect 24811 24837 24820 24871
rect 24768 24828 24820 24837
rect 25504 24828 25556 24880
rect 21824 24803 21876 24812
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 22100 24803 22152 24812
rect 22100 24769 22109 24803
rect 22109 24769 22143 24803
rect 22143 24769 22152 24803
rect 22100 24760 22152 24769
rect 19340 24692 19392 24744
rect 20904 24692 20956 24744
rect 15752 24624 15804 24676
rect 2044 24556 2096 24608
rect 2964 24556 3016 24608
rect 3424 24556 3476 24608
rect 6092 24556 6144 24608
rect 6552 24556 6604 24608
rect 6920 24556 6972 24608
rect 7472 24556 7524 24608
rect 8116 24556 8168 24608
rect 9220 24599 9272 24608
rect 9220 24565 9229 24599
rect 9229 24565 9263 24599
rect 9263 24565 9272 24599
rect 9220 24556 9272 24565
rect 9312 24556 9364 24608
rect 10508 24556 10560 24608
rect 15568 24556 15620 24608
rect 21272 24599 21324 24608
rect 21272 24565 21281 24599
rect 21281 24565 21315 24599
rect 21315 24565 21324 24599
rect 21272 24556 21324 24565
rect 22008 24735 22060 24744
rect 22008 24701 22017 24735
rect 22017 24701 22051 24735
rect 22051 24701 22060 24735
rect 22652 24803 22704 24812
rect 22652 24769 22661 24803
rect 22661 24769 22695 24803
rect 22695 24769 22704 24803
rect 22652 24760 22704 24769
rect 23296 24803 23348 24812
rect 23296 24769 23330 24803
rect 23330 24769 23348 24803
rect 23296 24760 23348 24769
rect 24216 24760 24268 24812
rect 26424 24760 26476 24812
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 27436 24760 27488 24769
rect 28632 24760 28684 24812
rect 22008 24692 22060 24701
rect 22468 24735 22520 24744
rect 22468 24701 22477 24735
rect 22477 24701 22511 24735
rect 22511 24701 22520 24735
rect 22468 24692 22520 24701
rect 22928 24692 22980 24744
rect 26976 24735 27028 24744
rect 26976 24701 26985 24735
rect 26985 24701 27019 24735
rect 27019 24701 27028 24735
rect 26976 24692 27028 24701
rect 26700 24624 26752 24676
rect 27160 24624 27212 24676
rect 29092 24735 29144 24744
rect 29092 24701 29101 24735
rect 29101 24701 29135 24735
rect 29135 24701 29144 24735
rect 29092 24692 29144 24701
rect 29552 24735 29604 24744
rect 29552 24701 29561 24735
rect 29561 24701 29595 24735
rect 29595 24701 29604 24735
rect 29552 24692 29604 24701
rect 30840 24803 30892 24812
rect 30840 24769 30849 24803
rect 30849 24769 30883 24803
rect 30883 24769 30892 24803
rect 30840 24760 30892 24769
rect 31116 24803 31168 24812
rect 31116 24769 31125 24803
rect 31125 24769 31159 24803
rect 31159 24769 31168 24803
rect 31116 24760 31168 24769
rect 31576 24871 31628 24880
rect 31576 24837 31585 24871
rect 31585 24837 31619 24871
rect 31619 24837 31628 24871
rect 31576 24828 31628 24837
rect 32128 24803 32180 24812
rect 32128 24769 32137 24803
rect 32137 24769 32171 24803
rect 32171 24769 32180 24803
rect 32128 24760 32180 24769
rect 31576 24692 31628 24744
rect 32680 24803 32732 24812
rect 32680 24769 32689 24803
rect 32689 24769 32723 24803
rect 32723 24769 32732 24803
rect 32680 24760 32732 24769
rect 29000 24624 29052 24676
rect 32220 24624 32272 24676
rect 32312 24624 32364 24676
rect 22284 24599 22336 24608
rect 22284 24565 22293 24599
rect 22293 24565 22327 24599
rect 22327 24565 22336 24599
rect 22284 24556 22336 24565
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 25228 24556 25280 24608
rect 26240 24599 26292 24608
rect 26240 24565 26249 24599
rect 26249 24565 26283 24599
rect 26283 24565 26292 24599
rect 26240 24556 26292 24565
rect 32128 24556 32180 24608
rect 33600 24871 33652 24880
rect 33600 24837 33609 24871
rect 33609 24837 33643 24871
rect 33643 24837 33652 24871
rect 33600 24828 33652 24837
rect 33784 24760 33836 24812
rect 34704 24896 34756 24948
rect 35440 24896 35492 24948
rect 35992 24939 36044 24948
rect 35992 24905 36001 24939
rect 36001 24905 36035 24939
rect 36035 24905 36044 24939
rect 35992 24896 36044 24905
rect 33692 24624 33744 24676
rect 33876 24624 33928 24676
rect 33784 24556 33836 24608
rect 34796 24760 34848 24812
rect 35440 24760 35492 24812
rect 36820 24803 36872 24812
rect 36820 24769 36829 24803
rect 36829 24769 36863 24803
rect 36863 24769 36872 24803
rect 36820 24760 36872 24769
rect 37004 24803 37056 24812
rect 37004 24769 37013 24803
rect 37013 24769 37047 24803
rect 37047 24769 37056 24803
rect 37004 24760 37056 24769
rect 34888 24667 34940 24676
rect 34888 24633 34897 24667
rect 34897 24633 34931 24667
rect 34931 24633 34940 24667
rect 34888 24624 34940 24633
rect 35532 24692 35584 24744
rect 37096 24624 37148 24676
rect 35440 24599 35492 24608
rect 35440 24565 35449 24599
rect 35449 24565 35483 24599
rect 35483 24565 35492 24599
rect 35440 24556 35492 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3240 24395 3292 24404
rect 3240 24361 3249 24395
rect 3249 24361 3283 24395
rect 3283 24361 3292 24395
rect 3240 24352 3292 24361
rect 3976 24352 4028 24404
rect 5632 24395 5684 24404
rect 5632 24361 5641 24395
rect 5641 24361 5675 24395
rect 5675 24361 5684 24395
rect 5632 24352 5684 24361
rect 7288 24352 7340 24404
rect 7380 24395 7432 24404
rect 7380 24361 7389 24395
rect 7389 24361 7423 24395
rect 7423 24361 7432 24395
rect 7380 24352 7432 24361
rect 7840 24395 7892 24404
rect 7840 24361 7849 24395
rect 7849 24361 7883 24395
rect 7883 24361 7892 24395
rect 7840 24352 7892 24361
rect 9312 24352 9364 24404
rect 9496 24352 9548 24404
rect 12072 24352 12124 24404
rect 4988 24327 5040 24336
rect 4988 24293 4997 24327
rect 4997 24293 5031 24327
rect 5031 24293 5040 24327
rect 4988 24284 5040 24293
rect 2964 24191 3016 24200
rect 2964 24157 2973 24191
rect 2973 24157 3007 24191
rect 3007 24157 3016 24191
rect 2964 24148 3016 24157
rect 3424 24216 3476 24268
rect 4712 24259 4764 24268
rect 4712 24225 4721 24259
rect 4721 24225 4755 24259
rect 4755 24225 4764 24259
rect 4712 24216 4764 24225
rect 6552 24259 6604 24268
rect 6552 24225 6561 24259
rect 6561 24225 6595 24259
rect 6595 24225 6604 24259
rect 6552 24216 6604 24225
rect 3332 24191 3384 24200
rect 3332 24157 3341 24191
rect 3341 24157 3375 24191
rect 3375 24157 3384 24191
rect 3332 24148 3384 24157
rect 3148 24080 3200 24132
rect 3424 24055 3476 24064
rect 3424 24021 3433 24055
rect 3433 24021 3467 24055
rect 3467 24021 3476 24055
rect 3424 24012 3476 24021
rect 3608 24080 3660 24132
rect 6184 24148 6236 24200
rect 6920 24191 6972 24200
rect 6920 24157 6929 24191
rect 6929 24157 6963 24191
rect 6963 24157 6972 24191
rect 6920 24148 6972 24157
rect 8760 24284 8812 24336
rect 7288 24259 7340 24268
rect 7288 24225 7297 24259
rect 7297 24225 7331 24259
rect 7331 24225 7340 24259
rect 7288 24216 7340 24225
rect 7472 24259 7524 24268
rect 7472 24225 7481 24259
rect 7481 24225 7515 24259
rect 7515 24225 7524 24259
rect 7472 24216 7524 24225
rect 8208 24259 8260 24268
rect 8208 24225 8217 24259
rect 8217 24225 8251 24259
rect 8251 24225 8260 24259
rect 8208 24216 8260 24225
rect 9864 24216 9916 24268
rect 10232 24259 10284 24268
rect 10232 24225 10241 24259
rect 10241 24225 10275 24259
rect 10275 24225 10284 24259
rect 10232 24216 10284 24225
rect 10508 24259 10560 24268
rect 10508 24225 10517 24259
rect 10517 24225 10551 24259
rect 10551 24225 10560 24259
rect 10508 24216 10560 24225
rect 13912 24352 13964 24404
rect 14280 24352 14332 24404
rect 14372 24352 14424 24404
rect 15752 24352 15804 24404
rect 19147 24352 19199 24404
rect 19248 24352 19300 24404
rect 19340 24352 19392 24404
rect 19800 24352 19852 24404
rect 19892 24395 19944 24404
rect 19892 24361 19901 24395
rect 19901 24361 19935 24395
rect 19935 24361 19944 24395
rect 19892 24352 19944 24361
rect 21088 24352 21140 24404
rect 21916 24352 21968 24404
rect 23296 24352 23348 24404
rect 25044 24352 25096 24404
rect 25688 24395 25740 24404
rect 25688 24361 25697 24395
rect 25697 24361 25731 24395
rect 25731 24361 25740 24395
rect 25688 24352 25740 24361
rect 26332 24352 26384 24404
rect 27988 24352 28040 24404
rect 28632 24395 28684 24404
rect 28632 24361 28641 24395
rect 28641 24361 28675 24395
rect 28675 24361 28684 24395
rect 28632 24352 28684 24361
rect 29552 24395 29604 24404
rect 7656 24191 7708 24200
rect 7656 24157 7665 24191
rect 7665 24157 7699 24191
rect 7699 24157 7708 24191
rect 7656 24148 7708 24157
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 9220 24148 9272 24200
rect 12992 24148 13044 24200
rect 13636 24191 13688 24200
rect 13636 24157 13645 24191
rect 13645 24157 13679 24191
rect 13679 24157 13688 24191
rect 13636 24148 13688 24157
rect 15108 24259 15160 24268
rect 15108 24225 15117 24259
rect 15117 24225 15151 24259
rect 15151 24225 15160 24259
rect 15108 24216 15160 24225
rect 15568 24259 15620 24268
rect 15568 24225 15577 24259
rect 15577 24225 15611 24259
rect 15611 24225 15620 24259
rect 15568 24216 15620 24225
rect 16304 24284 16356 24336
rect 14832 24148 14884 24200
rect 16304 24148 16356 24200
rect 16488 24148 16540 24200
rect 17500 24284 17552 24336
rect 19524 24284 19576 24336
rect 20076 24284 20128 24336
rect 21640 24284 21692 24336
rect 22008 24284 22060 24336
rect 22376 24284 22428 24336
rect 18144 24148 18196 24200
rect 18420 24216 18472 24268
rect 18512 24259 18564 24268
rect 18512 24225 18521 24259
rect 18521 24225 18555 24259
rect 18555 24225 18564 24259
rect 18512 24216 18564 24225
rect 20444 24216 20496 24268
rect 7012 24123 7064 24132
rect 7012 24089 7021 24123
rect 7021 24089 7055 24123
rect 7055 24089 7064 24123
rect 7012 24080 7064 24089
rect 7472 24080 7524 24132
rect 8300 24080 8352 24132
rect 9036 24080 9088 24132
rect 11796 24080 11848 24132
rect 15016 24080 15068 24132
rect 17776 24080 17828 24132
rect 18420 24080 18472 24132
rect 18880 24193 18932 24200
rect 18880 24159 18889 24193
rect 18889 24159 18923 24193
rect 18923 24159 18932 24193
rect 18880 24148 18932 24159
rect 19064 24191 19116 24200
rect 19064 24157 19073 24191
rect 19073 24157 19107 24191
rect 19107 24157 19116 24191
rect 19064 24148 19116 24157
rect 19156 24148 19208 24200
rect 20168 24191 20220 24200
rect 20168 24157 20177 24191
rect 20177 24157 20211 24191
rect 20211 24157 20220 24191
rect 20168 24148 20220 24157
rect 20812 24148 20864 24200
rect 19248 24080 19300 24132
rect 20076 24080 20128 24132
rect 21916 24259 21968 24268
rect 21916 24225 21925 24259
rect 21925 24225 21959 24259
rect 21959 24225 21968 24259
rect 21916 24216 21968 24225
rect 21824 24148 21876 24200
rect 22284 24148 22336 24200
rect 25228 24216 25280 24268
rect 26240 24284 26292 24336
rect 28264 24284 28316 24336
rect 29552 24361 29561 24395
rect 29561 24361 29595 24395
rect 29595 24361 29604 24395
rect 29552 24352 29604 24361
rect 31576 24352 31628 24404
rect 32680 24395 32732 24404
rect 32680 24361 32689 24395
rect 32689 24361 32723 24395
rect 32723 24361 32732 24395
rect 32680 24352 32732 24361
rect 33876 24395 33928 24404
rect 33876 24361 33885 24395
rect 33885 24361 33919 24395
rect 33919 24361 33928 24395
rect 33876 24352 33928 24361
rect 35532 24395 35584 24404
rect 35532 24361 35541 24395
rect 35541 24361 35575 24395
rect 35575 24361 35584 24395
rect 35532 24352 35584 24361
rect 37004 24352 37056 24404
rect 22100 24080 22152 24132
rect 25596 24191 25648 24200
rect 25596 24157 25605 24191
rect 25605 24157 25639 24191
rect 25639 24157 25648 24191
rect 25596 24148 25648 24157
rect 27252 24216 27304 24268
rect 23664 24080 23716 24132
rect 24768 24080 24820 24132
rect 26700 24148 26752 24200
rect 27436 24148 27488 24200
rect 28816 24259 28868 24268
rect 28816 24225 28825 24259
rect 28825 24225 28859 24259
rect 28859 24225 28868 24259
rect 28816 24216 28868 24225
rect 29460 24216 29512 24268
rect 6368 24012 6420 24064
rect 8760 24012 8812 24064
rect 14740 24012 14792 24064
rect 15200 24012 15252 24064
rect 16396 24012 16448 24064
rect 16580 24055 16632 24064
rect 16580 24021 16589 24055
rect 16589 24021 16623 24055
rect 16623 24021 16632 24055
rect 16580 24012 16632 24021
rect 18604 24012 18656 24064
rect 18880 24012 18932 24064
rect 21364 24012 21416 24064
rect 21640 24012 21692 24064
rect 22468 24012 22520 24064
rect 22836 24012 22888 24064
rect 25596 24012 25648 24064
rect 27160 24080 27212 24132
rect 26424 24012 26476 24064
rect 26700 24055 26752 24064
rect 26700 24021 26709 24055
rect 26709 24021 26743 24055
rect 26743 24021 26752 24055
rect 26700 24012 26752 24021
rect 27712 24012 27764 24064
rect 30196 24191 30248 24200
rect 30196 24157 30205 24191
rect 30205 24157 30239 24191
rect 30239 24157 30248 24191
rect 30196 24148 30248 24157
rect 30380 24191 30432 24200
rect 30380 24157 30389 24191
rect 30389 24157 30423 24191
rect 30423 24157 30432 24191
rect 30380 24148 30432 24157
rect 29368 24080 29420 24132
rect 31576 24080 31628 24132
rect 28816 24012 28868 24064
rect 28908 24012 28960 24064
rect 30012 24012 30064 24064
rect 32312 24148 32364 24200
rect 33692 24216 33744 24268
rect 36176 24284 36228 24336
rect 36820 24284 36872 24336
rect 32864 24148 32916 24200
rect 33784 24191 33836 24200
rect 33784 24157 33793 24191
rect 33793 24157 33827 24191
rect 33827 24157 33836 24191
rect 33784 24148 33836 24157
rect 34520 24148 34572 24200
rect 36360 24148 36412 24200
rect 36636 24080 36688 24132
rect 37924 24080 37976 24132
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 2964 23808 3016 23860
rect 5172 23808 5224 23860
rect 8208 23808 8260 23860
rect 8300 23808 8352 23860
rect 8576 23851 8628 23860
rect 8576 23817 8585 23851
rect 8585 23817 8619 23851
rect 8619 23817 8628 23851
rect 8576 23808 8628 23817
rect 9036 23808 9088 23860
rect 9588 23808 9640 23860
rect 3056 23740 3108 23792
rect 2964 23672 3016 23724
rect 3332 23672 3384 23724
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 1676 23647 1728 23656
rect 1676 23613 1685 23647
rect 1685 23613 1719 23647
rect 1719 23613 1728 23647
rect 1676 23604 1728 23613
rect 3608 23647 3660 23656
rect 3608 23613 3617 23647
rect 3617 23613 3651 23647
rect 3651 23613 3660 23647
rect 3608 23604 3660 23613
rect 8852 23740 8904 23792
rect 10232 23740 10284 23792
rect 10784 23740 10836 23792
rect 8392 23715 8444 23724
rect 5356 23604 5408 23656
rect 6000 23604 6052 23656
rect 7012 23604 7064 23656
rect 3976 23511 4028 23520
rect 3976 23477 3985 23511
rect 3985 23477 4019 23511
rect 4019 23477 4028 23511
rect 3976 23468 4028 23477
rect 8392 23681 8410 23715
rect 8410 23681 8444 23715
rect 8392 23672 8444 23681
rect 8944 23715 8996 23724
rect 8944 23681 8953 23715
rect 8953 23681 8987 23715
rect 8987 23681 8996 23715
rect 8944 23672 8996 23681
rect 9036 23672 9088 23724
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 9588 23715 9640 23724
rect 9588 23681 9597 23715
rect 9597 23681 9631 23715
rect 9631 23681 9640 23715
rect 9588 23672 9640 23681
rect 9772 23715 9824 23724
rect 9772 23681 9781 23715
rect 9781 23681 9815 23715
rect 9815 23681 9824 23715
rect 9772 23672 9824 23681
rect 10140 23604 10192 23656
rect 11152 23672 11204 23724
rect 13912 23808 13964 23860
rect 13452 23783 13504 23792
rect 13452 23749 13461 23783
rect 13461 23749 13495 23783
rect 13495 23749 13504 23783
rect 13452 23740 13504 23749
rect 14740 23808 14792 23860
rect 14832 23851 14884 23860
rect 14832 23817 14841 23851
rect 14841 23817 14875 23851
rect 14875 23817 14884 23851
rect 14832 23808 14884 23817
rect 18512 23851 18564 23860
rect 18512 23817 18521 23851
rect 18521 23817 18555 23851
rect 18555 23817 18564 23851
rect 18512 23808 18564 23817
rect 19248 23808 19300 23860
rect 15200 23740 15252 23792
rect 14372 23715 14424 23724
rect 14372 23681 14381 23715
rect 14381 23681 14415 23715
rect 14415 23681 14424 23715
rect 14372 23672 14424 23681
rect 12624 23604 12676 23656
rect 9128 23536 9180 23588
rect 12992 23536 13044 23588
rect 15108 23672 15160 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 17500 23715 17552 23724
rect 17500 23681 17509 23715
rect 17509 23681 17543 23715
rect 17543 23681 17552 23715
rect 17500 23672 17552 23681
rect 17960 23783 18012 23792
rect 17960 23749 17969 23783
rect 17969 23749 18003 23783
rect 18003 23749 18012 23783
rect 17960 23740 18012 23749
rect 18696 23740 18748 23792
rect 19064 23740 19116 23792
rect 20076 23808 20128 23860
rect 20352 23808 20404 23860
rect 20628 23808 20680 23860
rect 22008 23808 22060 23860
rect 22560 23808 22612 23860
rect 29000 23851 29052 23860
rect 29000 23817 29009 23851
rect 29009 23817 29043 23851
rect 29043 23817 29052 23851
rect 29000 23808 29052 23817
rect 30196 23808 30248 23860
rect 31576 23808 31628 23860
rect 32864 23851 32916 23860
rect 32864 23817 32873 23851
rect 32873 23817 32907 23851
rect 32907 23817 32916 23851
rect 32864 23808 32916 23817
rect 33692 23808 33744 23860
rect 33784 23808 33836 23860
rect 34520 23851 34572 23860
rect 34520 23817 34529 23851
rect 34529 23817 34563 23851
rect 34563 23817 34572 23851
rect 34520 23808 34572 23817
rect 34796 23808 34848 23860
rect 36360 23851 36412 23860
rect 36360 23817 36369 23851
rect 36369 23817 36403 23851
rect 36403 23817 36412 23851
rect 36360 23808 36412 23817
rect 37924 23851 37976 23860
rect 37924 23817 37933 23851
rect 37933 23817 37967 23851
rect 37967 23817 37976 23851
rect 37924 23808 37976 23817
rect 14188 23536 14240 23588
rect 14464 23536 14516 23588
rect 16580 23604 16632 23656
rect 18880 23672 18932 23724
rect 20168 23740 20220 23792
rect 18144 23604 18196 23656
rect 18788 23647 18840 23656
rect 18788 23613 18797 23647
rect 18797 23613 18831 23647
rect 18831 23613 18840 23647
rect 18788 23604 18840 23613
rect 15016 23579 15068 23588
rect 15016 23545 15025 23579
rect 15025 23545 15059 23579
rect 15059 23545 15068 23579
rect 15016 23536 15068 23545
rect 19340 23672 19392 23724
rect 19984 23715 20036 23724
rect 19984 23681 19993 23715
rect 19993 23681 20027 23715
rect 20027 23681 20036 23715
rect 19984 23672 20036 23681
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 22836 23740 22888 23792
rect 28540 23740 28592 23792
rect 30012 23740 30064 23792
rect 30380 23783 30432 23792
rect 30380 23749 30389 23783
rect 30389 23749 30423 23783
rect 30423 23749 30432 23783
rect 30380 23740 30432 23749
rect 33048 23740 33100 23792
rect 21088 23672 21140 23724
rect 21364 23715 21416 23724
rect 21364 23681 21373 23715
rect 21373 23681 21407 23715
rect 21407 23681 21416 23715
rect 21364 23672 21416 23681
rect 21824 23715 21876 23724
rect 21824 23681 21833 23715
rect 21833 23681 21867 23715
rect 21867 23681 21876 23715
rect 21824 23672 21876 23681
rect 22468 23672 22520 23724
rect 24768 23672 24820 23724
rect 25320 23672 25372 23724
rect 25504 23715 25556 23724
rect 25504 23681 25513 23715
rect 25513 23681 25547 23715
rect 25547 23681 25556 23715
rect 25504 23672 25556 23681
rect 8484 23468 8536 23520
rect 8944 23468 8996 23520
rect 11152 23468 11204 23520
rect 16120 23468 16172 23520
rect 16856 23468 16908 23520
rect 18052 23468 18104 23520
rect 18696 23511 18748 23520
rect 18696 23477 18705 23511
rect 18705 23477 18739 23511
rect 18739 23477 18748 23511
rect 18696 23468 18748 23477
rect 19340 23536 19392 23588
rect 20812 23604 20864 23656
rect 26240 23604 26292 23656
rect 27160 23672 27212 23724
rect 27528 23604 27580 23656
rect 20444 23468 20496 23520
rect 20628 23468 20680 23520
rect 22100 23536 22152 23588
rect 24308 23579 24360 23588
rect 24308 23545 24317 23579
rect 24317 23545 24351 23579
rect 24351 23545 24360 23579
rect 24308 23536 24360 23545
rect 25596 23536 25648 23588
rect 26884 23536 26936 23588
rect 28908 23672 28960 23724
rect 29276 23715 29328 23724
rect 29276 23681 29285 23715
rect 29285 23681 29319 23715
rect 29319 23681 29328 23715
rect 29276 23672 29328 23681
rect 29368 23715 29420 23724
rect 29368 23681 29377 23715
rect 29377 23681 29411 23715
rect 29411 23681 29420 23715
rect 29368 23672 29420 23681
rect 29460 23715 29512 23724
rect 29460 23681 29469 23715
rect 29469 23681 29503 23715
rect 29503 23681 29512 23715
rect 29460 23672 29512 23681
rect 30196 23715 30248 23724
rect 30196 23681 30205 23715
rect 30205 23681 30239 23715
rect 30239 23681 30248 23715
rect 30196 23672 30248 23681
rect 30104 23604 30156 23656
rect 31576 23715 31628 23724
rect 31576 23681 31585 23715
rect 31585 23681 31619 23715
rect 31619 23681 31628 23715
rect 31576 23672 31628 23681
rect 32128 23672 32180 23724
rect 36636 23783 36688 23792
rect 36636 23749 36645 23783
rect 36645 23749 36679 23783
rect 36679 23749 36688 23783
rect 36636 23740 36688 23749
rect 34336 23715 34388 23724
rect 34336 23681 34345 23715
rect 34345 23681 34379 23715
rect 34379 23681 34388 23715
rect 34336 23672 34388 23681
rect 34612 23715 34664 23724
rect 34612 23681 34621 23715
rect 34621 23681 34655 23715
rect 34655 23681 34664 23715
rect 34612 23672 34664 23681
rect 34796 23672 34848 23724
rect 35440 23672 35492 23724
rect 36268 23715 36320 23724
rect 36268 23681 36277 23715
rect 36277 23681 36311 23715
rect 36311 23681 36320 23715
rect 36268 23672 36320 23681
rect 37280 23715 37332 23724
rect 23940 23468 23992 23520
rect 24492 23511 24544 23520
rect 24492 23477 24501 23511
rect 24501 23477 24535 23511
rect 24535 23477 24544 23511
rect 24492 23468 24544 23477
rect 24952 23468 25004 23520
rect 26608 23468 26660 23520
rect 27804 23468 27856 23520
rect 37280 23681 37289 23715
rect 37289 23681 37323 23715
rect 37323 23681 37332 23715
rect 37280 23672 37332 23681
rect 37464 23715 37516 23724
rect 37464 23681 37473 23715
rect 37473 23681 37507 23715
rect 37507 23681 37516 23715
rect 37464 23672 37516 23681
rect 36636 23604 36688 23656
rect 36912 23468 36964 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1676 23264 1728 23316
rect 5172 23307 5224 23316
rect 5172 23273 5181 23307
rect 5181 23273 5215 23307
rect 5215 23273 5224 23307
rect 5172 23264 5224 23273
rect 2044 23060 2096 23112
rect 3424 23196 3476 23248
rect 6828 23264 6880 23316
rect 6460 23196 6512 23248
rect 8760 23196 8812 23248
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 3976 23060 4028 23112
rect 4896 23060 4948 23112
rect 5172 23060 5224 23112
rect 5724 23060 5776 23112
rect 6000 23103 6052 23112
rect 6000 23069 6009 23103
rect 6009 23069 6043 23103
rect 6043 23069 6052 23103
rect 6000 23060 6052 23069
rect 6092 23103 6144 23112
rect 6092 23069 6101 23103
rect 6101 23069 6135 23103
rect 6135 23069 6144 23103
rect 6092 23060 6144 23069
rect 6368 23060 6420 23112
rect 6460 23103 6512 23112
rect 6460 23069 6469 23103
rect 6469 23069 6503 23103
rect 6503 23069 6512 23103
rect 6460 23060 6512 23069
rect 6644 23103 6696 23112
rect 6644 23069 6653 23103
rect 6653 23069 6687 23103
rect 6687 23069 6696 23103
rect 6644 23060 6696 23069
rect 6184 22992 6236 23044
rect 6828 23103 6880 23112
rect 6828 23069 6837 23103
rect 6837 23069 6871 23103
rect 6871 23069 6880 23103
rect 6828 23060 6880 23069
rect 8484 23060 8536 23112
rect 9220 23264 9272 23316
rect 18604 23264 18656 23316
rect 20536 23307 20588 23316
rect 20536 23273 20545 23307
rect 20545 23273 20579 23307
rect 20579 23273 20588 23307
rect 20536 23264 20588 23273
rect 28172 23264 28224 23316
rect 28264 23307 28316 23316
rect 28264 23273 28273 23307
rect 28273 23273 28307 23307
rect 28307 23273 28316 23307
rect 28264 23264 28316 23273
rect 31576 23264 31628 23316
rect 32128 23307 32180 23316
rect 32128 23273 32137 23307
rect 32137 23273 32171 23307
rect 32171 23273 32180 23307
rect 32128 23264 32180 23273
rect 33048 23264 33100 23316
rect 36268 23264 36320 23316
rect 36912 23307 36964 23316
rect 36912 23273 36921 23307
rect 36921 23273 36955 23307
rect 36955 23273 36964 23307
rect 36912 23264 36964 23273
rect 37280 23264 37332 23316
rect 10232 23128 10284 23180
rect 10508 23128 10560 23180
rect 21916 23196 21968 23248
rect 23204 23196 23256 23248
rect 16028 23060 16080 23112
rect 17684 23128 17736 23180
rect 18788 23128 18840 23180
rect 18880 23103 18932 23112
rect 18880 23069 18889 23103
rect 18889 23069 18923 23103
rect 18923 23069 18932 23103
rect 18880 23060 18932 23069
rect 19340 23103 19392 23112
rect 19340 23069 19349 23103
rect 19349 23069 19383 23103
rect 19383 23069 19392 23103
rect 19340 23060 19392 23069
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 9220 23035 9272 23044
rect 9220 23001 9229 23035
rect 9229 23001 9263 23035
rect 9263 23001 9272 23035
rect 9220 22992 9272 23001
rect 9680 22992 9732 23044
rect 16580 22992 16632 23044
rect 19984 23103 20036 23112
rect 19984 23069 19993 23103
rect 19993 23069 20027 23103
rect 20027 23069 20036 23103
rect 19984 23060 20036 23069
rect 20076 23060 20128 23112
rect 20812 23128 20864 23180
rect 22836 23171 22888 23180
rect 21088 23103 21140 23112
rect 21088 23069 21097 23103
rect 21097 23069 21131 23103
rect 21131 23069 21140 23103
rect 21088 23060 21140 23069
rect 20996 23035 21048 23044
rect 20996 23001 21005 23035
rect 21005 23001 21039 23035
rect 21039 23001 21048 23035
rect 20996 22992 21048 23001
rect 22836 23137 22845 23171
rect 22845 23137 22879 23171
rect 22879 23137 22888 23171
rect 22836 23128 22888 23137
rect 24400 23171 24452 23180
rect 24400 23137 24409 23171
rect 24409 23137 24443 23171
rect 24443 23137 24452 23171
rect 24400 23128 24452 23137
rect 26240 23128 26292 23180
rect 23940 23103 23992 23112
rect 23940 23069 23949 23103
rect 23949 23069 23983 23103
rect 23983 23069 23992 23103
rect 23940 23060 23992 23069
rect 24308 23060 24360 23112
rect 26424 23103 26476 23112
rect 26424 23069 26433 23103
rect 26433 23069 26467 23103
rect 26467 23069 26476 23103
rect 26424 23060 26476 23069
rect 26608 23060 26660 23112
rect 26792 23060 26844 23112
rect 27896 23196 27948 23248
rect 30104 23239 30156 23248
rect 30104 23205 30113 23239
rect 30113 23205 30147 23239
rect 30147 23205 30156 23239
rect 30104 23196 30156 23205
rect 37464 23196 37516 23248
rect 24952 22992 25004 23044
rect 25412 22992 25464 23044
rect 2320 22924 2372 22976
rect 3148 22924 3200 22976
rect 4068 22924 4120 22976
rect 5172 22924 5224 22976
rect 5632 22967 5684 22976
rect 5632 22933 5641 22967
rect 5641 22933 5675 22967
rect 5675 22933 5684 22967
rect 5632 22924 5684 22933
rect 5724 22924 5776 22976
rect 7012 22924 7064 22976
rect 8576 22924 8628 22976
rect 8668 22924 8720 22976
rect 12072 22967 12124 22976
rect 12072 22933 12081 22967
rect 12081 22933 12115 22967
rect 12115 22933 12124 22967
rect 12072 22924 12124 22933
rect 15752 22967 15804 22976
rect 15752 22933 15761 22967
rect 15761 22933 15795 22967
rect 15795 22933 15804 22967
rect 15752 22924 15804 22933
rect 16120 22967 16172 22976
rect 16120 22933 16129 22967
rect 16129 22933 16163 22967
rect 16163 22933 16172 22967
rect 16120 22924 16172 22933
rect 18144 22924 18196 22976
rect 19248 22924 19300 22976
rect 24492 22924 24544 22976
rect 27252 23060 27304 23112
rect 30288 23128 30340 23180
rect 27804 23103 27856 23112
rect 27804 23069 27813 23103
rect 27813 23069 27847 23103
rect 27847 23069 27856 23103
rect 27804 23060 27856 23069
rect 27896 23103 27948 23112
rect 27896 23069 27905 23103
rect 27905 23069 27939 23103
rect 27939 23069 27948 23103
rect 27896 23060 27948 23069
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 28448 23103 28500 23112
rect 28448 23069 28457 23103
rect 28457 23069 28491 23103
rect 28491 23069 28500 23103
rect 28448 23060 28500 23069
rect 28540 23103 28592 23112
rect 28540 23069 28549 23103
rect 28549 23069 28583 23103
rect 28583 23069 28592 23103
rect 28540 23060 28592 23069
rect 30840 23060 30892 23112
rect 36636 23128 36688 23180
rect 31760 23103 31812 23112
rect 31760 23069 31769 23103
rect 31769 23069 31803 23103
rect 31803 23069 31812 23103
rect 31760 23060 31812 23069
rect 32128 23103 32180 23112
rect 32128 23069 32137 23103
rect 32137 23069 32171 23103
rect 32171 23069 32180 23103
rect 32128 23060 32180 23069
rect 33140 23103 33192 23112
rect 33140 23069 33149 23103
rect 33149 23069 33183 23103
rect 33183 23069 33192 23103
rect 33140 23060 33192 23069
rect 33232 23103 33284 23112
rect 33232 23069 33241 23103
rect 33241 23069 33275 23103
rect 33275 23069 33284 23103
rect 33232 23060 33284 23069
rect 36728 23103 36780 23112
rect 36728 23069 36737 23103
rect 36737 23069 36771 23103
rect 36771 23069 36780 23103
rect 36728 23060 36780 23069
rect 36912 23103 36964 23112
rect 36912 23069 36921 23103
rect 36921 23069 36955 23103
rect 36955 23069 36964 23103
rect 36912 23060 36964 23069
rect 37188 23103 37240 23112
rect 37188 23069 37197 23103
rect 37197 23069 37231 23103
rect 37231 23069 37240 23103
rect 37188 23060 37240 23069
rect 37372 23060 37424 23112
rect 37648 23060 37700 23112
rect 37924 23103 37976 23112
rect 37924 23069 37933 23103
rect 37933 23069 37967 23103
rect 37967 23069 37976 23103
rect 37924 23060 37976 23069
rect 37372 22924 37424 22976
rect 38108 22924 38160 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 5632 22720 5684 22772
rect 2320 22695 2372 22704
rect 2320 22661 2329 22695
rect 2329 22661 2363 22695
rect 2363 22661 2372 22695
rect 2320 22652 2372 22661
rect 3056 22652 3108 22704
rect 4068 22652 4120 22704
rect 1400 22516 1452 22568
rect 2044 22559 2096 22568
rect 2044 22525 2053 22559
rect 2053 22525 2087 22559
rect 2087 22525 2096 22559
rect 3884 22559 3936 22568
rect 2044 22516 2096 22525
rect 3884 22525 3893 22559
rect 3893 22525 3927 22559
rect 3927 22525 3936 22559
rect 3884 22516 3936 22525
rect 4712 22516 4764 22568
rect 4804 22516 4856 22568
rect 5908 22584 5960 22636
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 6644 22652 6696 22704
rect 6828 22720 6880 22772
rect 8392 22720 8444 22772
rect 8760 22720 8812 22772
rect 9220 22720 9272 22772
rect 11796 22720 11848 22772
rect 7012 22695 7064 22704
rect 7012 22661 7021 22695
rect 7021 22661 7055 22695
rect 7055 22661 7064 22695
rect 7012 22652 7064 22661
rect 8024 22652 8076 22704
rect 8668 22695 8720 22704
rect 8668 22661 8677 22695
rect 8677 22661 8711 22695
rect 8711 22661 8720 22695
rect 8668 22652 8720 22661
rect 14556 22720 14608 22772
rect 19616 22720 19668 22772
rect 19984 22720 20036 22772
rect 18788 22652 18840 22704
rect 20996 22763 21048 22772
rect 20996 22729 21005 22763
rect 21005 22729 21039 22763
rect 21039 22729 21048 22763
rect 20996 22720 21048 22729
rect 22284 22720 22336 22772
rect 25504 22720 25556 22772
rect 26792 22763 26844 22772
rect 26792 22729 26801 22763
rect 26801 22729 26835 22763
rect 26835 22729 26844 22763
rect 26792 22720 26844 22729
rect 27712 22720 27764 22772
rect 28816 22720 28868 22772
rect 29368 22720 29420 22772
rect 30196 22763 30248 22772
rect 30196 22729 30205 22763
rect 30205 22729 30239 22763
rect 30239 22729 30248 22763
rect 30196 22720 30248 22729
rect 30288 22763 30340 22772
rect 30288 22729 30297 22763
rect 30297 22729 30331 22763
rect 30331 22729 30340 22763
rect 30288 22720 30340 22729
rect 30840 22763 30892 22772
rect 30840 22729 30849 22763
rect 30849 22729 30883 22763
rect 30883 22729 30892 22763
rect 30840 22720 30892 22729
rect 32128 22763 32180 22772
rect 32128 22729 32137 22763
rect 32137 22729 32171 22763
rect 32171 22729 32180 22763
rect 32128 22720 32180 22729
rect 33232 22720 33284 22772
rect 11336 22584 11388 22636
rect 12072 22584 12124 22636
rect 19156 22584 19208 22636
rect 21364 22652 21416 22704
rect 5724 22559 5776 22568
rect 5724 22525 5733 22559
rect 5733 22525 5767 22559
rect 5767 22525 5776 22559
rect 5724 22516 5776 22525
rect 7472 22516 7524 22568
rect 13728 22516 13780 22568
rect 20260 22584 20312 22636
rect 23204 22695 23256 22704
rect 23204 22661 23213 22695
rect 23213 22661 23247 22695
rect 23247 22661 23256 22695
rect 23204 22652 23256 22661
rect 23664 22652 23716 22704
rect 24768 22652 24820 22704
rect 18696 22448 18748 22500
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 3976 22380 4028 22432
rect 5356 22380 5408 22432
rect 5908 22380 5960 22432
rect 9588 22380 9640 22432
rect 12992 22380 13044 22432
rect 19340 22380 19392 22432
rect 21180 22423 21232 22432
rect 21180 22389 21189 22423
rect 21189 22389 21223 22423
rect 21223 22389 21232 22423
rect 22928 22559 22980 22568
rect 22928 22525 22937 22559
rect 22937 22525 22971 22559
rect 22971 22525 22980 22559
rect 22928 22516 22980 22525
rect 26424 22516 26476 22568
rect 26608 22627 26660 22636
rect 26608 22593 26617 22627
rect 26617 22593 26651 22627
rect 26651 22593 26660 22627
rect 26608 22584 26660 22593
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 28540 22652 28592 22704
rect 26700 22516 26752 22568
rect 27344 22559 27396 22568
rect 27344 22525 27353 22559
rect 27353 22525 27387 22559
rect 27387 22525 27396 22559
rect 27344 22516 27396 22525
rect 27712 22516 27764 22568
rect 28080 22559 28132 22568
rect 28080 22525 28089 22559
rect 28089 22525 28123 22559
rect 28123 22525 28132 22559
rect 28080 22516 28132 22525
rect 28632 22627 28684 22636
rect 28632 22593 28641 22627
rect 28641 22593 28675 22627
rect 28675 22593 28684 22627
rect 28632 22584 28684 22593
rect 28908 22584 28960 22636
rect 29184 22695 29236 22704
rect 29184 22661 29193 22695
rect 29193 22661 29227 22695
rect 29227 22661 29236 22695
rect 29184 22652 29236 22661
rect 29000 22516 29052 22568
rect 30380 22584 30432 22636
rect 21180 22380 21232 22389
rect 22652 22448 22704 22500
rect 26884 22448 26936 22500
rect 27436 22448 27488 22500
rect 22376 22380 22428 22432
rect 23664 22380 23716 22432
rect 24308 22380 24360 22432
rect 26976 22380 27028 22432
rect 27344 22423 27396 22432
rect 27344 22389 27353 22423
rect 27353 22389 27387 22423
rect 27387 22389 27396 22423
rect 27344 22380 27396 22389
rect 28816 22448 28868 22500
rect 30104 22516 30156 22568
rect 32036 22516 32088 22568
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 33048 22652 33100 22704
rect 32864 22584 32916 22636
rect 34336 22720 34388 22772
rect 34612 22720 34664 22772
rect 34796 22763 34848 22772
rect 34796 22729 34805 22763
rect 34805 22729 34839 22763
rect 34839 22729 34848 22763
rect 34796 22720 34848 22729
rect 36636 22720 36688 22772
rect 36728 22720 36780 22772
rect 37832 22763 37884 22772
rect 37832 22729 37841 22763
rect 37841 22729 37875 22763
rect 37875 22729 37884 22763
rect 37832 22720 37884 22729
rect 37924 22763 37976 22772
rect 37924 22729 37933 22763
rect 37933 22729 37967 22763
rect 37967 22729 37976 22763
rect 37924 22720 37976 22729
rect 34428 22627 34480 22636
rect 34428 22593 34437 22627
rect 34437 22593 34471 22627
rect 34471 22593 34480 22627
rect 34428 22584 34480 22593
rect 34612 22627 34664 22636
rect 34612 22593 34621 22627
rect 34621 22593 34655 22627
rect 34655 22593 34664 22627
rect 34612 22584 34664 22593
rect 35348 22627 35400 22636
rect 35348 22593 35357 22627
rect 35357 22593 35391 22627
rect 35391 22593 35400 22627
rect 35348 22584 35400 22593
rect 35900 22584 35952 22636
rect 37280 22652 37332 22704
rect 31760 22448 31812 22500
rect 33968 22516 34020 22568
rect 35440 22448 35492 22500
rect 36452 22627 36504 22636
rect 36452 22593 36461 22627
rect 36461 22593 36495 22627
rect 36495 22593 36504 22627
rect 36452 22584 36504 22593
rect 36636 22584 36688 22636
rect 37556 22584 37608 22636
rect 37464 22516 37516 22568
rect 36636 22448 36688 22500
rect 38016 22652 38068 22704
rect 38384 22652 38436 22704
rect 29184 22380 29236 22432
rect 32864 22380 32916 22432
rect 35348 22380 35400 22432
rect 38108 22423 38160 22432
rect 38108 22389 38117 22423
rect 38117 22389 38151 22423
rect 38151 22389 38160 22423
rect 38108 22380 38160 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5172 22176 5224 22228
rect 5448 22176 5500 22228
rect 5908 22219 5960 22228
rect 3884 22040 3936 22092
rect 4620 22040 4672 22092
rect 5908 22185 5938 22219
rect 5938 22185 5960 22219
rect 5908 22176 5960 22185
rect 7472 22176 7524 22228
rect 14280 22176 14332 22228
rect 14556 22176 14608 22228
rect 15108 22176 15160 22228
rect 15752 22176 15804 22228
rect 20444 22176 20496 22228
rect 26976 22176 27028 22228
rect 27436 22176 27488 22228
rect 28080 22176 28132 22228
rect 28632 22219 28684 22228
rect 28632 22185 28641 22219
rect 28641 22185 28675 22219
rect 28675 22185 28684 22219
rect 28632 22176 28684 22185
rect 30104 22219 30156 22228
rect 30104 22185 30113 22219
rect 30113 22185 30147 22219
rect 30147 22185 30156 22219
rect 30104 22176 30156 22185
rect 32036 22219 32088 22228
rect 32036 22185 32045 22219
rect 32045 22185 32079 22219
rect 32079 22185 32088 22219
rect 32036 22176 32088 22185
rect 32312 22176 32364 22228
rect 33140 22176 33192 22228
rect 34428 22219 34480 22228
rect 34428 22185 34437 22219
rect 34437 22185 34471 22219
rect 34471 22185 34480 22219
rect 34428 22176 34480 22185
rect 34612 22176 34664 22228
rect 36452 22176 36504 22228
rect 37556 22176 37608 22228
rect 8852 22108 8904 22160
rect 20904 22108 20956 22160
rect 21640 22108 21692 22160
rect 3792 21972 3844 22024
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 8484 22040 8536 22092
rect 9956 22040 10008 22092
rect 11244 22040 11296 22092
rect 11704 22040 11756 22092
rect 12532 22040 12584 22092
rect 5632 22015 5684 22024
rect 5632 21981 5641 22015
rect 5641 21981 5675 22015
rect 5675 21981 5684 22015
rect 5632 21972 5684 21981
rect 9036 21972 9088 22024
rect 13728 22040 13780 22092
rect 16120 22040 16172 22092
rect 19248 22040 19300 22092
rect 20812 22040 20864 22092
rect 22928 22040 22980 22092
rect 27896 22040 27948 22092
rect 14188 21972 14240 22024
rect 17408 21972 17460 22024
rect 20076 22015 20128 22024
rect 20076 21981 20080 22015
rect 20080 21981 20114 22015
rect 20114 21981 20128 22015
rect 20076 21972 20128 21981
rect 2872 21879 2924 21888
rect 2872 21845 2881 21879
rect 2881 21845 2915 21879
rect 2915 21845 2924 21879
rect 2872 21836 2924 21845
rect 3700 21836 3752 21888
rect 3976 21836 4028 21888
rect 9680 21904 9732 21956
rect 11244 21904 11296 21956
rect 11796 21947 11848 21956
rect 11796 21913 11805 21947
rect 11805 21913 11839 21947
rect 11839 21913 11848 21947
rect 11796 21904 11848 21913
rect 12440 21947 12492 21956
rect 12440 21913 12449 21947
rect 12449 21913 12483 21947
rect 12483 21913 12492 21947
rect 12440 21904 12492 21913
rect 11060 21836 11112 21888
rect 11704 21836 11756 21888
rect 16672 21904 16724 21956
rect 18696 21947 18748 21956
rect 18696 21913 18705 21947
rect 18705 21913 18739 21947
rect 18739 21913 18748 21947
rect 18696 21904 18748 21913
rect 20628 21972 20680 22024
rect 20996 21972 21048 22024
rect 21364 22015 21416 22024
rect 21364 21981 21381 22015
rect 21381 21981 21416 22015
rect 21364 21972 21416 21981
rect 21640 22015 21692 22024
rect 21640 21981 21649 22015
rect 21649 21981 21683 22015
rect 21683 21981 21692 22015
rect 21640 21972 21692 21981
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 26608 21972 26660 22024
rect 28816 22040 28868 22092
rect 30196 22040 30248 22092
rect 35256 22040 35308 22092
rect 37280 22083 37332 22092
rect 37280 22049 37289 22083
rect 37289 22049 37323 22083
rect 37323 22049 37332 22083
rect 37280 22040 37332 22049
rect 18052 21836 18104 21888
rect 19892 21879 19944 21888
rect 19892 21845 19901 21879
rect 19901 21845 19935 21879
rect 19935 21845 19944 21879
rect 19892 21836 19944 21845
rect 20076 21836 20128 21888
rect 20720 21904 20772 21956
rect 21456 21947 21508 21956
rect 21456 21913 21465 21947
rect 21465 21913 21499 21947
rect 21499 21913 21508 21947
rect 21456 21904 21508 21913
rect 22100 21904 22152 21956
rect 20904 21836 20956 21888
rect 21824 21836 21876 21888
rect 24308 21904 24360 21956
rect 25872 21904 25924 21956
rect 28448 22015 28500 22024
rect 28448 21981 28457 22015
rect 28457 21981 28491 22015
rect 28491 21981 28500 22015
rect 28448 21972 28500 21981
rect 28632 22015 28684 22024
rect 28632 21981 28641 22015
rect 28641 21981 28675 22015
rect 28675 21981 28684 22015
rect 28632 21972 28684 21981
rect 29644 21972 29696 22024
rect 28816 21904 28868 21956
rect 29460 21904 29512 21956
rect 32680 22015 32732 22024
rect 32680 21981 32689 22015
rect 32689 21981 32723 22015
rect 32723 21981 32732 22015
rect 32680 21972 32732 21981
rect 32864 22015 32916 22024
rect 32864 21981 32873 22015
rect 32873 21981 32907 22015
rect 32907 21981 32916 22015
rect 32864 21972 32916 21981
rect 34428 21972 34480 22024
rect 35348 22015 35400 22024
rect 35348 21981 35357 22015
rect 35357 21981 35391 22015
rect 35391 21981 35400 22015
rect 35348 21972 35400 21981
rect 37096 21972 37148 22024
rect 37372 22015 37424 22024
rect 37372 21981 37381 22015
rect 37381 21981 37415 22015
rect 37415 21981 37424 22015
rect 37372 21972 37424 21981
rect 33048 21947 33100 21956
rect 33048 21913 33057 21947
rect 33057 21913 33091 21947
rect 33091 21913 33100 21947
rect 33048 21904 33100 21913
rect 25780 21836 25832 21888
rect 28356 21836 28408 21888
rect 34704 21836 34756 21888
rect 37556 21904 37608 21956
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 4712 21632 4764 21684
rect 6184 21632 6236 21684
rect 8944 21632 8996 21684
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12440 21632 12492 21684
rect 13360 21632 13412 21684
rect 14096 21632 14148 21684
rect 15108 21632 15160 21684
rect 17408 21632 17460 21684
rect 18696 21632 18748 21684
rect 21732 21632 21784 21684
rect 26792 21632 26844 21684
rect 28356 21632 28408 21684
rect 28908 21632 28960 21684
rect 33968 21675 34020 21684
rect 33968 21641 33977 21675
rect 33977 21641 34011 21675
rect 34011 21641 34020 21675
rect 33968 21632 34020 21641
rect 35256 21632 35308 21684
rect 35348 21675 35400 21684
rect 35348 21641 35357 21675
rect 35357 21641 35391 21675
rect 35391 21641 35400 21675
rect 35348 21632 35400 21641
rect 3976 21607 4028 21616
rect 3976 21573 3985 21607
rect 3985 21573 4019 21607
rect 4019 21573 4028 21607
rect 3976 21564 4028 21573
rect 4620 21564 4672 21616
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 5356 21496 5408 21548
rect 5724 21539 5776 21548
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 9680 21564 9732 21616
rect 9956 21564 10008 21616
rect 12164 21607 12216 21616
rect 12164 21573 12173 21607
rect 12173 21573 12207 21607
rect 12207 21573 12216 21607
rect 12164 21564 12216 21573
rect 12992 21564 13044 21616
rect 16672 21564 16724 21616
rect 20720 21564 20772 21616
rect 6460 21496 6512 21548
rect 11612 21496 11664 21548
rect 5540 21428 5592 21480
rect 8576 21471 8628 21480
rect 8576 21437 8585 21471
rect 8585 21437 8619 21471
rect 8619 21437 8628 21471
rect 8576 21428 8628 21437
rect 10508 21471 10560 21480
rect 10508 21437 10517 21471
rect 10517 21437 10551 21471
rect 10551 21437 10560 21471
rect 10508 21428 10560 21437
rect 10600 21428 10652 21480
rect 12716 21496 12768 21548
rect 13452 21496 13504 21548
rect 13636 21539 13688 21548
rect 13636 21505 13645 21539
rect 13645 21505 13679 21539
rect 13679 21505 13688 21539
rect 13636 21496 13688 21505
rect 5448 21360 5500 21412
rect 6000 21360 6052 21412
rect 13544 21428 13596 21480
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 14188 21360 14240 21412
rect 4160 21292 4212 21344
rect 4804 21292 4856 21344
rect 7932 21292 7984 21344
rect 10692 21292 10744 21344
rect 12992 21292 13044 21344
rect 13360 21292 13412 21344
rect 14464 21471 14516 21480
rect 14464 21437 14473 21471
rect 14473 21437 14507 21471
rect 14507 21437 14516 21471
rect 14464 21428 14516 21437
rect 15200 21428 15252 21480
rect 20904 21496 20956 21548
rect 21732 21496 21784 21548
rect 21916 21496 21968 21548
rect 22376 21496 22428 21548
rect 17040 21471 17092 21480
rect 17040 21437 17049 21471
rect 17049 21437 17083 21471
rect 17083 21437 17092 21471
rect 17040 21428 17092 21437
rect 17960 21428 18012 21480
rect 18144 21428 18196 21480
rect 21640 21428 21692 21480
rect 22100 21471 22152 21480
rect 22100 21437 22109 21471
rect 22109 21437 22143 21471
rect 22143 21437 22152 21471
rect 22100 21428 22152 21437
rect 22560 21428 22612 21480
rect 21824 21360 21876 21412
rect 25964 21564 26016 21616
rect 29920 21564 29972 21616
rect 25136 21471 25188 21480
rect 25136 21437 25145 21471
rect 25145 21437 25179 21471
rect 25179 21437 25188 21471
rect 25136 21428 25188 21437
rect 25780 21539 25832 21548
rect 25780 21505 25789 21539
rect 25789 21505 25823 21539
rect 25823 21505 25832 21539
rect 25780 21496 25832 21505
rect 25872 21539 25924 21548
rect 25872 21505 25881 21539
rect 25881 21505 25915 21539
rect 25915 21505 25924 21539
rect 25872 21496 25924 21505
rect 26976 21539 27028 21548
rect 15568 21292 15620 21344
rect 20352 21335 20404 21344
rect 20352 21301 20361 21335
rect 20361 21301 20395 21335
rect 20395 21301 20404 21335
rect 20352 21292 20404 21301
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 21548 21292 21600 21344
rect 22008 21292 22060 21344
rect 22560 21335 22612 21344
rect 22560 21301 22569 21335
rect 22569 21301 22603 21335
rect 22603 21301 22612 21335
rect 22560 21292 22612 21301
rect 23848 21292 23900 21344
rect 26240 21360 26292 21412
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27804 21496 27856 21548
rect 28632 21496 28684 21548
rect 29276 21539 29328 21548
rect 29276 21505 29285 21539
rect 29285 21505 29319 21539
rect 29319 21505 29328 21539
rect 29276 21496 29328 21505
rect 29460 21539 29512 21548
rect 29460 21505 29469 21539
rect 29469 21505 29503 21539
rect 29503 21505 29512 21539
rect 29460 21496 29512 21505
rect 29644 21496 29696 21548
rect 30196 21539 30248 21548
rect 30196 21505 30205 21539
rect 30205 21505 30239 21539
rect 30239 21505 30248 21539
rect 30196 21496 30248 21505
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 33876 21539 33928 21548
rect 33876 21505 33885 21539
rect 33885 21505 33919 21539
rect 33919 21505 33928 21539
rect 33876 21496 33928 21505
rect 34336 21564 34388 21616
rect 28448 21428 28500 21480
rect 29000 21360 29052 21412
rect 31760 21428 31812 21480
rect 32680 21471 32732 21480
rect 32680 21437 32689 21471
rect 32689 21437 32723 21471
rect 32723 21437 32732 21471
rect 32680 21428 32732 21437
rect 36728 21496 36780 21548
rect 26700 21292 26752 21344
rect 27252 21292 27304 21344
rect 29184 21292 29236 21344
rect 30380 21335 30432 21344
rect 30380 21301 30389 21335
rect 30389 21301 30423 21335
rect 30423 21301 30432 21335
rect 30380 21292 30432 21301
rect 36360 21292 36412 21344
rect 38200 21292 38252 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 9404 21088 9456 21140
rect 13452 21131 13504 21140
rect 13452 21097 13461 21131
rect 13461 21097 13495 21131
rect 13495 21097 13504 21131
rect 13452 21088 13504 21097
rect 13544 21088 13596 21140
rect 13728 21088 13780 21140
rect 14188 21088 14240 21140
rect 5632 20995 5684 21004
rect 5632 20961 5641 20995
rect 5641 20961 5675 20995
rect 5675 20961 5684 20995
rect 5632 20952 5684 20961
rect 2872 20927 2924 20936
rect 2872 20893 2881 20927
rect 2881 20893 2915 20927
rect 2915 20893 2924 20927
rect 2872 20884 2924 20893
rect 3884 20884 3936 20936
rect 8484 20952 8536 21004
rect 10692 20995 10744 21004
rect 10692 20961 10701 20995
rect 10701 20961 10735 20995
rect 10735 20961 10744 20995
rect 10692 20952 10744 20961
rect 3700 20816 3752 20868
rect 4804 20816 4856 20868
rect 5356 20859 5408 20868
rect 5356 20825 5365 20859
rect 5365 20825 5399 20859
rect 5399 20825 5408 20859
rect 5356 20816 5408 20825
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 9680 20884 9732 20936
rect 10416 20927 10468 20936
rect 10416 20893 10425 20927
rect 10425 20893 10459 20927
rect 10459 20893 10468 20927
rect 10416 20884 10468 20893
rect 12164 20884 12216 20936
rect 13084 20952 13136 21004
rect 13820 21020 13872 21072
rect 14464 21088 14516 21140
rect 15936 21088 15988 21140
rect 12992 20884 13044 20936
rect 13360 20884 13412 20936
rect 15200 20995 15252 21004
rect 15200 20961 15209 20995
rect 15209 20961 15243 20995
rect 15243 20961 15252 20995
rect 15200 20952 15252 20961
rect 16672 21020 16724 21072
rect 11244 20816 11296 20868
rect 13636 20816 13688 20868
rect 13728 20816 13780 20868
rect 2780 20748 2832 20800
rect 3424 20791 3476 20800
rect 3424 20757 3433 20791
rect 3433 20757 3467 20791
rect 3467 20757 3476 20791
rect 3424 20748 3476 20757
rect 4712 20748 4764 20800
rect 7748 20791 7800 20800
rect 7748 20757 7757 20791
rect 7757 20757 7791 20791
rect 7791 20757 7800 20791
rect 7748 20748 7800 20757
rect 12164 20791 12216 20800
rect 12164 20757 12173 20791
rect 12173 20757 12207 20791
rect 12207 20757 12216 20791
rect 12164 20748 12216 20757
rect 12716 20748 12768 20800
rect 15568 20927 15620 20936
rect 15568 20893 15577 20927
rect 15577 20893 15611 20927
rect 15611 20893 15620 20927
rect 15568 20884 15620 20893
rect 16856 20952 16908 21004
rect 17132 21088 17184 21140
rect 17960 21131 18012 21140
rect 17960 21097 17969 21131
rect 17969 21097 18003 21131
rect 18003 21097 18012 21131
rect 17960 21088 18012 21097
rect 19340 21088 19392 21140
rect 20996 21131 21048 21140
rect 20996 21097 21005 21131
rect 21005 21097 21039 21131
rect 21039 21097 21048 21131
rect 20996 21088 21048 21097
rect 21732 21131 21784 21140
rect 21732 21097 21741 21131
rect 21741 21097 21775 21131
rect 21775 21097 21784 21131
rect 21732 21088 21784 21097
rect 22376 21131 22428 21140
rect 22376 21097 22385 21131
rect 22385 21097 22419 21131
rect 22419 21097 22428 21131
rect 22376 21088 22428 21097
rect 25136 21088 25188 21140
rect 26884 21088 26936 21140
rect 28172 21088 28224 21140
rect 29368 21088 29420 21140
rect 31760 21131 31812 21140
rect 31760 21097 31769 21131
rect 31769 21097 31803 21131
rect 31803 21097 31812 21131
rect 31760 21088 31812 21097
rect 33048 21088 33100 21140
rect 33876 21088 33928 21140
rect 34336 21131 34388 21140
rect 34336 21097 34345 21131
rect 34345 21097 34379 21131
rect 34379 21097 34388 21131
rect 34336 21088 34388 21097
rect 35992 21088 36044 21140
rect 36728 21131 36780 21140
rect 36728 21097 36737 21131
rect 36737 21097 36771 21131
rect 36771 21097 36780 21131
rect 36728 21088 36780 21097
rect 37556 21131 37608 21140
rect 37556 21097 37565 21131
rect 37565 21097 37599 21131
rect 37599 21097 37608 21131
rect 37556 21088 37608 21097
rect 17040 21020 17092 21072
rect 21180 21020 21232 21072
rect 22652 21020 22704 21072
rect 17868 20995 17920 21004
rect 17868 20961 17877 20995
rect 17877 20961 17911 20995
rect 17911 20961 17920 20995
rect 17868 20952 17920 20961
rect 18788 20952 18840 21004
rect 19248 20995 19300 21004
rect 19248 20961 19257 20995
rect 19257 20961 19291 20995
rect 19291 20961 19300 20995
rect 19248 20952 19300 20961
rect 21272 20952 21324 21004
rect 21456 20952 21508 21004
rect 15568 20748 15620 20800
rect 16396 20791 16448 20800
rect 16396 20757 16405 20791
rect 16405 20757 16439 20791
rect 16439 20757 16448 20791
rect 16396 20748 16448 20757
rect 16856 20791 16908 20800
rect 16856 20757 16865 20791
rect 16865 20757 16899 20791
rect 16899 20757 16908 20791
rect 16856 20748 16908 20757
rect 16948 20748 17000 20800
rect 21824 20927 21876 20936
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 24400 20995 24452 21004
rect 24400 20961 24409 20995
rect 24409 20961 24443 20995
rect 24443 20961 24452 20995
rect 24400 20952 24452 20961
rect 28080 21020 28132 21072
rect 29000 21020 29052 21072
rect 27068 20952 27120 21004
rect 22468 20884 22520 20936
rect 23020 20927 23072 20936
rect 23020 20893 23029 20927
rect 23029 20893 23063 20927
rect 23063 20893 23072 20927
rect 23020 20884 23072 20893
rect 23296 20927 23348 20936
rect 23296 20893 23305 20927
rect 23305 20893 23339 20927
rect 23339 20893 23348 20927
rect 23296 20884 23348 20893
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 26976 20884 27028 20936
rect 18236 20816 18288 20868
rect 18144 20748 18196 20800
rect 18512 20748 18564 20800
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 19524 20859 19576 20868
rect 19524 20825 19533 20859
rect 19533 20825 19567 20859
rect 19567 20825 19576 20859
rect 19524 20816 19576 20825
rect 20996 20816 21048 20868
rect 23480 20816 23532 20868
rect 25504 20816 25556 20868
rect 27804 20884 27856 20936
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 29276 21020 29328 21072
rect 28816 20927 28868 20936
rect 28816 20893 28825 20927
rect 28825 20893 28859 20927
rect 28859 20893 28868 20927
rect 28816 20884 28868 20893
rect 28908 20927 28960 20936
rect 28908 20893 28917 20927
rect 28917 20893 28951 20927
rect 28951 20893 28960 20927
rect 28908 20884 28960 20893
rect 29000 20927 29052 20936
rect 29000 20893 29009 20927
rect 29009 20893 29043 20927
rect 29043 20893 29052 20927
rect 29000 20884 29052 20893
rect 29184 20927 29236 20936
rect 29184 20893 29193 20927
rect 29193 20893 29227 20927
rect 29227 20893 29236 20927
rect 29184 20884 29236 20893
rect 29460 20884 29512 20936
rect 30380 20884 30432 20936
rect 30840 20952 30892 21004
rect 37924 21020 37976 21072
rect 31392 20927 31444 20936
rect 31392 20893 31401 20927
rect 31401 20893 31435 20927
rect 31435 20893 31444 20927
rect 31392 20884 31444 20893
rect 31576 20927 31628 20936
rect 31576 20893 31585 20927
rect 31585 20893 31619 20927
rect 31619 20893 31628 20927
rect 31576 20884 31628 20893
rect 27620 20816 27672 20868
rect 32312 20927 32364 20936
rect 32312 20893 32321 20927
rect 32321 20893 32355 20927
rect 32355 20893 32364 20927
rect 32312 20884 32364 20893
rect 33876 20927 33928 20936
rect 33876 20893 33885 20927
rect 33885 20893 33919 20927
rect 33919 20893 33928 20927
rect 33876 20884 33928 20893
rect 35440 20884 35492 20936
rect 35992 20927 36044 20936
rect 35992 20893 36001 20927
rect 36001 20893 36035 20927
rect 36035 20893 36044 20927
rect 35992 20884 36044 20893
rect 31944 20859 31996 20868
rect 31944 20825 31953 20859
rect 31953 20825 31987 20859
rect 31987 20825 31996 20859
rect 31944 20816 31996 20825
rect 32588 20816 32640 20868
rect 22192 20791 22244 20800
rect 22192 20757 22201 20791
rect 22201 20757 22235 20791
rect 22235 20757 22244 20791
rect 22192 20748 22244 20757
rect 26332 20748 26384 20800
rect 28448 20791 28500 20800
rect 28448 20757 28457 20791
rect 28457 20757 28491 20791
rect 28491 20757 28500 20791
rect 28448 20748 28500 20757
rect 30196 20791 30248 20800
rect 30196 20757 30205 20791
rect 30205 20757 30239 20791
rect 30239 20757 30248 20791
rect 30196 20748 30248 20757
rect 31576 20748 31628 20800
rect 32312 20748 32364 20800
rect 33048 20859 33100 20868
rect 33048 20825 33057 20859
rect 33057 20825 33091 20859
rect 33091 20825 33100 20859
rect 33048 20816 33100 20825
rect 35992 20748 36044 20800
rect 36544 20884 36596 20936
rect 36728 20884 36780 20936
rect 37832 20927 37884 20936
rect 37832 20893 37841 20927
rect 37841 20893 37875 20927
rect 37875 20893 37884 20927
rect 37832 20884 37884 20893
rect 38108 20927 38160 20936
rect 38108 20893 38117 20927
rect 38117 20893 38151 20927
rect 38151 20893 38160 20927
rect 38108 20884 38160 20893
rect 38200 20927 38252 20936
rect 38200 20893 38209 20927
rect 38209 20893 38243 20927
rect 38243 20893 38252 20927
rect 38200 20884 38252 20893
rect 38384 20927 38436 20936
rect 38384 20893 38393 20927
rect 38393 20893 38427 20927
rect 38427 20893 38436 20927
rect 38384 20884 38436 20893
rect 37740 20859 37792 20868
rect 37740 20825 37749 20859
rect 37749 20825 37783 20859
rect 37783 20825 37792 20859
rect 37740 20816 37792 20825
rect 36452 20748 36504 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 3424 20544 3476 20596
rect 2780 20476 2832 20528
rect 4804 20476 4856 20528
rect 5356 20587 5408 20596
rect 5356 20553 5365 20587
rect 5365 20553 5399 20587
rect 5399 20553 5408 20587
rect 5356 20544 5408 20553
rect 8576 20544 8628 20596
rect 8024 20476 8076 20528
rect 9588 20544 9640 20596
rect 11612 20587 11664 20596
rect 11612 20553 11621 20587
rect 11621 20553 11655 20587
rect 11655 20553 11664 20587
rect 11612 20544 11664 20553
rect 12164 20544 12216 20596
rect 9404 20519 9456 20528
rect 9404 20485 9413 20519
rect 9413 20485 9447 20519
rect 9447 20485 9456 20519
rect 9404 20476 9456 20485
rect 2044 20408 2096 20460
rect 5540 20451 5592 20460
rect 5540 20417 5549 20451
rect 5549 20417 5583 20451
rect 5583 20417 5592 20451
rect 5540 20408 5592 20417
rect 3700 20204 3752 20256
rect 4712 20340 4764 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 3884 20272 3936 20324
rect 7748 20451 7800 20460
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 12900 20544 12952 20596
rect 13728 20544 13780 20596
rect 16856 20544 16908 20596
rect 17500 20544 17552 20596
rect 18236 20544 18288 20596
rect 19524 20544 19576 20596
rect 25872 20544 25924 20596
rect 25964 20587 26016 20596
rect 25964 20553 25973 20587
rect 25973 20553 26007 20587
rect 26007 20553 26016 20587
rect 25964 20544 26016 20553
rect 26608 20544 26660 20596
rect 27528 20544 27580 20596
rect 34428 20587 34480 20596
rect 34428 20553 34437 20587
rect 34437 20553 34471 20587
rect 34471 20553 34480 20587
rect 34428 20544 34480 20553
rect 35440 20544 35492 20596
rect 36176 20544 36228 20596
rect 37832 20587 37884 20596
rect 37832 20553 37841 20587
rect 37841 20553 37875 20587
rect 37875 20553 37884 20587
rect 37832 20544 37884 20553
rect 12532 20408 12584 20460
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 7472 20340 7524 20392
rect 7656 20340 7708 20392
rect 4068 20247 4120 20256
rect 4068 20213 4077 20247
rect 4077 20213 4111 20247
rect 4111 20213 4120 20247
rect 4068 20204 4120 20213
rect 4988 20247 5040 20256
rect 4988 20213 4997 20247
rect 4997 20213 5031 20247
rect 5031 20213 5040 20247
rect 4988 20204 5040 20213
rect 6644 20204 6696 20256
rect 13452 20204 13504 20256
rect 13912 20383 13964 20392
rect 13912 20349 13921 20383
rect 13921 20349 13955 20383
rect 13955 20349 13964 20383
rect 13912 20340 13964 20349
rect 15660 20340 15712 20392
rect 16580 20408 16632 20460
rect 17316 20340 17368 20392
rect 17960 20476 18012 20528
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 18880 20408 18932 20460
rect 19248 20476 19300 20528
rect 20352 20476 20404 20528
rect 21180 20519 21232 20528
rect 21180 20485 21189 20519
rect 21189 20485 21223 20519
rect 21223 20485 21232 20519
rect 21180 20476 21232 20485
rect 21548 20476 21600 20528
rect 20996 20408 21048 20460
rect 18144 20315 18196 20324
rect 18144 20281 18153 20315
rect 18153 20281 18187 20315
rect 18187 20281 18196 20315
rect 18144 20272 18196 20281
rect 18788 20272 18840 20324
rect 14372 20204 14424 20256
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 17408 20247 17460 20256
rect 17408 20213 17417 20247
rect 17417 20213 17451 20247
rect 17451 20213 17460 20247
rect 17408 20204 17460 20213
rect 19800 20340 19852 20392
rect 20076 20340 20128 20392
rect 21548 20340 21600 20392
rect 21916 20383 21968 20392
rect 21916 20349 21925 20383
rect 21925 20349 21959 20383
rect 21959 20349 21968 20383
rect 21916 20340 21968 20349
rect 22284 20340 22336 20392
rect 23848 20519 23900 20528
rect 23848 20485 23857 20519
rect 23857 20485 23891 20519
rect 23891 20485 23900 20519
rect 23848 20476 23900 20485
rect 24308 20476 24360 20528
rect 25504 20519 25556 20528
rect 25504 20485 25513 20519
rect 25513 20485 25547 20519
rect 25547 20485 25556 20519
rect 25504 20476 25556 20485
rect 22652 20408 22704 20460
rect 21640 20315 21692 20324
rect 21640 20281 21649 20315
rect 21649 20281 21683 20315
rect 21683 20281 21692 20315
rect 21640 20272 21692 20281
rect 23020 20340 23072 20392
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 23480 20451 23532 20460
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 23480 20408 23532 20417
rect 26240 20408 26292 20460
rect 26332 20451 26384 20460
rect 26332 20417 26341 20451
rect 26341 20417 26375 20451
rect 26375 20417 26384 20451
rect 26332 20408 26384 20417
rect 29276 20476 29328 20528
rect 31852 20476 31904 20528
rect 33048 20476 33100 20528
rect 36084 20476 36136 20528
rect 23388 20383 23440 20392
rect 23388 20349 23397 20383
rect 23397 20349 23431 20383
rect 23431 20349 23440 20383
rect 23388 20340 23440 20349
rect 19340 20204 19392 20256
rect 19524 20204 19576 20256
rect 21916 20204 21968 20256
rect 22376 20204 22428 20256
rect 22560 20247 22612 20256
rect 22560 20213 22569 20247
rect 22569 20213 22603 20247
rect 22603 20213 22612 20247
rect 22560 20204 22612 20213
rect 22744 20247 22796 20256
rect 22744 20213 22753 20247
rect 22753 20213 22787 20247
rect 22787 20213 22796 20247
rect 22744 20204 22796 20213
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 26056 20340 26108 20392
rect 27252 20451 27304 20460
rect 27252 20417 27261 20451
rect 27261 20417 27295 20451
rect 27295 20417 27304 20451
rect 27252 20408 27304 20417
rect 27620 20408 27672 20460
rect 29000 20408 29052 20460
rect 29368 20408 29420 20460
rect 29552 20408 29604 20460
rect 27804 20340 27856 20392
rect 28356 20340 28408 20392
rect 29736 20340 29788 20392
rect 31944 20408 31996 20460
rect 33600 20383 33652 20392
rect 33600 20349 33609 20383
rect 33609 20349 33643 20383
rect 33643 20349 33652 20383
rect 33600 20340 33652 20349
rect 33968 20451 34020 20460
rect 33968 20417 33977 20451
rect 33977 20417 34011 20451
rect 34011 20417 34020 20451
rect 33968 20408 34020 20417
rect 33876 20383 33928 20392
rect 33876 20349 33885 20383
rect 33885 20349 33919 20383
rect 33919 20349 33928 20383
rect 33876 20340 33928 20349
rect 34152 20408 34204 20460
rect 33692 20272 33744 20324
rect 35808 20383 35860 20392
rect 35808 20349 35817 20383
rect 35817 20349 35851 20383
rect 35851 20349 35860 20383
rect 35808 20340 35860 20349
rect 36176 20408 36228 20460
rect 37464 20519 37516 20528
rect 37464 20485 37473 20519
rect 37473 20485 37507 20519
rect 37507 20485 37516 20519
rect 37464 20476 37516 20485
rect 37648 20519 37700 20528
rect 37648 20485 37657 20519
rect 37657 20485 37691 20519
rect 37691 20485 37700 20519
rect 37648 20476 37700 20485
rect 35992 20340 36044 20392
rect 36360 20272 36412 20324
rect 24952 20204 25004 20256
rect 26792 20247 26844 20256
rect 26792 20213 26801 20247
rect 26801 20213 26835 20247
rect 26835 20213 26844 20247
rect 26792 20204 26844 20213
rect 29644 20204 29696 20256
rect 30104 20204 30156 20256
rect 31576 20247 31628 20256
rect 31576 20213 31585 20247
rect 31585 20213 31619 20247
rect 31619 20213 31628 20247
rect 31576 20204 31628 20213
rect 35900 20247 35952 20256
rect 35900 20213 35909 20247
rect 35909 20213 35943 20247
rect 35943 20213 35952 20247
rect 35900 20204 35952 20213
rect 35992 20247 36044 20256
rect 35992 20213 36001 20247
rect 36001 20213 36035 20247
rect 36035 20213 36044 20247
rect 35992 20204 36044 20213
rect 36728 20247 36780 20256
rect 36728 20213 36737 20247
rect 36737 20213 36771 20247
rect 36771 20213 36780 20247
rect 36728 20204 36780 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3700 20000 3752 20052
rect 3792 20043 3844 20052
rect 3792 20009 3801 20043
rect 3801 20009 3835 20043
rect 3835 20009 3844 20043
rect 3792 20000 3844 20009
rect 5540 20000 5592 20052
rect 7748 20000 7800 20052
rect 8484 20000 8536 20052
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 3884 19932 3936 19984
rect 2044 19864 2096 19916
rect 5632 19864 5684 19916
rect 6644 19907 6696 19916
rect 6644 19873 6653 19907
rect 6653 19873 6687 19907
rect 6687 19873 6696 19907
rect 6644 19864 6696 19873
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 12532 19907 12584 19916
rect 12532 19873 12541 19907
rect 12541 19873 12575 19907
rect 12575 19873 12584 19907
rect 12532 19864 12584 19873
rect 13452 19907 13504 19916
rect 13452 19873 13461 19907
rect 13461 19873 13495 19907
rect 13495 19873 13504 19907
rect 13452 19864 13504 19873
rect 14096 19932 14148 19984
rect 16672 20000 16724 20052
rect 17960 20000 18012 20052
rect 19800 20043 19852 20052
rect 19800 20009 19809 20043
rect 19809 20009 19843 20043
rect 19843 20009 19852 20043
rect 19800 20000 19852 20009
rect 21456 20000 21508 20052
rect 21732 20043 21784 20052
rect 21732 20009 21741 20043
rect 21741 20009 21775 20043
rect 21775 20009 21784 20043
rect 21732 20000 21784 20009
rect 15660 19864 15712 19916
rect 16396 19864 16448 19916
rect 18604 19864 18656 19916
rect 2780 19796 2832 19848
rect 3976 19839 4028 19848
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 4712 19796 4764 19848
rect 8576 19796 8628 19848
rect 1676 19771 1728 19780
rect 1676 19737 1685 19771
rect 1685 19737 1719 19771
rect 1719 19737 1728 19771
rect 1676 19728 1728 19737
rect 3516 19728 3568 19780
rect 3884 19728 3936 19780
rect 4988 19728 5040 19780
rect 6000 19771 6052 19780
rect 6000 19737 6009 19771
rect 6009 19737 6043 19771
rect 6043 19737 6052 19771
rect 6000 19728 6052 19737
rect 7932 19728 7984 19780
rect 11796 19728 11848 19780
rect 12256 19771 12308 19780
rect 12256 19737 12265 19771
rect 12265 19737 12299 19771
rect 12299 19737 12308 19771
rect 12256 19728 12308 19737
rect 14648 19796 14700 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 17500 19728 17552 19780
rect 17684 19728 17736 19780
rect 18696 19796 18748 19848
rect 21640 19864 21692 19916
rect 23388 20000 23440 20052
rect 28080 20043 28132 20052
rect 28080 20009 28089 20043
rect 28089 20009 28123 20043
rect 28123 20009 28132 20043
rect 28080 20000 28132 20009
rect 29184 20043 29236 20052
rect 29184 20009 29193 20043
rect 29193 20009 29227 20043
rect 29227 20009 29236 20043
rect 29184 20000 29236 20009
rect 29644 20000 29696 20052
rect 23664 19932 23716 19984
rect 29828 19932 29880 19984
rect 31852 19932 31904 19984
rect 33600 19975 33652 19984
rect 33600 19941 33609 19975
rect 33609 19941 33643 19975
rect 33643 19941 33652 19975
rect 33600 19932 33652 19941
rect 33968 19932 34020 19984
rect 35808 19932 35860 19984
rect 23480 19864 23532 19916
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 18880 19728 18932 19780
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 22744 19796 22796 19848
rect 22928 19796 22980 19848
rect 23204 19796 23256 19848
rect 24032 19796 24084 19848
rect 29368 19907 29420 19916
rect 29368 19873 29377 19907
rect 29377 19873 29411 19907
rect 29411 19873 29420 19907
rect 29368 19864 29420 19873
rect 29552 19907 29604 19916
rect 29552 19873 29561 19907
rect 29561 19873 29595 19907
rect 29595 19873 29604 19907
rect 29552 19864 29604 19873
rect 30012 19907 30064 19916
rect 30012 19873 30021 19907
rect 30021 19873 30055 19907
rect 30055 19873 30064 19907
rect 30012 19864 30064 19873
rect 30196 19864 30248 19916
rect 26056 19839 26108 19848
rect 26056 19805 26065 19839
rect 26065 19805 26099 19839
rect 26099 19805 26108 19839
rect 26056 19796 26108 19805
rect 26240 19839 26292 19848
rect 26240 19805 26249 19839
rect 26249 19805 26283 19839
rect 26283 19805 26292 19839
rect 26240 19796 26292 19805
rect 26332 19839 26384 19848
rect 26332 19805 26341 19839
rect 26341 19805 26375 19839
rect 26375 19805 26384 19839
rect 26332 19796 26384 19805
rect 27620 19796 27672 19848
rect 27804 19839 27856 19848
rect 27804 19805 27813 19839
rect 27813 19805 27847 19839
rect 27847 19805 27856 19839
rect 27804 19796 27856 19805
rect 22192 19728 22244 19780
rect 3424 19703 3476 19712
rect 3424 19669 3451 19703
rect 3451 19669 3476 19703
rect 3424 19660 3476 19669
rect 4712 19660 4764 19712
rect 5264 19660 5316 19712
rect 7472 19660 7524 19712
rect 9772 19660 9824 19712
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 11888 19660 11940 19712
rect 12440 19660 12492 19712
rect 14004 19660 14056 19712
rect 14740 19660 14792 19712
rect 18788 19660 18840 19712
rect 21456 19660 21508 19712
rect 23940 19728 23992 19780
rect 27712 19771 27764 19780
rect 27712 19737 27721 19771
rect 27721 19737 27755 19771
rect 27755 19737 27764 19771
rect 27712 19728 27764 19737
rect 28816 19839 28868 19848
rect 28816 19805 28825 19839
rect 28825 19805 28859 19839
rect 28859 19805 28868 19839
rect 28816 19796 28868 19805
rect 29000 19796 29052 19848
rect 29644 19796 29696 19848
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 29828 19796 29880 19848
rect 29460 19728 29512 19780
rect 31208 19728 31260 19780
rect 31576 19796 31628 19848
rect 32588 19839 32640 19848
rect 32588 19805 32591 19839
rect 32591 19805 32625 19839
rect 32625 19805 32640 19839
rect 32588 19796 32640 19805
rect 32680 19796 32732 19848
rect 35992 19907 36044 19916
rect 35992 19873 36001 19907
rect 36001 19873 36035 19907
rect 36035 19873 36044 19907
rect 35992 19864 36044 19873
rect 34152 19796 34204 19848
rect 35900 19796 35952 19848
rect 32128 19728 32180 19780
rect 32312 19728 32364 19780
rect 34336 19728 34388 19780
rect 36084 19728 36136 19780
rect 36268 19839 36320 19848
rect 36268 19805 36277 19839
rect 36277 19805 36311 19839
rect 36311 19805 36320 19839
rect 36268 19796 36320 19805
rect 36452 20043 36504 20052
rect 36452 20009 36461 20043
rect 36461 20009 36495 20043
rect 36495 20009 36504 20043
rect 36452 20000 36504 20009
rect 36728 20000 36780 20052
rect 36544 19864 36596 19916
rect 37924 19864 37976 19916
rect 36452 19728 36504 19780
rect 23204 19660 23256 19712
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 26884 19660 26936 19712
rect 27160 19660 27212 19712
rect 27988 19660 28040 19712
rect 29552 19660 29604 19712
rect 29920 19703 29972 19712
rect 29920 19669 29929 19703
rect 29929 19669 29963 19703
rect 29963 19669 29972 19703
rect 29920 19660 29972 19669
rect 33232 19660 33284 19712
rect 33784 19660 33836 19712
rect 35440 19660 35492 19712
rect 36176 19660 36228 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 112 19388 164 19440
rect 2872 19388 2924 19440
rect 3424 19363 3476 19372
rect 1676 19252 1728 19304
rect 3424 19329 3433 19363
rect 3433 19329 3467 19363
rect 3467 19329 3476 19363
rect 3424 19320 3476 19329
rect 3516 19363 3568 19372
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 4068 19388 4120 19440
rect 7932 19388 7984 19440
rect 5724 19320 5776 19372
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 8484 19320 8536 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12256 19320 12308 19372
rect 12992 19388 13044 19440
rect 5264 19295 5316 19304
rect 5264 19261 5273 19295
rect 5273 19261 5307 19295
rect 5307 19261 5316 19295
rect 5264 19252 5316 19261
rect 9220 19252 9272 19304
rect 9772 19295 9824 19304
rect 9772 19261 9781 19295
rect 9781 19261 9815 19295
rect 9815 19261 9824 19295
rect 9772 19252 9824 19261
rect 10324 19252 10376 19304
rect 10968 19252 11020 19304
rect 6000 19184 6052 19236
rect 10784 19184 10836 19236
rect 12900 19363 12952 19372
rect 12900 19329 12909 19363
rect 12909 19329 12943 19363
rect 12943 19329 12952 19363
rect 12900 19320 12952 19329
rect 14372 19388 14424 19440
rect 18788 19431 18840 19440
rect 18788 19397 18797 19431
rect 18797 19397 18831 19431
rect 18831 19397 18840 19431
rect 18788 19388 18840 19397
rect 20812 19388 20864 19440
rect 26056 19456 26108 19508
rect 27068 19456 27120 19508
rect 22928 19388 22980 19440
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 14004 19320 14056 19372
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 13452 19252 13504 19304
rect 12440 19184 12492 19236
rect 14004 19184 14056 19236
rect 14740 19363 14792 19372
rect 14740 19329 14749 19363
rect 14749 19329 14783 19363
rect 14783 19329 14792 19363
rect 14740 19320 14792 19329
rect 16120 19320 16172 19372
rect 15476 19252 15528 19304
rect 16580 19320 16632 19372
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 18512 19363 18564 19372
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 17960 19252 18012 19304
rect 23020 19320 23072 19372
rect 24216 19388 24268 19440
rect 23940 19363 23992 19372
rect 23940 19329 23949 19363
rect 23949 19329 23983 19363
rect 23983 19329 23992 19363
rect 23940 19320 23992 19329
rect 24032 19363 24084 19372
rect 24032 19329 24041 19363
rect 24041 19329 24075 19363
rect 24075 19329 24084 19363
rect 24032 19320 24084 19329
rect 26792 19388 26844 19440
rect 29000 19456 29052 19508
rect 19800 19295 19852 19304
rect 19800 19261 19809 19295
rect 19809 19261 19843 19295
rect 19843 19261 19852 19295
rect 19800 19252 19852 19261
rect 24860 19252 24912 19304
rect 25320 19363 25372 19372
rect 25320 19329 25329 19363
rect 25329 19329 25363 19363
rect 25363 19329 25372 19363
rect 25320 19320 25372 19329
rect 25780 19363 25832 19372
rect 25780 19329 25789 19363
rect 25789 19329 25823 19363
rect 25823 19329 25832 19363
rect 25780 19320 25832 19329
rect 25964 19363 26016 19372
rect 25964 19329 25973 19363
rect 25973 19329 26007 19363
rect 26007 19329 26016 19363
rect 25964 19320 26016 19329
rect 26700 19320 26752 19372
rect 25412 19252 25464 19304
rect 26332 19184 26384 19236
rect 6920 19116 6972 19168
rect 13360 19116 13412 19168
rect 15016 19116 15068 19168
rect 17040 19116 17092 19168
rect 19340 19116 19392 19168
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 23664 19116 23716 19168
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 27528 19363 27580 19372
rect 27528 19329 27537 19363
rect 27537 19329 27571 19363
rect 27571 19329 27580 19363
rect 27528 19320 27580 19329
rect 28172 19431 28224 19440
rect 28172 19397 28181 19431
rect 28181 19397 28215 19431
rect 28215 19397 28224 19431
rect 28172 19388 28224 19397
rect 31760 19456 31812 19508
rect 32128 19456 32180 19508
rect 29644 19388 29696 19440
rect 29920 19431 29972 19440
rect 29920 19397 29929 19431
rect 29929 19397 29963 19431
rect 29963 19397 29972 19431
rect 29920 19388 29972 19397
rect 30104 19431 30156 19440
rect 30104 19397 30113 19431
rect 30113 19397 30147 19431
rect 30147 19397 30156 19431
rect 30104 19388 30156 19397
rect 31576 19388 31628 19440
rect 32588 19456 32640 19508
rect 33324 19456 33376 19508
rect 33600 19456 33652 19508
rect 34152 19456 34204 19508
rect 35440 19456 35492 19508
rect 35716 19456 35768 19508
rect 36268 19456 36320 19508
rect 36636 19456 36688 19508
rect 32680 19431 32732 19440
rect 32680 19397 32689 19431
rect 32689 19397 32723 19431
rect 32723 19397 32732 19431
rect 32680 19388 32732 19397
rect 27896 19363 27948 19372
rect 27896 19329 27906 19363
rect 27906 19329 27940 19363
rect 27940 19329 27948 19363
rect 27896 19320 27948 19329
rect 27068 19252 27120 19304
rect 27620 19252 27672 19304
rect 29092 19363 29144 19372
rect 29092 19329 29101 19363
rect 29101 19329 29135 19363
rect 29135 19329 29144 19363
rect 29092 19320 29144 19329
rect 29460 19363 29512 19372
rect 29460 19329 29469 19363
rect 29469 19329 29503 19363
rect 29503 19329 29512 19363
rect 29460 19320 29512 19329
rect 29276 19252 29328 19304
rect 28080 19184 28132 19236
rect 29828 19320 29880 19372
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 33232 19363 33284 19372
rect 33232 19329 33241 19363
rect 33241 19329 33275 19363
rect 33275 19329 33284 19363
rect 33232 19320 33284 19329
rect 33508 19363 33560 19372
rect 33508 19329 33517 19363
rect 33517 19329 33551 19363
rect 33551 19329 33560 19363
rect 33508 19320 33560 19329
rect 33784 19363 33836 19372
rect 33784 19329 33793 19363
rect 33793 19329 33827 19363
rect 33827 19329 33836 19363
rect 33784 19320 33836 19329
rect 34796 19320 34848 19372
rect 36084 19388 36136 19440
rect 36912 19431 36964 19440
rect 36912 19397 36921 19431
rect 36921 19397 36955 19431
rect 36955 19397 36964 19431
rect 36912 19388 36964 19397
rect 34336 19252 34388 19304
rect 33140 19184 33192 19236
rect 35992 19363 36044 19372
rect 35992 19329 36001 19363
rect 36001 19329 36035 19363
rect 36035 19329 36044 19363
rect 35992 19320 36044 19329
rect 36268 19363 36320 19372
rect 36268 19329 36277 19363
rect 36277 19329 36311 19363
rect 36311 19329 36320 19363
rect 36268 19320 36320 19329
rect 36360 19320 36412 19372
rect 36820 19363 36872 19372
rect 36820 19329 36829 19363
rect 36829 19329 36863 19363
rect 36863 19329 36872 19363
rect 36820 19320 36872 19329
rect 37004 19320 37056 19372
rect 37372 19252 37424 19304
rect 38384 19252 38436 19304
rect 27804 19116 27856 19168
rect 28816 19116 28868 19168
rect 29184 19116 29236 19168
rect 31392 19116 31444 19168
rect 32772 19159 32824 19168
rect 32772 19125 32781 19159
rect 32781 19125 32815 19159
rect 32815 19125 32824 19159
rect 32772 19116 32824 19125
rect 33048 19159 33100 19168
rect 33048 19125 33057 19159
rect 33057 19125 33091 19159
rect 33091 19125 33100 19159
rect 33048 19116 33100 19125
rect 34152 19116 34204 19168
rect 34704 19116 34756 19168
rect 36636 19184 36688 19236
rect 36176 19116 36228 19168
rect 37004 19116 37056 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3516 18912 3568 18964
rect 3976 18912 4028 18964
rect 4528 18844 4580 18896
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 13176 18912 13228 18964
rect 14648 18955 14700 18964
rect 14648 18921 14657 18955
rect 14657 18921 14691 18955
rect 14691 18921 14700 18955
rect 14648 18912 14700 18921
rect 15844 18912 15896 18964
rect 17132 18912 17184 18964
rect 17408 18912 17460 18964
rect 23940 18912 23992 18964
rect 25780 18912 25832 18964
rect 27712 18912 27764 18964
rect 29092 18912 29144 18964
rect 10968 18844 11020 18896
rect 13360 18844 13412 18896
rect 6920 18819 6972 18828
rect 6920 18785 6929 18819
rect 6929 18785 6963 18819
rect 6963 18785 6972 18819
rect 6920 18776 6972 18785
rect 3240 18751 3292 18760
rect 3240 18717 3249 18751
rect 3249 18717 3283 18751
rect 3283 18717 3292 18751
rect 3240 18708 3292 18717
rect 3700 18708 3752 18760
rect 3976 18708 4028 18760
rect 4344 18751 4396 18760
rect 4344 18717 4353 18751
rect 4353 18717 4387 18751
rect 4387 18717 4396 18751
rect 4344 18708 4396 18717
rect 4528 18708 4580 18760
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 8024 18708 8076 18760
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 8668 18751 8720 18760
rect 8668 18717 8677 18751
rect 8677 18717 8711 18751
rect 8711 18717 8720 18751
rect 8668 18708 8720 18717
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 14004 18776 14056 18828
rect 6828 18640 6880 18692
rect 9404 18683 9456 18692
rect 9404 18649 9413 18683
rect 9413 18649 9447 18683
rect 9447 18649 9456 18683
rect 9404 18640 9456 18649
rect 10416 18640 10468 18692
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 13636 18751 13688 18760
rect 13636 18717 13645 18751
rect 13645 18717 13679 18751
rect 13679 18717 13688 18751
rect 13636 18708 13688 18717
rect 13912 18708 13964 18760
rect 14096 18751 14148 18760
rect 14096 18717 14105 18751
rect 14105 18717 14139 18751
rect 14139 18717 14148 18751
rect 14096 18708 14148 18717
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 15200 18751 15252 18760
rect 15200 18717 15209 18751
rect 15209 18717 15243 18751
rect 15243 18717 15252 18751
rect 15200 18708 15252 18717
rect 18696 18844 18748 18896
rect 27068 18844 27120 18896
rect 31760 18887 31812 18896
rect 31760 18853 31769 18887
rect 31769 18853 31803 18887
rect 31803 18853 31812 18887
rect 31760 18844 31812 18853
rect 32496 18844 32548 18896
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 16764 18819 16816 18828
rect 16764 18785 16773 18819
rect 16773 18785 16807 18819
rect 16807 18785 16816 18819
rect 16764 18776 16816 18785
rect 17592 18776 17644 18828
rect 16028 18708 16080 18760
rect 17408 18708 17460 18760
rect 18880 18776 18932 18828
rect 19340 18776 19392 18828
rect 22008 18776 22060 18828
rect 22468 18776 22520 18828
rect 23388 18776 23440 18828
rect 25964 18776 26016 18828
rect 18420 18708 18472 18760
rect 16304 18640 16356 18692
rect 17040 18683 17092 18692
rect 17040 18649 17065 18683
rect 17065 18649 17092 18683
rect 17040 18640 17092 18649
rect 17592 18683 17644 18692
rect 17592 18649 17601 18683
rect 17601 18649 17635 18683
rect 17635 18649 17644 18683
rect 17592 18640 17644 18649
rect 17776 18640 17828 18692
rect 4620 18572 4672 18624
rect 4804 18572 4856 18624
rect 8300 18572 8352 18624
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 13268 18572 13320 18624
rect 15292 18615 15344 18624
rect 15292 18581 15301 18615
rect 15301 18581 15335 18615
rect 15335 18581 15344 18615
rect 15292 18572 15344 18581
rect 15752 18615 15804 18624
rect 15752 18581 15761 18615
rect 15761 18581 15795 18615
rect 15795 18581 15804 18615
rect 15752 18572 15804 18581
rect 17868 18615 17920 18624
rect 17868 18581 17877 18615
rect 17877 18581 17911 18615
rect 17911 18581 17920 18615
rect 17868 18572 17920 18581
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 20812 18708 20864 18760
rect 21272 18708 21324 18760
rect 21732 18751 21784 18760
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 21456 18683 21508 18692
rect 21456 18649 21465 18683
rect 21465 18649 21499 18683
rect 21499 18649 21508 18683
rect 21916 18708 21968 18760
rect 21456 18640 21508 18649
rect 22744 18708 22796 18760
rect 23204 18708 23256 18760
rect 23940 18708 23992 18760
rect 24124 18751 24176 18760
rect 24124 18717 24133 18751
rect 24133 18717 24167 18751
rect 24167 18717 24176 18751
rect 24124 18708 24176 18717
rect 24860 18751 24912 18760
rect 24860 18717 24869 18751
rect 24869 18717 24903 18751
rect 24903 18717 24912 18751
rect 24860 18708 24912 18717
rect 25320 18751 25372 18760
rect 25320 18717 25329 18751
rect 25329 18717 25363 18751
rect 25363 18717 25372 18751
rect 25320 18708 25372 18717
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 26884 18751 26936 18760
rect 26884 18717 26893 18751
rect 26893 18717 26927 18751
rect 26927 18717 26936 18751
rect 26884 18708 26936 18717
rect 21732 18572 21784 18624
rect 27252 18776 27304 18828
rect 27804 18776 27856 18828
rect 27344 18751 27396 18760
rect 27344 18717 27353 18751
rect 27353 18717 27387 18751
rect 27387 18717 27396 18751
rect 27344 18708 27396 18717
rect 27896 18708 27948 18760
rect 28080 18708 28132 18760
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 26976 18683 27028 18692
rect 26976 18649 26985 18683
rect 26985 18649 27019 18683
rect 27019 18649 27028 18683
rect 26976 18640 27028 18649
rect 27712 18640 27764 18692
rect 31024 18776 31076 18828
rect 31484 18776 31536 18828
rect 33140 18819 33192 18828
rect 33140 18785 33149 18819
rect 33149 18785 33183 18819
rect 33183 18785 33192 18819
rect 33140 18776 33192 18785
rect 28448 18708 28500 18760
rect 28816 18751 28868 18760
rect 28816 18717 28825 18751
rect 28825 18717 28859 18751
rect 28859 18717 28868 18751
rect 28816 18708 28868 18717
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 29184 18751 29236 18760
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 29552 18751 29604 18760
rect 29552 18717 29561 18751
rect 29561 18717 29595 18751
rect 29595 18717 29604 18751
rect 29552 18708 29604 18717
rect 30196 18708 30248 18760
rect 32128 18751 32180 18760
rect 32128 18717 32137 18751
rect 32137 18717 32171 18751
rect 32171 18717 32180 18751
rect 32128 18708 32180 18717
rect 32220 18708 32272 18760
rect 32772 18751 32824 18760
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 33508 18912 33560 18964
rect 34428 18912 34480 18964
rect 35716 18912 35768 18964
rect 33416 18844 33468 18896
rect 36084 18912 36136 18964
rect 33508 18708 33560 18760
rect 29092 18683 29144 18692
rect 29092 18649 29101 18683
rect 29101 18649 29135 18683
rect 29135 18649 29144 18683
rect 29092 18640 29144 18649
rect 29276 18640 29328 18692
rect 30840 18640 30892 18692
rect 31484 18640 31536 18692
rect 23756 18615 23808 18624
rect 23756 18581 23765 18615
rect 23765 18581 23799 18615
rect 23799 18581 23808 18615
rect 23756 18572 23808 18581
rect 24124 18615 24176 18624
rect 24124 18581 24133 18615
rect 24133 18581 24167 18615
rect 24167 18581 24176 18615
rect 24124 18572 24176 18581
rect 28908 18572 28960 18624
rect 29368 18615 29420 18624
rect 29368 18581 29377 18615
rect 29377 18581 29411 18615
rect 29411 18581 29420 18615
rect 29368 18572 29420 18581
rect 29644 18615 29696 18624
rect 29644 18581 29653 18615
rect 29653 18581 29687 18615
rect 29687 18581 29696 18615
rect 29644 18572 29696 18581
rect 29920 18572 29972 18624
rect 32588 18640 32640 18692
rect 33692 18683 33744 18692
rect 33692 18649 33701 18683
rect 33701 18649 33735 18683
rect 33735 18649 33744 18683
rect 33692 18640 33744 18649
rect 34152 18819 34204 18828
rect 34152 18785 34161 18819
rect 34161 18785 34195 18819
rect 34195 18785 34204 18819
rect 34152 18776 34204 18785
rect 34980 18776 35032 18828
rect 36176 18887 36228 18896
rect 36176 18853 36185 18887
rect 36185 18853 36219 18887
rect 36219 18853 36228 18887
rect 36176 18844 36228 18853
rect 36360 18776 36412 18828
rect 37280 18887 37332 18896
rect 37280 18853 37289 18887
rect 37289 18853 37323 18887
rect 37323 18853 37332 18887
rect 37280 18844 37332 18853
rect 37740 18844 37792 18896
rect 34428 18640 34480 18692
rect 36636 18751 36688 18760
rect 36636 18717 36645 18751
rect 36645 18717 36679 18751
rect 36679 18717 36688 18751
rect 36636 18708 36688 18717
rect 37464 18708 37516 18760
rect 33600 18572 33652 18624
rect 34612 18572 34664 18624
rect 34704 18572 34756 18624
rect 35256 18572 35308 18624
rect 37096 18683 37148 18692
rect 37096 18649 37105 18683
rect 37105 18649 37139 18683
rect 37139 18649 37148 18683
rect 37096 18640 37148 18649
rect 37280 18572 37332 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 4528 18411 4580 18420
rect 4528 18377 4537 18411
rect 4537 18377 4571 18411
rect 4571 18377 4580 18411
rect 4528 18368 4580 18377
rect 2872 18232 2924 18284
rect 4712 18300 4764 18352
rect 3792 18232 3844 18284
rect 4436 18232 4488 18284
rect 4896 18275 4948 18284
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 4896 18232 4948 18241
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 7564 18300 7616 18352
rect 7932 18300 7984 18352
rect 8484 18368 8536 18420
rect 8668 18368 8720 18420
rect 9404 18368 9456 18420
rect 10324 18368 10376 18420
rect 13820 18368 13872 18420
rect 15200 18368 15252 18420
rect 16764 18368 16816 18420
rect 17592 18368 17644 18420
rect 1400 18164 1452 18216
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 3240 18207 3292 18216
rect 3240 18173 3249 18207
rect 3249 18173 3283 18207
rect 3283 18173 3292 18207
rect 3240 18164 3292 18173
rect 2964 18096 3016 18148
rect 3424 18096 3476 18148
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 4068 18096 4120 18148
rect 8300 18275 8352 18284
rect 8300 18241 8309 18275
rect 8309 18241 8343 18275
rect 8343 18241 8352 18275
rect 8300 18232 8352 18241
rect 8760 18232 8812 18284
rect 10876 18232 10928 18284
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 13360 18232 13412 18284
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 14924 18300 14976 18352
rect 15292 18300 15344 18352
rect 17132 18343 17184 18352
rect 17132 18309 17141 18343
rect 17141 18309 17175 18343
rect 17175 18309 17184 18343
rect 17132 18300 17184 18309
rect 17684 18300 17736 18352
rect 17868 18300 17920 18352
rect 7472 18164 7524 18216
rect 9128 18164 9180 18216
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 11888 18164 11940 18216
rect 12532 18164 12584 18216
rect 12992 18096 13044 18148
rect 13452 18139 13504 18148
rect 13452 18105 13461 18139
rect 13461 18105 13495 18139
rect 13495 18105 13504 18139
rect 13452 18096 13504 18105
rect 13728 18164 13780 18216
rect 14004 18207 14056 18216
rect 14004 18173 14013 18207
rect 14013 18173 14047 18207
rect 14047 18173 14056 18207
rect 14004 18164 14056 18173
rect 14188 18164 14240 18216
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 16120 18232 16172 18284
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 17776 18232 17828 18284
rect 17960 18275 18012 18284
rect 17960 18241 17969 18275
rect 17969 18241 18003 18275
rect 18003 18241 18012 18275
rect 17960 18232 18012 18241
rect 15016 18164 15068 18216
rect 17316 18164 17368 18216
rect 19524 18300 19576 18352
rect 22928 18368 22980 18420
rect 24860 18368 24912 18420
rect 25320 18368 25372 18420
rect 28264 18368 28316 18420
rect 28816 18368 28868 18420
rect 23480 18300 23532 18352
rect 20076 18232 20128 18284
rect 22468 18232 22520 18284
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 27252 18300 27304 18352
rect 24860 18232 24912 18284
rect 21272 18164 21324 18216
rect 23940 18207 23992 18216
rect 23940 18173 23949 18207
rect 23949 18173 23983 18207
rect 23983 18173 23992 18207
rect 23940 18164 23992 18173
rect 3976 18028 4028 18080
rect 4344 18028 4396 18080
rect 5080 18028 5132 18080
rect 6552 18028 6604 18080
rect 7564 18028 7616 18080
rect 11980 18028 12032 18080
rect 13544 18028 13596 18080
rect 14556 18071 14608 18080
rect 14556 18037 14565 18071
rect 14565 18037 14599 18071
rect 14599 18037 14608 18071
rect 14556 18028 14608 18037
rect 17684 18096 17736 18148
rect 16028 18028 16080 18080
rect 16948 18028 17000 18080
rect 23756 18096 23808 18148
rect 25504 18164 25556 18216
rect 26148 18232 26200 18284
rect 28172 18232 28224 18284
rect 28264 18232 28316 18284
rect 29184 18300 29236 18352
rect 27712 18164 27764 18216
rect 28448 18164 28500 18216
rect 29000 18275 29052 18284
rect 29000 18241 29009 18275
rect 29009 18241 29043 18275
rect 29043 18241 29052 18275
rect 29000 18232 29052 18241
rect 29368 18232 29420 18284
rect 30656 18300 30708 18352
rect 31392 18343 31444 18352
rect 31392 18309 31401 18343
rect 31401 18309 31435 18343
rect 31435 18309 31444 18343
rect 31392 18300 31444 18309
rect 32128 18300 32180 18352
rect 29092 18207 29144 18216
rect 29092 18173 29101 18207
rect 29101 18173 29135 18207
rect 29135 18173 29144 18207
rect 29092 18164 29144 18173
rect 30932 18164 30984 18216
rect 32036 18232 32088 18284
rect 33048 18232 33100 18284
rect 33416 18275 33468 18284
rect 33416 18241 33425 18275
rect 33425 18241 33459 18275
rect 33459 18241 33468 18275
rect 33416 18232 33468 18241
rect 33232 18207 33284 18216
rect 19616 18028 19668 18080
rect 21916 18028 21968 18080
rect 25412 18028 25464 18080
rect 28724 18028 28776 18080
rect 31668 18096 31720 18148
rect 33232 18173 33241 18207
rect 33241 18173 33275 18207
rect 33275 18173 33284 18207
rect 33232 18164 33284 18173
rect 33600 18207 33652 18216
rect 33600 18173 33609 18207
rect 33609 18173 33643 18207
rect 33643 18173 33652 18207
rect 33600 18164 33652 18173
rect 34428 18368 34480 18420
rect 37372 18368 37424 18420
rect 34520 18300 34572 18352
rect 34612 18275 34664 18284
rect 34612 18241 34621 18275
rect 34621 18241 34655 18275
rect 34655 18241 34664 18275
rect 34612 18232 34664 18241
rect 34704 18232 34756 18284
rect 34980 18275 35032 18284
rect 34980 18241 34989 18275
rect 34989 18241 35023 18275
rect 35023 18241 35032 18275
rect 34980 18232 35032 18241
rect 35256 18275 35308 18284
rect 35256 18241 35265 18275
rect 35265 18241 35299 18275
rect 35299 18241 35308 18275
rect 35256 18232 35308 18241
rect 34428 18164 34480 18216
rect 33508 18028 33560 18080
rect 34244 18028 34296 18080
rect 35808 18028 35860 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1768 17824 1820 17876
rect 4712 17824 4764 17876
rect 4988 17824 5040 17876
rect 5356 17824 5408 17876
rect 8760 17867 8812 17876
rect 8760 17833 8769 17867
rect 8769 17833 8803 17867
rect 8803 17833 8812 17867
rect 8760 17824 8812 17833
rect 11888 17824 11940 17876
rect 5080 17799 5132 17808
rect 5080 17765 5089 17799
rect 5089 17765 5123 17799
rect 5123 17765 5132 17799
rect 5080 17756 5132 17765
rect 12624 17824 12676 17876
rect 12900 17824 12952 17876
rect 13820 17824 13872 17876
rect 14924 17824 14976 17876
rect 15752 17824 15804 17876
rect 18420 17867 18472 17876
rect 18420 17833 18429 17867
rect 18429 17833 18463 17867
rect 18463 17833 18472 17867
rect 18420 17824 18472 17833
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 24860 17824 24912 17876
rect 27252 17867 27304 17876
rect 27252 17833 27261 17867
rect 27261 17833 27295 17867
rect 27295 17833 27304 17867
rect 27252 17824 27304 17833
rect 27988 17824 28040 17876
rect 30196 17824 30248 17876
rect 30840 17824 30892 17876
rect 30932 17867 30984 17876
rect 30932 17833 30941 17867
rect 30941 17833 30975 17867
rect 30975 17833 30984 17867
rect 30932 17824 30984 17833
rect 6552 17731 6604 17740
rect 6552 17697 6561 17731
rect 6561 17697 6595 17731
rect 6595 17697 6604 17731
rect 6552 17688 6604 17697
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 7932 17731 7984 17740
rect 7932 17697 7941 17731
rect 7941 17697 7975 17731
rect 7975 17697 7984 17731
rect 7932 17688 7984 17697
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 4160 17620 4212 17672
rect 4436 17663 4488 17672
rect 4436 17629 4445 17663
rect 4445 17629 4479 17663
rect 4479 17629 4488 17663
rect 4436 17620 4488 17629
rect 7564 17620 7616 17672
rect 12532 17688 12584 17740
rect 4528 17552 4580 17604
rect 5080 17552 5132 17604
rect 5908 17552 5960 17604
rect 10416 17620 10468 17672
rect 9220 17552 9272 17604
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 9312 17552 9364 17561
rect 4896 17484 4948 17536
rect 5264 17484 5316 17536
rect 7012 17484 7064 17536
rect 7656 17484 7708 17536
rect 8116 17484 8168 17536
rect 11152 17595 11204 17604
rect 11152 17561 11161 17595
rect 11161 17561 11195 17595
rect 11195 17561 11204 17595
rect 11152 17552 11204 17561
rect 11796 17552 11848 17604
rect 10876 17484 10928 17536
rect 12900 17620 12952 17672
rect 26792 17756 26844 17808
rect 28264 17756 28316 17808
rect 30288 17756 30340 17808
rect 33232 17867 33284 17876
rect 33232 17833 33241 17867
rect 33241 17833 33275 17867
rect 33275 17833 33284 17867
rect 33232 17824 33284 17833
rect 33324 17824 33376 17876
rect 33600 17824 33652 17876
rect 37096 17824 37148 17876
rect 13820 17688 13872 17740
rect 14740 17688 14792 17740
rect 17960 17688 18012 17740
rect 19432 17688 19484 17740
rect 23572 17688 23624 17740
rect 25596 17688 25648 17740
rect 34520 17756 34572 17808
rect 32128 17731 32180 17740
rect 13544 17620 13596 17672
rect 15476 17620 15528 17672
rect 18696 17620 18748 17672
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 23940 17663 23992 17672
rect 23940 17629 23949 17663
rect 23949 17629 23983 17663
rect 23983 17629 23992 17663
rect 23940 17620 23992 17629
rect 24124 17620 24176 17672
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 13084 17552 13136 17604
rect 14004 17552 14056 17604
rect 13728 17484 13780 17536
rect 16948 17595 17000 17604
rect 16948 17561 16957 17595
rect 16957 17561 16991 17595
rect 16991 17561 17000 17595
rect 16948 17552 17000 17561
rect 16120 17484 16172 17536
rect 19340 17552 19392 17604
rect 21272 17552 21324 17604
rect 21548 17595 21600 17604
rect 21548 17561 21557 17595
rect 21557 17561 21591 17595
rect 21591 17561 21600 17595
rect 21548 17552 21600 17561
rect 22100 17552 22152 17604
rect 22836 17552 22888 17604
rect 23848 17552 23900 17604
rect 24492 17552 24544 17604
rect 17960 17484 18012 17536
rect 23756 17484 23808 17536
rect 24124 17484 24176 17536
rect 24860 17484 24912 17536
rect 25228 17620 25280 17672
rect 25504 17620 25556 17672
rect 26148 17663 26200 17672
rect 26148 17629 26157 17663
rect 26157 17629 26191 17663
rect 26191 17629 26200 17663
rect 26148 17620 26200 17629
rect 26608 17663 26660 17672
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 26792 17663 26844 17672
rect 26792 17629 26801 17663
rect 26801 17629 26835 17663
rect 26835 17629 26844 17663
rect 26792 17620 26844 17629
rect 27804 17620 27856 17672
rect 27988 17620 28040 17672
rect 28172 17663 28224 17672
rect 28172 17629 28181 17663
rect 28181 17629 28215 17663
rect 28215 17629 28224 17663
rect 28172 17620 28224 17629
rect 28264 17663 28316 17672
rect 28264 17629 28273 17663
rect 28273 17629 28307 17663
rect 28307 17629 28316 17663
rect 28264 17620 28316 17629
rect 28356 17552 28408 17604
rect 28724 17663 28776 17672
rect 28724 17629 28733 17663
rect 28733 17629 28767 17663
rect 28767 17629 28776 17663
rect 28724 17620 28776 17629
rect 28908 17663 28960 17672
rect 28908 17629 28917 17663
rect 28917 17629 28951 17663
rect 28951 17629 28960 17663
rect 28908 17620 28960 17629
rect 29000 17663 29052 17672
rect 29000 17629 29009 17663
rect 29009 17629 29043 17663
rect 29043 17629 29052 17663
rect 29000 17620 29052 17629
rect 29092 17663 29144 17672
rect 29092 17629 29101 17663
rect 29101 17629 29135 17663
rect 29135 17629 29144 17663
rect 29092 17620 29144 17629
rect 29644 17620 29696 17672
rect 30012 17663 30064 17672
rect 30012 17629 30021 17663
rect 30021 17629 30055 17663
rect 30055 17629 30064 17663
rect 30012 17620 30064 17629
rect 30196 17663 30248 17672
rect 30196 17629 30205 17663
rect 30205 17629 30239 17663
rect 30239 17629 30248 17663
rect 30196 17620 30248 17629
rect 29184 17552 29236 17604
rect 30380 17663 30432 17672
rect 30380 17629 30389 17663
rect 30389 17629 30423 17663
rect 30423 17629 30432 17663
rect 32128 17697 32137 17731
rect 32137 17697 32171 17731
rect 32171 17697 32180 17731
rect 32128 17688 32180 17697
rect 32220 17731 32272 17740
rect 32220 17697 32229 17731
rect 32229 17697 32263 17731
rect 32263 17697 32272 17731
rect 32220 17688 32272 17697
rect 32312 17688 32364 17740
rect 34796 17688 34848 17740
rect 35808 17731 35860 17740
rect 35808 17697 35817 17731
rect 35817 17697 35851 17731
rect 35851 17697 35860 17731
rect 35808 17688 35860 17697
rect 30380 17620 30432 17629
rect 30656 17620 30708 17672
rect 30932 17620 30984 17672
rect 31668 17620 31720 17672
rect 32036 17663 32088 17672
rect 32036 17629 32045 17663
rect 32045 17629 32079 17663
rect 32079 17629 32088 17663
rect 32036 17620 32088 17629
rect 31024 17552 31076 17604
rect 32404 17663 32456 17672
rect 32404 17629 32413 17663
rect 32413 17629 32447 17663
rect 32447 17629 32456 17663
rect 32404 17620 32456 17629
rect 32496 17620 32548 17672
rect 33324 17663 33376 17672
rect 33324 17629 33333 17663
rect 33333 17629 33367 17663
rect 33367 17629 33376 17663
rect 33324 17620 33376 17629
rect 26884 17484 26936 17536
rect 28264 17484 28316 17536
rect 29460 17484 29512 17536
rect 30196 17484 30248 17536
rect 30564 17484 30616 17536
rect 32680 17527 32732 17536
rect 32680 17493 32689 17527
rect 32689 17493 32723 17527
rect 32723 17493 32732 17527
rect 32680 17484 32732 17493
rect 34428 17620 34480 17672
rect 34612 17620 34664 17672
rect 34704 17552 34756 17604
rect 36176 17552 36228 17604
rect 34796 17484 34848 17536
rect 37648 17484 37700 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 5264 17280 5316 17332
rect 5448 17280 5500 17332
rect 7840 17280 7892 17332
rect 9312 17280 9364 17332
rect 10876 17323 10928 17332
rect 10876 17289 10885 17323
rect 10885 17289 10919 17323
rect 10919 17289 10928 17323
rect 10876 17280 10928 17289
rect 11152 17280 11204 17332
rect 11980 17323 12032 17332
rect 11980 17289 11989 17323
rect 11989 17289 12023 17323
rect 12023 17289 12032 17323
rect 11980 17280 12032 17289
rect 13636 17280 13688 17332
rect 13820 17323 13872 17332
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 14556 17280 14608 17332
rect 21548 17280 21600 17332
rect 22836 17280 22888 17332
rect 24860 17280 24912 17332
rect 24952 17280 25004 17332
rect 26608 17280 26660 17332
rect 28172 17280 28224 17332
rect 28356 17280 28408 17332
rect 29920 17280 29972 17332
rect 3240 17212 3292 17264
rect 3884 17212 3936 17264
rect 4436 17255 4488 17264
rect 4436 17221 4445 17255
rect 4445 17221 4479 17255
rect 4479 17221 4488 17255
rect 4436 17212 4488 17221
rect 8116 17212 8168 17264
rect 9128 17255 9180 17264
rect 9128 17221 9137 17255
rect 9137 17221 9171 17255
rect 9171 17221 9180 17255
rect 9128 17212 9180 17221
rect 9220 17212 9272 17264
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 5724 17144 5776 17196
rect 3148 17076 3200 17128
rect 3792 17076 3844 17128
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 2964 17008 3016 17060
rect 5908 17076 5960 17128
rect 2412 16983 2464 16992
rect 2412 16949 2421 16983
rect 2421 16949 2455 16983
rect 2455 16949 2464 16983
rect 2412 16940 2464 16949
rect 2780 16983 2832 16992
rect 2780 16949 2789 16983
rect 2789 16949 2823 16983
rect 2823 16949 2832 16983
rect 2780 16940 2832 16949
rect 2872 16983 2924 16992
rect 2872 16949 2881 16983
rect 2881 16949 2915 16983
rect 2915 16949 2924 16983
rect 2872 16940 2924 16949
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 4712 16940 4764 16992
rect 5540 16940 5592 16992
rect 6736 16983 6788 16992
rect 6736 16949 6745 16983
rect 6745 16949 6779 16983
rect 6779 16949 6788 16983
rect 6736 16940 6788 16949
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 13084 17144 13136 17196
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 7656 17076 7708 17128
rect 9680 17076 9732 17128
rect 10692 17076 10744 17128
rect 15936 17212 15988 17264
rect 18788 17255 18840 17264
rect 18788 17221 18797 17255
rect 18797 17221 18831 17255
rect 18831 17221 18840 17255
rect 18788 17212 18840 17221
rect 18972 17255 19024 17264
rect 18972 17221 18997 17255
rect 18997 17221 19024 17255
rect 18972 17212 19024 17221
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 15200 17187 15252 17196
rect 15200 17153 15209 17187
rect 15209 17153 15243 17187
rect 15243 17153 15252 17187
rect 15200 17144 15252 17153
rect 18420 17187 18472 17196
rect 18420 17153 18429 17187
rect 18429 17153 18463 17187
rect 18463 17153 18472 17187
rect 18420 17144 18472 17153
rect 19892 17187 19944 17196
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 23480 17144 23532 17196
rect 19524 17076 19576 17128
rect 20168 17119 20220 17128
rect 20168 17085 20177 17119
rect 20177 17085 20211 17119
rect 20211 17085 20220 17119
rect 20168 17076 20220 17085
rect 21088 17076 21140 17128
rect 23204 17076 23256 17128
rect 23572 17076 23624 17128
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 24124 17144 24176 17196
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 24768 17187 24820 17196
rect 24768 17153 24777 17187
rect 24777 17153 24811 17187
rect 24811 17153 24820 17187
rect 24768 17144 24820 17153
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 25596 17187 25648 17196
rect 25596 17153 25605 17187
rect 25605 17153 25639 17187
rect 25639 17153 25648 17187
rect 25596 17144 25648 17153
rect 11336 17008 11388 17060
rect 19984 17008 20036 17060
rect 26792 17144 26844 17196
rect 26884 17144 26936 17196
rect 26056 17076 26108 17128
rect 29092 17187 29144 17196
rect 29092 17153 29101 17187
rect 29101 17153 29135 17187
rect 29135 17153 29144 17187
rect 29092 17144 29144 17153
rect 29184 17119 29236 17128
rect 29184 17085 29193 17119
rect 29193 17085 29227 17119
rect 29227 17085 29236 17119
rect 29184 17076 29236 17085
rect 29460 17187 29512 17196
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 31024 17212 31076 17264
rect 29920 17187 29972 17196
rect 29920 17153 29930 17187
rect 29930 17153 29964 17187
rect 29964 17153 29972 17187
rect 29920 17144 29972 17153
rect 30196 17187 30248 17196
rect 30196 17153 30205 17187
rect 30205 17153 30239 17187
rect 30239 17153 30248 17187
rect 30196 17144 30248 17153
rect 30288 17187 30340 17196
rect 30288 17153 30302 17187
rect 30302 17153 30336 17187
rect 30336 17153 30340 17187
rect 30288 17144 30340 17153
rect 30656 17187 30708 17196
rect 30656 17153 30665 17187
rect 30665 17153 30699 17187
rect 30699 17153 30708 17187
rect 30656 17144 30708 17153
rect 26148 17008 26200 17060
rect 32404 17280 32456 17332
rect 32496 17212 32548 17264
rect 36636 17280 36688 17332
rect 32220 17144 32272 17196
rect 9772 16940 9824 16992
rect 15936 16940 15988 16992
rect 18236 16940 18288 16992
rect 18696 16940 18748 16992
rect 19156 16983 19208 16992
rect 19156 16949 19165 16983
rect 19165 16949 19199 16983
rect 19199 16949 19208 16983
rect 19156 16940 19208 16949
rect 19524 16940 19576 16992
rect 20260 16940 20312 16992
rect 24860 16940 24912 16992
rect 25872 16940 25924 16992
rect 30012 16940 30064 16992
rect 30104 16940 30156 16992
rect 31300 16940 31352 16992
rect 31392 16983 31444 16992
rect 31392 16949 31401 16983
rect 31401 16949 31435 16983
rect 31435 16949 31444 16983
rect 31392 16940 31444 16949
rect 31760 16983 31812 16992
rect 31760 16949 31769 16983
rect 31769 16949 31803 16983
rect 31803 16949 31812 16983
rect 31760 16940 31812 16949
rect 32588 17187 32640 17196
rect 32588 17153 32597 17187
rect 32597 17153 32631 17187
rect 32631 17153 32640 17187
rect 32588 17144 32640 17153
rect 33140 17187 33192 17196
rect 33140 17153 33149 17187
rect 33149 17153 33183 17187
rect 33183 17153 33192 17187
rect 33140 17144 33192 17153
rect 34428 17212 34480 17264
rect 32956 17076 33008 17128
rect 33692 17144 33744 17196
rect 34244 17187 34296 17196
rect 34244 17153 34253 17187
rect 34253 17153 34287 17187
rect 34287 17153 34296 17187
rect 34244 17144 34296 17153
rect 35992 17144 36044 17196
rect 34612 17119 34664 17128
rect 34612 17085 34621 17119
rect 34621 17085 34655 17119
rect 34655 17085 34664 17119
rect 34612 17076 34664 17085
rect 33416 17051 33468 17060
rect 33416 17017 33425 17051
rect 33425 17017 33459 17051
rect 33459 17017 33468 17051
rect 33416 17008 33468 17017
rect 34520 17008 34572 17060
rect 33692 16940 33744 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3148 16736 3200 16788
rect 7012 16779 7064 16788
rect 7012 16745 7021 16779
rect 7021 16745 7055 16779
rect 7055 16745 7064 16779
rect 7012 16736 7064 16745
rect 12716 16736 12768 16788
rect 15016 16736 15068 16788
rect 17224 16736 17276 16788
rect 18604 16736 18656 16788
rect 18788 16736 18840 16788
rect 25228 16736 25280 16788
rect 29184 16736 29236 16788
rect 30288 16736 30340 16788
rect 5356 16668 5408 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 4068 16600 4120 16652
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 9772 16600 9824 16652
rect 1676 16507 1728 16516
rect 1676 16473 1685 16507
rect 1685 16473 1719 16507
rect 1719 16473 1728 16507
rect 1676 16464 1728 16473
rect 2688 16464 2740 16516
rect 2504 16396 2556 16448
rect 3240 16507 3292 16516
rect 3240 16473 3249 16507
rect 3249 16473 3283 16507
rect 3283 16473 3292 16507
rect 3240 16464 3292 16473
rect 9220 16532 9272 16584
rect 11336 16575 11388 16584
rect 11336 16541 11345 16575
rect 11345 16541 11379 16575
rect 11379 16541 11388 16575
rect 11336 16532 11388 16541
rect 13728 16600 13780 16652
rect 15752 16668 15804 16720
rect 24860 16711 24912 16720
rect 24860 16677 24869 16711
rect 24869 16677 24903 16711
rect 24903 16677 24912 16711
rect 24860 16668 24912 16677
rect 25688 16668 25740 16720
rect 26056 16668 26108 16720
rect 28632 16668 28684 16720
rect 30932 16711 30984 16720
rect 30932 16677 30941 16711
rect 30941 16677 30975 16711
rect 30975 16677 30984 16711
rect 30932 16668 30984 16677
rect 13268 16575 13320 16584
rect 13268 16541 13277 16575
rect 13277 16541 13311 16575
rect 13311 16541 13320 16575
rect 13268 16532 13320 16541
rect 13820 16532 13872 16584
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 15568 16575 15620 16584
rect 15568 16541 15577 16575
rect 15577 16541 15611 16575
rect 15611 16541 15620 16575
rect 15568 16532 15620 16541
rect 5264 16464 5316 16516
rect 5908 16464 5960 16516
rect 6368 16464 6420 16516
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 3148 16396 3200 16405
rect 4160 16396 4212 16448
rect 8024 16464 8076 16516
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 19524 16643 19576 16652
rect 19524 16609 19533 16643
rect 19533 16609 19567 16643
rect 19567 16609 19576 16643
rect 19524 16600 19576 16609
rect 20260 16600 20312 16652
rect 16304 16575 16356 16584
rect 16304 16541 16313 16575
rect 16313 16541 16347 16575
rect 16347 16541 16356 16575
rect 16304 16532 16356 16541
rect 19064 16532 19116 16584
rect 23020 16600 23072 16652
rect 24032 16600 24084 16652
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 9404 16396 9456 16448
rect 9864 16396 9916 16448
rect 17960 16464 18012 16516
rect 22008 16532 22060 16584
rect 22100 16532 22152 16584
rect 25136 16575 25188 16584
rect 25136 16541 25145 16575
rect 25145 16541 25179 16575
rect 25179 16541 25188 16575
rect 25136 16532 25188 16541
rect 25412 16600 25464 16652
rect 26792 16643 26844 16652
rect 26792 16609 26801 16643
rect 26801 16609 26835 16643
rect 26835 16609 26844 16643
rect 26792 16600 26844 16609
rect 28080 16600 28132 16652
rect 30104 16643 30156 16652
rect 30104 16609 30113 16643
rect 30113 16609 30147 16643
rect 30147 16609 30156 16643
rect 30104 16600 30156 16609
rect 33140 16736 33192 16788
rect 34796 16736 34848 16788
rect 31300 16668 31352 16720
rect 32496 16711 32548 16720
rect 32496 16677 32505 16711
rect 32505 16677 32539 16711
rect 32539 16677 32548 16711
rect 32496 16668 32548 16677
rect 31760 16600 31812 16652
rect 19432 16464 19484 16516
rect 19984 16464 20036 16516
rect 22560 16507 22612 16516
rect 22560 16473 22569 16507
rect 22569 16473 22603 16507
rect 22603 16473 22612 16507
rect 22560 16464 22612 16473
rect 23020 16464 23072 16516
rect 23940 16464 23992 16516
rect 11428 16396 11480 16448
rect 15936 16396 15988 16448
rect 21088 16396 21140 16448
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 24032 16439 24084 16448
rect 24032 16405 24041 16439
rect 24041 16405 24075 16439
rect 24075 16405 24084 16439
rect 24032 16396 24084 16405
rect 27988 16464 28040 16516
rect 29000 16464 29052 16516
rect 29368 16464 29420 16516
rect 31392 16575 31444 16584
rect 31392 16541 31401 16575
rect 31401 16541 31435 16575
rect 31435 16541 31444 16575
rect 31392 16532 31444 16541
rect 32404 16600 32456 16652
rect 32680 16600 32732 16652
rect 32772 16575 32824 16584
rect 32772 16541 32781 16575
rect 32781 16541 32815 16575
rect 32815 16541 32824 16575
rect 32772 16532 32824 16541
rect 29460 16396 29512 16448
rect 30472 16396 30524 16448
rect 30564 16439 30616 16448
rect 30564 16405 30573 16439
rect 30573 16405 30607 16439
rect 30607 16405 30616 16439
rect 30564 16396 30616 16405
rect 30656 16396 30708 16448
rect 33324 16464 33376 16516
rect 31668 16396 31720 16448
rect 36176 16464 36228 16516
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 2872 16192 2924 16244
rect 1676 16124 1728 16176
rect 2504 16124 2556 16176
rect 2412 16099 2464 16108
rect 2412 16065 2421 16099
rect 2421 16065 2455 16099
rect 2455 16065 2464 16099
rect 2412 16056 2464 16065
rect 2780 16056 2832 16108
rect 4160 16192 4212 16244
rect 5448 16192 5500 16244
rect 7564 16192 7616 16244
rect 9404 16192 9456 16244
rect 11336 16192 11388 16244
rect 4068 16124 4120 16176
rect 5080 16056 5132 16108
rect 2964 15988 3016 16040
rect 3240 15852 3292 15904
rect 4896 15852 4948 15904
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 6828 16124 6880 16176
rect 9128 16124 9180 16176
rect 10048 16124 10100 16176
rect 7932 16056 7984 16108
rect 6368 15988 6420 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 15292 16192 15344 16244
rect 15568 16235 15620 16244
rect 15568 16201 15577 16235
rect 15577 16201 15611 16235
rect 15611 16201 15620 16235
rect 15568 16192 15620 16201
rect 17316 16235 17368 16244
rect 17316 16201 17325 16235
rect 17325 16201 17359 16235
rect 17359 16201 17368 16235
rect 17316 16192 17368 16201
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 19892 16192 19944 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 21180 16192 21232 16244
rect 22560 16192 22612 16244
rect 24032 16192 24084 16244
rect 25136 16192 25188 16244
rect 13084 16124 13136 16176
rect 13636 15988 13688 16040
rect 13820 16056 13872 16108
rect 15844 16124 15896 16176
rect 14740 16099 14792 16108
rect 14740 16065 14749 16099
rect 14749 16065 14783 16099
rect 14783 16065 14792 16099
rect 14740 16056 14792 16065
rect 15200 16056 15252 16108
rect 16028 16099 16080 16108
rect 16028 16065 16037 16099
rect 16037 16065 16071 16099
rect 16071 16065 16080 16099
rect 16028 16056 16080 16065
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15108 15920 15160 15972
rect 15384 15988 15436 16040
rect 15660 15920 15712 15972
rect 16672 16099 16724 16108
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 16764 16056 16816 16108
rect 16396 15988 16448 16040
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18788 16056 18840 16108
rect 20260 16099 20312 16108
rect 20260 16065 20269 16099
rect 20269 16065 20303 16099
rect 20303 16065 20312 16099
rect 20260 16056 20312 16065
rect 19616 15988 19668 16040
rect 20168 15988 20220 16040
rect 21088 16124 21140 16176
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 24124 16124 24176 16176
rect 20536 15988 20588 16040
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 28080 16235 28132 16244
rect 28080 16201 28089 16235
rect 28089 16201 28123 16235
rect 28123 16201 28132 16235
rect 28080 16192 28132 16201
rect 28264 16235 28316 16244
rect 28264 16201 28273 16235
rect 28273 16201 28307 16235
rect 28307 16201 28316 16235
rect 28264 16192 28316 16201
rect 19340 15920 19392 15972
rect 13544 15852 13596 15904
rect 13820 15852 13872 15904
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 15200 15852 15252 15904
rect 16212 15852 16264 15904
rect 23204 15920 23256 15972
rect 25228 16031 25280 16040
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 31392 16192 31444 16244
rect 32220 16192 32272 16244
rect 31208 16124 31260 16176
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 31668 16124 31720 16176
rect 29460 16056 29512 16065
rect 27988 15988 28040 16040
rect 29000 15988 29052 16040
rect 29092 16031 29144 16040
rect 29092 15997 29101 16031
rect 29101 15997 29135 16031
rect 29135 15997 29144 16031
rect 29092 15988 29144 15997
rect 29552 15988 29604 16040
rect 30472 16031 30524 16040
rect 30472 15997 30481 16031
rect 30481 15997 30515 16031
rect 30515 15997 30524 16031
rect 30472 15988 30524 15997
rect 35348 16056 35400 16108
rect 32864 15988 32916 16040
rect 34612 15988 34664 16040
rect 34796 15988 34848 16040
rect 27804 15920 27856 15972
rect 28632 15963 28684 15972
rect 28632 15929 28641 15963
rect 28641 15929 28675 15963
rect 28675 15929 28684 15963
rect 28632 15920 28684 15929
rect 33140 15920 33192 15972
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 26884 15852 26936 15904
rect 30656 15852 30708 15904
rect 32956 15852 33008 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2504 15648 2556 15700
rect 4620 15648 4672 15700
rect 5264 15648 5316 15700
rect 7012 15648 7064 15700
rect 10876 15648 10928 15700
rect 4252 15580 4304 15632
rect 5080 15580 5132 15632
rect 13268 15691 13320 15700
rect 13268 15657 13277 15691
rect 13277 15657 13311 15691
rect 13311 15657 13320 15691
rect 13268 15648 13320 15657
rect 15384 15648 15436 15700
rect 16028 15648 16080 15700
rect 16948 15648 17000 15700
rect 18420 15648 18472 15700
rect 23112 15648 23164 15700
rect 13636 15623 13688 15632
rect 4068 15512 4120 15564
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 2964 15444 3016 15496
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 5356 15512 5408 15564
rect 5264 15444 5316 15496
rect 9220 15444 9272 15496
rect 13636 15589 13645 15623
rect 13645 15589 13679 15623
rect 13679 15589 13688 15623
rect 13636 15580 13688 15589
rect 16396 15623 16448 15632
rect 16396 15589 16405 15623
rect 16405 15589 16439 15623
rect 16439 15589 16448 15623
rect 16396 15580 16448 15589
rect 16672 15623 16724 15632
rect 16672 15589 16681 15623
rect 16681 15589 16715 15623
rect 16715 15589 16724 15623
rect 16672 15580 16724 15589
rect 16856 15580 16908 15632
rect 25228 15623 25280 15632
rect 25228 15589 25237 15623
rect 25237 15589 25271 15623
rect 25271 15589 25280 15623
rect 25228 15580 25280 15589
rect 12716 15512 12768 15564
rect 14372 15555 14424 15564
rect 14372 15521 14381 15555
rect 14381 15521 14415 15555
rect 14415 15521 14424 15555
rect 14372 15512 14424 15521
rect 14832 15512 14884 15564
rect 16028 15555 16080 15564
rect 16028 15521 16037 15555
rect 16037 15521 16071 15555
rect 16071 15521 16080 15555
rect 16028 15512 16080 15521
rect 3148 15376 3200 15428
rect 2412 15308 2464 15360
rect 4896 15308 4948 15360
rect 12900 15444 12952 15496
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 15476 15444 15528 15496
rect 15752 15444 15804 15496
rect 16212 15487 16264 15496
rect 16212 15453 16221 15487
rect 16221 15453 16255 15487
rect 16255 15453 16264 15487
rect 16212 15444 16264 15453
rect 18052 15512 18104 15564
rect 20720 15512 20772 15564
rect 24124 15512 24176 15564
rect 25688 15555 25740 15564
rect 25688 15521 25697 15555
rect 25697 15521 25731 15555
rect 25731 15521 25740 15555
rect 25688 15512 25740 15521
rect 27804 15623 27856 15632
rect 27804 15589 27813 15623
rect 27813 15589 27847 15623
rect 27847 15589 27856 15623
rect 27804 15580 27856 15589
rect 11060 15419 11112 15428
rect 11060 15385 11069 15419
rect 11069 15385 11103 15419
rect 11103 15385 11112 15419
rect 11060 15376 11112 15385
rect 11796 15376 11848 15428
rect 12716 15376 12768 15428
rect 12992 15376 13044 15428
rect 16764 15376 16816 15428
rect 17132 15376 17184 15428
rect 18880 15444 18932 15496
rect 19064 15444 19116 15496
rect 18696 15376 18748 15428
rect 15660 15308 15712 15360
rect 19248 15419 19300 15428
rect 19248 15385 19257 15419
rect 19257 15385 19291 15419
rect 19291 15385 19300 15419
rect 19248 15376 19300 15385
rect 22008 15376 22060 15428
rect 22100 15376 22152 15428
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 26884 15444 26936 15496
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 32864 15512 32916 15564
rect 37280 15487 37332 15496
rect 37280 15453 37289 15487
rect 37289 15453 37323 15487
rect 37323 15453 37332 15487
rect 37280 15444 37332 15453
rect 28172 15419 28224 15428
rect 28172 15385 28181 15419
rect 28181 15385 28215 15419
rect 28215 15385 28224 15419
rect 28172 15376 28224 15385
rect 32956 15376 33008 15428
rect 34428 15376 34480 15428
rect 34520 15376 34572 15428
rect 35440 15419 35492 15428
rect 35440 15385 35449 15419
rect 35449 15385 35483 15419
rect 35483 15385 35492 15419
rect 35440 15376 35492 15385
rect 18880 15308 18932 15360
rect 19432 15308 19484 15360
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 23664 15351 23716 15360
rect 23664 15317 23673 15351
rect 23673 15317 23707 15351
rect 23707 15317 23716 15351
rect 23664 15308 23716 15317
rect 23940 15308 23992 15360
rect 24124 15351 24176 15360
rect 24124 15317 24133 15351
rect 24133 15317 24167 15351
rect 24167 15317 24176 15351
rect 24124 15308 24176 15317
rect 24400 15351 24452 15360
rect 24400 15317 24409 15351
rect 24409 15317 24443 15351
rect 24443 15317 24452 15351
rect 24400 15308 24452 15317
rect 27620 15351 27672 15360
rect 27620 15317 27629 15351
rect 27629 15317 27663 15351
rect 27663 15317 27672 15351
rect 27620 15308 27672 15317
rect 27712 15351 27764 15360
rect 27712 15317 27721 15351
rect 27721 15317 27755 15351
rect 27755 15317 27764 15351
rect 27712 15308 27764 15317
rect 30104 15308 30156 15360
rect 34704 15308 34756 15360
rect 36636 15351 36688 15360
rect 36636 15317 36645 15351
rect 36645 15317 36679 15351
rect 36679 15317 36688 15351
rect 36636 15308 36688 15317
rect 38476 15351 38528 15360
rect 38476 15317 38485 15351
rect 38485 15317 38519 15351
rect 38519 15317 38528 15351
rect 38476 15308 38528 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 3608 15104 3660 15156
rect 5724 15104 5776 15156
rect 4620 15036 4672 15088
rect 5448 15036 5500 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 2780 14968 2832 15020
rect 2964 14968 3016 15020
rect 2228 14900 2280 14952
rect 4068 14900 4120 14952
rect 4528 14900 4580 14952
rect 3240 14807 3292 14816
rect 3240 14773 3249 14807
rect 3249 14773 3283 14807
rect 3283 14773 3292 14807
rect 3240 14764 3292 14773
rect 3700 14764 3752 14816
rect 4252 14764 4304 14816
rect 4620 14764 4672 14816
rect 5080 15011 5132 15020
rect 5080 14977 5089 15011
rect 5089 14977 5123 15011
rect 5123 14977 5132 15011
rect 5080 14968 5132 14977
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 5356 14900 5408 14952
rect 6552 14968 6604 15020
rect 8300 15104 8352 15156
rect 7472 15036 7524 15088
rect 9220 15104 9272 15156
rect 9864 15104 9916 15156
rect 10876 15104 10928 15156
rect 11060 15104 11112 15156
rect 11796 15104 11848 15156
rect 12256 15104 12308 15156
rect 13636 15104 13688 15156
rect 13820 15104 13872 15156
rect 14280 15104 14332 15156
rect 14740 15104 14792 15156
rect 10048 15036 10100 15088
rect 11428 15036 11480 15088
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 9588 14900 9640 14952
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 13084 15036 13136 15088
rect 12440 14968 12492 15020
rect 12716 15011 12768 15020
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 12348 14900 12400 14952
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 13636 14900 13688 14952
rect 14832 15036 14884 15088
rect 15476 15036 15528 15088
rect 18788 15104 18840 15156
rect 19524 15104 19576 15156
rect 20260 15104 20312 15156
rect 22008 15104 22060 15156
rect 20720 15036 20772 15088
rect 21272 15036 21324 15088
rect 24952 15104 25004 15156
rect 28172 15104 28224 15156
rect 29460 15104 29512 15156
rect 30104 15147 30156 15156
rect 30104 15113 30113 15147
rect 30113 15113 30147 15147
rect 30147 15113 30156 15147
rect 30104 15104 30156 15113
rect 23848 15036 23900 15088
rect 27988 15036 28040 15088
rect 33140 15079 33192 15088
rect 33140 15045 33149 15079
rect 33149 15045 33183 15079
rect 33183 15045 33192 15079
rect 33140 15036 33192 15045
rect 34428 15036 34480 15088
rect 35992 15104 36044 15156
rect 37464 15036 37516 15088
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 17960 14968 18012 15020
rect 18696 15011 18748 15020
rect 18696 14977 18705 15011
rect 18705 14977 18739 15011
rect 18739 14977 18748 15011
rect 18696 14968 18748 14977
rect 18972 14968 19024 15020
rect 19156 14968 19208 15020
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 19432 14968 19484 14977
rect 18880 14900 18932 14952
rect 19708 14968 19760 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20352 15011 20404 15020
rect 20352 14977 20361 15011
rect 20361 14977 20395 15011
rect 20395 14977 20404 15011
rect 20352 14968 20404 14977
rect 20812 14900 20864 14952
rect 22100 14900 22152 14952
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 19248 14875 19300 14884
rect 19248 14841 19257 14875
rect 19257 14841 19291 14875
rect 19291 14841 19300 14875
rect 19248 14832 19300 14841
rect 19984 14832 20036 14884
rect 5816 14764 5868 14816
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 18788 14764 18840 14816
rect 18880 14764 18932 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 23204 14764 23256 14816
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 26792 14968 26844 15020
rect 29828 14968 29880 15020
rect 30748 14968 30800 15020
rect 32864 15011 32916 15020
rect 32864 14977 32873 15011
rect 32873 14977 32907 15011
rect 32907 14977 32916 15011
rect 32864 14968 32916 14977
rect 36636 15011 36688 15020
rect 36636 14977 36645 15011
rect 36645 14977 36679 15011
rect 36679 14977 36688 15011
rect 36636 14968 36688 14977
rect 24124 14900 24176 14952
rect 25504 14900 25556 14952
rect 27712 14900 27764 14952
rect 34796 14943 34848 14952
rect 34796 14909 34805 14943
rect 34805 14909 34839 14943
rect 34839 14909 34848 14943
rect 34796 14900 34848 14909
rect 35440 14900 35492 14952
rect 36084 14832 36136 14884
rect 24032 14764 24084 14816
rect 24676 14764 24728 14816
rect 31024 14764 31076 14816
rect 34612 14807 34664 14816
rect 34612 14773 34621 14807
rect 34621 14773 34655 14807
rect 34655 14773 34664 14807
rect 34612 14764 34664 14773
rect 36544 14807 36596 14816
rect 36544 14773 36553 14807
rect 36553 14773 36587 14807
rect 36587 14773 36596 14807
rect 36544 14764 36596 14773
rect 37280 14764 37332 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 4804 14560 4856 14612
rect 5264 14560 5316 14612
rect 9588 14603 9640 14612
rect 9588 14569 9597 14603
rect 9597 14569 9631 14603
rect 9631 14569 9640 14603
rect 9588 14560 9640 14569
rect 11152 14560 11204 14612
rect 11428 14603 11480 14612
rect 11428 14569 11437 14603
rect 11437 14569 11471 14603
rect 11471 14569 11480 14603
rect 11428 14560 11480 14569
rect 12348 14560 12400 14612
rect 13912 14560 13964 14612
rect 18052 14560 18104 14612
rect 19340 14560 19392 14612
rect 19984 14560 20036 14612
rect 20352 14560 20404 14612
rect 22468 14560 22520 14612
rect 24400 14560 24452 14612
rect 3240 14424 3292 14476
rect 3608 14467 3660 14476
rect 3608 14433 3617 14467
rect 3617 14433 3651 14467
rect 3651 14433 3660 14467
rect 3608 14424 3660 14433
rect 1860 14399 1912 14408
rect 1860 14365 1869 14399
rect 1869 14365 1903 14399
rect 1903 14365 1912 14399
rect 1860 14356 1912 14365
rect 2412 14399 2464 14408
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 3056 14356 3108 14408
rect 4620 14492 4672 14544
rect 4712 14492 4764 14544
rect 4804 14467 4856 14476
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 8668 14492 8720 14544
rect 4804 14424 4856 14433
rect 5724 14424 5776 14476
rect 10692 14424 10744 14476
rect 3884 14356 3936 14408
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 4068 14288 4120 14340
rect 5356 14288 5408 14340
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 11336 14424 11388 14476
rect 12164 14424 12216 14476
rect 12992 14535 13044 14544
rect 12992 14501 13001 14535
rect 13001 14501 13035 14535
rect 13035 14501 13044 14535
rect 12992 14492 13044 14501
rect 25044 14560 25096 14612
rect 25504 14603 25556 14612
rect 25504 14569 25513 14603
rect 25513 14569 25547 14603
rect 25547 14569 25556 14603
rect 25504 14560 25556 14569
rect 26976 14560 27028 14612
rect 13636 14467 13688 14476
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 11060 14399 11112 14408
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 11060 14356 11112 14365
rect 12624 14356 12676 14408
rect 13820 14356 13872 14408
rect 13912 14399 13964 14408
rect 13912 14365 13921 14399
rect 13921 14365 13955 14399
rect 13955 14365 13964 14399
rect 13912 14356 13964 14365
rect 16212 14356 16264 14408
rect 18788 14467 18840 14476
rect 18788 14433 18797 14467
rect 18797 14433 18831 14467
rect 18831 14433 18840 14467
rect 18788 14424 18840 14433
rect 23480 14424 23532 14476
rect 25228 14492 25280 14544
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 19064 14399 19116 14408
rect 19064 14365 19073 14399
rect 19073 14365 19107 14399
rect 19107 14365 19116 14399
rect 19064 14356 19116 14365
rect 19156 14356 19208 14408
rect 22100 14356 22152 14408
rect 24768 14424 24820 14476
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 26884 14467 26936 14476
rect 26884 14433 26893 14467
rect 26893 14433 26927 14467
rect 26927 14433 26936 14467
rect 26884 14424 26936 14433
rect 27620 14424 27672 14476
rect 2688 14220 2740 14272
rect 3332 14220 3384 14272
rect 6184 14331 6236 14340
rect 6184 14297 6193 14331
rect 6193 14297 6227 14331
rect 6227 14297 6236 14331
rect 6184 14288 6236 14297
rect 7472 14288 7524 14340
rect 10508 14288 10560 14340
rect 12808 14288 12860 14340
rect 14188 14331 14240 14340
rect 14188 14297 14197 14331
rect 14197 14297 14231 14331
rect 14231 14297 14240 14331
rect 14188 14288 14240 14297
rect 16948 14288 17000 14340
rect 18144 14288 18196 14340
rect 21088 14288 21140 14340
rect 7656 14263 7708 14272
rect 7656 14229 7665 14263
rect 7665 14229 7699 14263
rect 7699 14229 7708 14263
rect 7656 14220 7708 14229
rect 10232 14220 10284 14272
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 13636 14220 13688 14272
rect 14740 14220 14792 14272
rect 17040 14220 17092 14272
rect 17776 14220 17828 14272
rect 18696 14220 18748 14272
rect 21548 14331 21600 14340
rect 21548 14297 21557 14331
rect 21557 14297 21591 14331
rect 21591 14297 21600 14331
rect 21548 14288 21600 14297
rect 23572 14331 23624 14340
rect 23572 14297 23581 14331
rect 23581 14297 23615 14331
rect 23615 14297 23624 14331
rect 23572 14288 23624 14297
rect 24032 14356 24084 14408
rect 24216 14399 24268 14408
rect 24216 14365 24225 14399
rect 24225 14365 24259 14399
rect 24259 14365 24268 14399
rect 24216 14356 24268 14365
rect 24308 14356 24360 14408
rect 26240 14356 26292 14408
rect 26516 14399 26568 14408
rect 26516 14365 26525 14399
rect 26525 14365 26559 14399
rect 26559 14365 26568 14399
rect 26516 14356 26568 14365
rect 29828 14560 29880 14612
rect 30840 14560 30892 14612
rect 34520 14560 34572 14612
rect 35440 14560 35492 14612
rect 30932 14492 30984 14544
rect 32864 14492 32916 14544
rect 34612 14492 34664 14544
rect 29552 14467 29604 14476
rect 29552 14433 29561 14467
rect 29561 14433 29595 14467
rect 29595 14433 29604 14467
rect 29552 14424 29604 14433
rect 30196 14424 30248 14476
rect 34704 14467 34756 14476
rect 34704 14433 34713 14467
rect 34713 14433 34747 14467
rect 34747 14433 34756 14467
rect 34704 14424 34756 14433
rect 34796 14424 34848 14476
rect 29368 14399 29420 14408
rect 29368 14365 29377 14399
rect 29377 14365 29411 14399
rect 29411 14365 29420 14399
rect 29368 14356 29420 14365
rect 35072 14399 35124 14408
rect 35072 14365 35081 14399
rect 35081 14365 35115 14399
rect 35115 14365 35124 14399
rect 35072 14356 35124 14365
rect 35992 14356 36044 14408
rect 36360 14399 36412 14408
rect 36360 14365 36369 14399
rect 36369 14365 36403 14399
rect 36403 14365 36412 14399
rect 36360 14356 36412 14365
rect 36728 14399 36780 14408
rect 36728 14365 36737 14399
rect 36737 14365 36771 14399
rect 36771 14365 36780 14399
rect 36728 14356 36780 14365
rect 24676 14331 24728 14340
rect 24676 14297 24685 14331
rect 24685 14297 24719 14331
rect 24719 14297 24728 14331
rect 24676 14288 24728 14297
rect 27068 14288 27120 14340
rect 27896 14288 27948 14340
rect 31116 14288 31168 14340
rect 31208 14288 31260 14340
rect 22008 14220 22060 14272
rect 24952 14220 25004 14272
rect 27528 14220 27580 14272
rect 28632 14263 28684 14272
rect 28632 14229 28641 14263
rect 28641 14229 28675 14263
rect 28675 14229 28684 14263
rect 28632 14220 28684 14229
rect 31300 14220 31352 14272
rect 34796 14288 34848 14340
rect 36084 14288 36136 14340
rect 36636 14331 36688 14340
rect 36636 14297 36645 14331
rect 36645 14297 36679 14331
rect 36679 14297 36688 14331
rect 36636 14288 36688 14297
rect 37464 14288 37516 14340
rect 37372 14220 37424 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 3608 14016 3660 14068
rect 3976 14016 4028 14068
rect 5356 14059 5408 14068
rect 2780 13948 2832 14000
rect 3700 13991 3752 14000
rect 3700 13957 3709 13991
rect 3709 13957 3743 13991
rect 3743 13957 3752 13991
rect 3700 13948 3752 13957
rect 4344 13948 4396 14000
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 6184 14016 6236 14068
rect 11060 14016 11112 14068
rect 12900 14016 12952 14068
rect 13728 14059 13780 14068
rect 13728 14025 13737 14059
rect 13737 14025 13771 14059
rect 13771 14025 13780 14059
rect 13728 14016 13780 14025
rect 1400 13880 1452 13932
rect 5632 13991 5684 14000
rect 5632 13957 5641 13991
rect 5641 13957 5675 13991
rect 5675 13957 5684 13991
rect 5632 13948 5684 13957
rect 5356 13880 5408 13932
rect 6552 13880 6604 13932
rect 7656 13880 7708 13932
rect 8300 13948 8352 14000
rect 9956 13948 10008 14000
rect 10232 13880 10284 13932
rect 10508 13880 10560 13932
rect 2780 13812 2832 13864
rect 4160 13812 4212 13864
rect 3332 13676 3384 13728
rect 4804 13719 4856 13728
rect 4804 13685 4813 13719
rect 4813 13685 4847 13719
rect 4847 13685 4856 13719
rect 4804 13676 4856 13685
rect 4896 13676 4948 13728
rect 11060 13880 11112 13932
rect 11796 13880 11848 13932
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 12900 13923 12952 13932
rect 12900 13889 12909 13923
rect 12909 13889 12943 13923
rect 12943 13889 12952 13923
rect 12900 13880 12952 13889
rect 14832 13948 14884 14000
rect 5264 13676 5316 13728
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 10048 13744 10100 13796
rect 12992 13812 13044 13864
rect 13360 13880 13412 13932
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 17684 14016 17736 14068
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 17960 14016 18012 14068
rect 18880 14016 18932 14068
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 20168 14016 20220 14068
rect 17040 13880 17092 13932
rect 19340 13948 19392 14000
rect 19432 13991 19484 14000
rect 19432 13957 19457 13991
rect 19457 13957 19484 13991
rect 19432 13948 19484 13957
rect 13360 13787 13412 13796
rect 13360 13753 13369 13787
rect 13369 13753 13403 13787
rect 13403 13753 13412 13787
rect 13360 13744 13412 13753
rect 17592 13812 17644 13864
rect 17960 13855 18012 13864
rect 17960 13821 17969 13855
rect 17969 13821 18003 13855
rect 18003 13821 18012 13855
rect 17960 13812 18012 13821
rect 18696 13880 18748 13932
rect 20260 13948 20312 14000
rect 21548 14016 21600 14068
rect 24308 14016 24360 14068
rect 24768 14016 24820 14068
rect 27068 14059 27120 14068
rect 27068 14025 27077 14059
rect 27077 14025 27111 14059
rect 27111 14025 27120 14059
rect 27068 14016 27120 14025
rect 27528 14016 27580 14068
rect 29368 14016 29420 14068
rect 31024 14059 31076 14068
rect 31024 14025 31033 14059
rect 31033 14025 31067 14059
rect 31067 14025 31076 14059
rect 31024 14016 31076 14025
rect 31208 14059 31260 14068
rect 31208 14025 31217 14059
rect 31217 14025 31251 14059
rect 31251 14025 31260 14059
rect 31208 14016 31260 14025
rect 35992 14059 36044 14068
rect 35992 14025 36001 14059
rect 36001 14025 36035 14059
rect 36035 14025 36044 14059
rect 35992 14016 36044 14025
rect 36636 14016 36688 14068
rect 37372 14016 37424 14068
rect 19984 13923 20036 13932
rect 19984 13889 19993 13923
rect 19993 13889 20027 13923
rect 20027 13889 20036 13923
rect 19984 13880 20036 13889
rect 20444 13880 20496 13932
rect 22100 13948 22152 14000
rect 23848 13948 23900 14000
rect 19524 13812 19576 13864
rect 19616 13812 19668 13864
rect 23480 13880 23532 13932
rect 24676 13991 24728 14000
rect 24676 13957 24685 13991
rect 24685 13957 24719 13991
rect 24719 13957 24728 13991
rect 24676 13948 24728 13957
rect 29828 13991 29880 14000
rect 29828 13957 29837 13991
rect 29837 13957 29871 13991
rect 29871 13957 29880 13991
rect 29828 13948 29880 13957
rect 22100 13855 22152 13864
rect 22100 13821 22109 13855
rect 22109 13821 22143 13855
rect 22143 13821 22152 13855
rect 22100 13812 22152 13821
rect 26700 13880 26752 13932
rect 28632 13880 28684 13932
rect 12440 13676 12492 13728
rect 13176 13676 13228 13728
rect 13636 13676 13688 13728
rect 14004 13719 14056 13728
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 16580 13676 16632 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 20720 13744 20772 13796
rect 23940 13744 23992 13796
rect 24860 13812 24912 13864
rect 27804 13812 27856 13864
rect 28540 13812 28592 13864
rect 26516 13744 26568 13796
rect 28172 13744 28224 13796
rect 34612 13948 34664 14000
rect 30932 13880 30984 13932
rect 31668 13880 31720 13932
rect 33508 13923 33560 13932
rect 33508 13889 33517 13923
rect 33517 13889 33551 13923
rect 33551 13889 33560 13923
rect 33508 13880 33560 13889
rect 35440 13880 35492 13932
rect 19616 13719 19668 13728
rect 19616 13685 19625 13719
rect 19625 13685 19659 13719
rect 19659 13685 19668 13719
rect 19616 13676 19668 13685
rect 20536 13719 20588 13728
rect 20536 13685 20545 13719
rect 20545 13685 20579 13719
rect 20579 13685 20588 13719
rect 20536 13676 20588 13685
rect 23664 13676 23716 13728
rect 24952 13676 25004 13728
rect 30196 13676 30248 13728
rect 30656 13787 30708 13796
rect 30656 13753 30665 13787
rect 30665 13753 30699 13787
rect 30699 13753 30708 13787
rect 30656 13744 30708 13753
rect 31760 13744 31812 13796
rect 35072 13812 35124 13864
rect 36360 13948 36412 14000
rect 35992 13923 36044 13932
rect 35992 13889 36001 13923
rect 36001 13889 36035 13923
rect 36035 13889 36044 13923
rect 35992 13880 36044 13889
rect 36084 13923 36136 13932
rect 36084 13889 36093 13923
rect 36093 13889 36127 13923
rect 36127 13889 36136 13923
rect 36084 13880 36136 13889
rect 37280 13744 37332 13796
rect 31576 13676 31628 13728
rect 32864 13676 32916 13728
rect 34704 13676 34756 13728
rect 35440 13676 35492 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2780 13472 2832 13524
rect 1860 13336 1912 13388
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 3884 13472 3936 13524
rect 3976 13515 4028 13524
rect 3976 13481 3985 13515
rect 3985 13481 4019 13515
rect 4019 13481 4028 13515
rect 3976 13472 4028 13481
rect 4988 13472 5040 13524
rect 12992 13515 13044 13524
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 15476 13472 15528 13524
rect 17592 13472 17644 13524
rect 17684 13472 17736 13524
rect 19432 13472 19484 13524
rect 20168 13472 20220 13524
rect 20720 13472 20772 13524
rect 21088 13472 21140 13524
rect 21916 13515 21968 13524
rect 21916 13481 21925 13515
rect 21925 13481 21959 13515
rect 21959 13481 21968 13515
rect 21916 13472 21968 13481
rect 22100 13515 22152 13524
rect 22100 13481 22109 13515
rect 22109 13481 22143 13515
rect 22143 13481 22152 13515
rect 22100 13472 22152 13481
rect 24952 13472 25004 13524
rect 25228 13515 25280 13524
rect 25228 13481 25237 13515
rect 25237 13481 25271 13515
rect 25271 13481 25280 13515
rect 25228 13472 25280 13481
rect 29828 13472 29880 13524
rect 31300 13472 31352 13524
rect 35992 13472 36044 13524
rect 36176 13472 36228 13524
rect 9220 13404 9272 13456
rect 13728 13404 13780 13456
rect 4620 13336 4672 13388
rect 10048 13336 10100 13388
rect 12348 13336 12400 13388
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 12624 13336 12676 13388
rect 2504 13200 2556 13252
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 10232 13268 10284 13320
rect 12532 13268 12584 13320
rect 13452 13336 13504 13388
rect 14740 13379 14792 13388
rect 14740 13345 14749 13379
rect 14749 13345 14783 13379
rect 14783 13345 14792 13379
rect 14740 13336 14792 13345
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 16580 13336 16632 13388
rect 4528 13200 4580 13252
rect 4620 13243 4672 13252
rect 4620 13209 4629 13243
rect 4629 13209 4663 13243
rect 4663 13209 4672 13243
rect 4620 13200 4672 13209
rect 4804 13132 4856 13184
rect 5448 13132 5500 13184
rect 9128 13200 9180 13252
rect 10140 13200 10192 13252
rect 6920 13132 6972 13184
rect 7656 13175 7708 13184
rect 7656 13141 7665 13175
rect 7665 13141 7699 13175
rect 7699 13141 7708 13175
rect 7656 13132 7708 13141
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 9680 13132 9732 13184
rect 11428 13132 11480 13184
rect 11796 13200 11848 13252
rect 12808 13200 12860 13252
rect 13268 13268 13320 13320
rect 13360 13268 13412 13320
rect 13820 13311 13872 13320
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 13820 13268 13872 13277
rect 14004 13268 14056 13320
rect 15108 13268 15160 13320
rect 14464 13200 14516 13252
rect 16028 13268 16080 13320
rect 18420 13268 18472 13320
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 19616 13268 19668 13320
rect 20260 13379 20312 13388
rect 20260 13345 20269 13379
rect 20269 13345 20303 13379
rect 20303 13345 20312 13379
rect 20260 13336 20312 13345
rect 24216 13404 24268 13456
rect 27896 13404 27948 13456
rect 28632 13404 28684 13456
rect 23940 13379 23992 13388
rect 20168 13268 20220 13320
rect 21548 13268 21600 13320
rect 23940 13345 23949 13379
rect 23949 13345 23983 13379
rect 23983 13345 23992 13379
rect 23940 13336 23992 13345
rect 23388 13268 23440 13320
rect 12440 13132 12492 13184
rect 12992 13132 13044 13184
rect 17684 13200 17736 13252
rect 18144 13200 18196 13252
rect 21180 13200 21232 13252
rect 21640 13200 21692 13252
rect 23664 13268 23716 13320
rect 24216 13268 24268 13320
rect 24952 13336 25004 13388
rect 28172 13336 28224 13388
rect 30380 13336 30432 13388
rect 32772 13336 32824 13388
rect 35992 13336 36044 13388
rect 36728 13379 36780 13388
rect 36728 13345 36737 13379
rect 36737 13345 36771 13379
rect 36771 13345 36780 13379
rect 36728 13336 36780 13345
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 23756 13200 23808 13252
rect 25136 13311 25188 13320
rect 25136 13277 25145 13311
rect 25145 13277 25179 13311
rect 25179 13277 25188 13311
rect 25136 13268 25188 13277
rect 26516 13311 26568 13320
rect 26516 13277 26525 13311
rect 26525 13277 26559 13311
rect 26559 13277 26568 13311
rect 26516 13268 26568 13277
rect 26608 13268 26660 13320
rect 14832 13175 14884 13184
rect 14832 13141 14841 13175
rect 14841 13141 14875 13175
rect 14875 13141 14884 13175
rect 14832 13132 14884 13141
rect 18696 13175 18748 13184
rect 18696 13141 18705 13175
rect 18705 13141 18739 13175
rect 18739 13141 18748 13175
rect 18696 13132 18748 13141
rect 19892 13175 19944 13184
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 23112 13175 23164 13184
rect 23112 13141 23121 13175
rect 23121 13141 23155 13175
rect 23155 13141 23164 13175
rect 23112 13132 23164 13141
rect 26700 13243 26752 13252
rect 26700 13209 26709 13243
rect 26709 13209 26743 13243
rect 26743 13209 26752 13243
rect 26700 13200 26752 13209
rect 27620 13243 27672 13252
rect 27620 13209 27629 13243
rect 27629 13209 27663 13243
rect 27663 13209 27672 13243
rect 27620 13200 27672 13209
rect 28632 13311 28684 13320
rect 28632 13277 28641 13311
rect 28641 13277 28675 13311
rect 28675 13277 28684 13311
rect 28632 13268 28684 13277
rect 34336 13268 34388 13320
rect 28724 13200 28776 13252
rect 29092 13200 29144 13252
rect 31116 13200 31168 13252
rect 31300 13200 31352 13252
rect 32864 13200 32916 13252
rect 26884 13132 26936 13184
rect 28264 13132 28316 13184
rect 29736 13175 29788 13184
rect 29736 13141 29745 13175
rect 29745 13141 29779 13175
rect 29779 13141 29788 13175
rect 29736 13132 29788 13141
rect 31208 13132 31260 13184
rect 33508 13132 33560 13184
rect 34704 13200 34756 13252
rect 37004 13243 37056 13252
rect 37004 13209 37013 13243
rect 37013 13209 37047 13243
rect 37047 13209 37056 13243
rect 37004 13200 37056 13209
rect 37464 13200 37516 13252
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 4528 12928 4580 12980
rect 4620 12928 4672 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 5540 12928 5592 12980
rect 9588 12928 9640 12980
rect 2780 12903 2832 12912
rect 2780 12869 2789 12903
rect 2789 12869 2823 12903
rect 2823 12869 2832 12903
rect 2780 12860 2832 12869
rect 4160 12860 4212 12912
rect 5448 12860 5500 12912
rect 6920 12903 6972 12912
rect 6920 12869 6929 12903
rect 6929 12869 6963 12903
rect 6963 12869 6972 12903
rect 6920 12860 6972 12869
rect 7472 12860 7524 12912
rect 9680 12903 9732 12912
rect 9680 12869 9689 12903
rect 9689 12869 9723 12903
rect 9723 12869 9732 12903
rect 9680 12860 9732 12869
rect 10140 12860 10192 12912
rect 12532 12928 12584 12980
rect 12900 12928 12952 12980
rect 19156 12928 19208 12980
rect 21548 12971 21600 12980
rect 21548 12937 21557 12971
rect 21557 12937 21591 12971
rect 21591 12937 21600 12971
rect 21548 12928 21600 12937
rect 21640 12928 21692 12980
rect 27620 12928 27672 12980
rect 28632 12928 28684 12980
rect 28816 12971 28868 12980
rect 28816 12937 28825 12971
rect 28825 12937 28859 12971
rect 28859 12937 28868 12971
rect 28816 12928 28868 12937
rect 30656 12971 30708 12980
rect 30656 12937 30665 12971
rect 30665 12937 30699 12971
rect 30699 12937 30708 12971
rect 30656 12928 30708 12937
rect 31116 12971 31168 12980
rect 31116 12937 31125 12971
rect 31125 12937 31159 12971
rect 31159 12937 31168 12971
rect 31116 12928 31168 12937
rect 31300 12928 31352 12980
rect 33416 12928 33468 12980
rect 35440 12928 35492 12980
rect 36360 12928 36412 12980
rect 12440 12860 12492 12912
rect 14924 12860 14976 12912
rect 15752 12860 15804 12912
rect 4620 12792 4672 12844
rect 4804 12792 4856 12844
rect 5264 12792 5316 12844
rect 5908 12792 5960 12844
rect 6184 12792 6236 12844
rect 8300 12792 8352 12844
rect 11428 12792 11480 12844
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 13544 12792 13596 12844
rect 17408 12860 17460 12912
rect 18052 12860 18104 12912
rect 16580 12792 16632 12844
rect 19432 12792 19484 12844
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 21088 12792 21140 12844
rect 23848 12792 23900 12844
rect 24952 12860 25004 12912
rect 26424 12903 26476 12912
rect 26424 12869 26433 12903
rect 26433 12869 26467 12903
rect 26467 12869 26476 12903
rect 26424 12860 26476 12869
rect 26700 12860 26752 12912
rect 27528 12860 27580 12912
rect 27896 12860 27948 12912
rect 29828 12860 29880 12912
rect 30380 12860 30432 12912
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 24676 12792 24728 12844
rect 25136 12792 25188 12844
rect 26516 12792 26568 12844
rect 26608 12835 26660 12844
rect 26608 12801 26617 12835
rect 26617 12801 26651 12835
rect 26651 12801 26660 12835
rect 26608 12792 26660 12801
rect 33232 12860 33284 12912
rect 37004 12971 37056 12980
rect 37004 12937 37013 12971
rect 37013 12937 37047 12971
rect 37047 12937 37056 12971
rect 37004 12928 37056 12937
rect 2504 12767 2556 12776
rect 2504 12733 2513 12767
rect 2513 12733 2547 12767
rect 2547 12733 2556 12767
rect 2504 12724 2556 12733
rect 4988 12724 5040 12776
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 14096 12767 14148 12776
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 20444 12724 20496 12776
rect 4804 12656 4856 12708
rect 8484 12656 8536 12708
rect 7472 12588 7524 12640
rect 8024 12588 8076 12640
rect 8576 12588 8628 12640
rect 19616 12656 19668 12708
rect 20260 12656 20312 12708
rect 20812 12656 20864 12708
rect 26240 12724 26292 12776
rect 27252 12767 27304 12776
rect 27252 12733 27261 12767
rect 27261 12733 27295 12767
rect 27295 12733 27304 12767
rect 27252 12724 27304 12733
rect 28540 12724 28592 12776
rect 10140 12588 10192 12640
rect 13452 12631 13504 12640
rect 13452 12597 13461 12631
rect 13461 12597 13495 12631
rect 13495 12597 13504 12631
rect 13452 12588 13504 12597
rect 19340 12631 19392 12640
rect 19340 12597 19349 12631
rect 19349 12597 19383 12631
rect 19383 12597 19392 12631
rect 19340 12588 19392 12597
rect 23480 12588 23532 12640
rect 26792 12631 26844 12640
rect 26792 12597 26801 12631
rect 26801 12597 26835 12631
rect 26835 12597 26844 12631
rect 26792 12588 26844 12597
rect 28724 12631 28776 12640
rect 28724 12597 28733 12631
rect 28733 12597 28767 12631
rect 28767 12597 28776 12631
rect 28724 12588 28776 12597
rect 30196 12588 30248 12640
rect 31116 12792 31168 12844
rect 31484 12835 31536 12844
rect 31484 12801 31493 12835
rect 31493 12801 31527 12835
rect 31527 12801 31536 12835
rect 31484 12792 31536 12801
rect 31576 12835 31628 12844
rect 31576 12801 31585 12835
rect 31585 12801 31619 12835
rect 31619 12801 31628 12835
rect 31576 12792 31628 12801
rect 31760 12835 31812 12844
rect 31760 12801 31769 12835
rect 31769 12801 31803 12835
rect 31803 12801 31812 12835
rect 31760 12792 31812 12801
rect 36084 12835 36136 12844
rect 36084 12801 36093 12835
rect 36093 12801 36127 12835
rect 36127 12801 36136 12835
rect 36084 12792 36136 12801
rect 36176 12835 36228 12844
rect 36176 12801 36185 12835
rect 36185 12801 36219 12835
rect 36219 12801 36228 12835
rect 36176 12792 36228 12801
rect 31208 12724 31260 12776
rect 32680 12699 32732 12708
rect 32680 12665 32689 12699
rect 32689 12665 32723 12699
rect 32723 12665 32732 12699
rect 32680 12656 32732 12665
rect 31300 12588 31352 12640
rect 34612 12656 34664 12708
rect 36268 12724 36320 12776
rect 36636 12835 36688 12844
rect 36636 12801 36645 12835
rect 36645 12801 36679 12835
rect 36679 12801 36688 12835
rect 36636 12792 36688 12801
rect 37004 12724 37056 12776
rect 37280 12767 37332 12776
rect 37280 12733 37289 12767
rect 37289 12733 37323 12767
rect 37323 12733 37332 12767
rect 37280 12724 37332 12733
rect 33140 12588 33192 12640
rect 36636 12588 36688 12640
rect 37832 12588 37884 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4712 12316 4764 12368
rect 5172 12384 5224 12436
rect 9128 12384 9180 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 13084 12384 13136 12436
rect 13360 12384 13412 12436
rect 15292 12384 15344 12436
rect 15660 12384 15712 12436
rect 5816 12359 5868 12368
rect 5816 12325 5825 12359
rect 5825 12325 5859 12359
rect 5859 12325 5868 12359
rect 5816 12316 5868 12325
rect 4804 12248 4856 12300
rect 10876 12316 10928 12368
rect 11244 12316 11296 12368
rect 7656 12248 7708 12300
rect 8116 12248 8168 12300
rect 13452 12316 13504 12368
rect 17132 12384 17184 12436
rect 20812 12384 20864 12436
rect 25136 12384 25188 12436
rect 26884 12384 26936 12436
rect 27252 12384 27304 12436
rect 28264 12384 28316 12436
rect 4344 12180 4396 12232
rect 3424 12112 3476 12164
rect 4436 12112 4488 12164
rect 5172 12180 5224 12232
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 7748 12180 7800 12232
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4528 12044 4580 12096
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 6460 12155 6512 12164
rect 6460 12121 6469 12155
rect 6469 12121 6503 12155
rect 6503 12121 6512 12155
rect 6460 12112 6512 12121
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 5356 12044 5408 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 8392 12044 8444 12096
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 12808 12248 12860 12300
rect 13728 12248 13780 12300
rect 13176 12180 13228 12232
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 8852 12044 8904 12096
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 13912 12112 13964 12164
rect 11612 12044 11664 12053
rect 11888 12087 11940 12096
rect 11888 12053 11897 12087
rect 11897 12053 11931 12087
rect 11931 12053 11940 12087
rect 11888 12044 11940 12053
rect 12256 12044 12308 12096
rect 12808 12044 12860 12096
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 13544 12044 13596 12096
rect 13728 12044 13780 12096
rect 15292 12180 15344 12232
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 18696 12248 18748 12300
rect 19616 12291 19668 12300
rect 19616 12257 19625 12291
rect 19625 12257 19659 12291
rect 19659 12257 19668 12291
rect 19616 12248 19668 12257
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 23480 12248 23532 12300
rect 19156 12180 19208 12232
rect 16948 12112 17000 12164
rect 18604 12112 18656 12164
rect 19064 12112 19116 12164
rect 20720 12180 20772 12232
rect 23388 12223 23440 12232
rect 23388 12189 23397 12223
rect 23397 12189 23431 12223
rect 23431 12189 23440 12223
rect 23388 12180 23440 12189
rect 24492 12316 24544 12368
rect 28540 12316 28592 12368
rect 23756 12180 23808 12232
rect 23940 12223 23992 12232
rect 23940 12189 23949 12223
rect 23949 12189 23983 12223
rect 23983 12189 23992 12223
rect 23940 12180 23992 12189
rect 24952 12248 25004 12300
rect 18420 12044 18472 12096
rect 20352 12044 20404 12096
rect 22008 12044 22060 12096
rect 23204 12044 23256 12096
rect 23848 12112 23900 12164
rect 24124 12155 24176 12164
rect 24124 12121 24133 12155
rect 24133 12121 24167 12155
rect 24167 12121 24176 12155
rect 24124 12112 24176 12121
rect 24676 12223 24728 12232
rect 24676 12189 24685 12223
rect 24685 12189 24719 12223
rect 24719 12189 24728 12223
rect 24676 12180 24728 12189
rect 24584 12112 24636 12164
rect 26516 12180 26568 12232
rect 30196 12384 30248 12436
rect 28724 12316 28776 12368
rect 28816 12359 28868 12368
rect 28816 12325 28825 12359
rect 28825 12325 28859 12359
rect 28859 12325 28868 12359
rect 28816 12316 28868 12325
rect 29828 12359 29880 12368
rect 29828 12325 29837 12359
rect 29837 12325 29871 12359
rect 29871 12325 29880 12359
rect 29828 12316 29880 12325
rect 24492 12087 24544 12096
rect 24492 12053 24501 12087
rect 24501 12053 24535 12087
rect 24535 12053 24544 12087
rect 24492 12044 24544 12053
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 25688 12087 25740 12096
rect 25688 12053 25697 12087
rect 25697 12053 25731 12087
rect 25731 12053 25740 12087
rect 25688 12044 25740 12053
rect 26792 12155 26844 12164
rect 26792 12121 26817 12155
rect 26817 12121 26844 12155
rect 26792 12112 26844 12121
rect 27528 12112 27580 12164
rect 29736 12180 29788 12232
rect 31208 12384 31260 12436
rect 33508 12384 33560 12436
rect 36268 12384 36320 12436
rect 31392 12316 31444 12368
rect 32680 12359 32732 12368
rect 32680 12325 32689 12359
rect 32689 12325 32723 12359
rect 32723 12325 32732 12359
rect 32680 12316 32732 12325
rect 32772 12291 32824 12300
rect 32772 12257 32781 12291
rect 32781 12257 32815 12291
rect 32815 12257 32824 12291
rect 32772 12248 32824 12257
rect 33140 12248 33192 12300
rect 33416 12248 33468 12300
rect 36084 12316 36136 12368
rect 36544 12316 36596 12368
rect 28356 12087 28408 12096
rect 28356 12053 28365 12087
rect 28365 12053 28399 12087
rect 28399 12053 28408 12087
rect 28356 12044 28408 12053
rect 30748 12223 30800 12232
rect 30748 12189 30757 12223
rect 30757 12189 30791 12223
rect 30791 12189 30800 12223
rect 30748 12180 30800 12189
rect 30932 12180 30984 12232
rect 31760 12223 31812 12232
rect 31760 12189 31769 12223
rect 31769 12189 31803 12223
rect 31803 12189 31812 12223
rect 31760 12180 31812 12189
rect 30840 12044 30892 12096
rect 31024 12112 31076 12164
rect 31300 12155 31352 12164
rect 31300 12121 31325 12155
rect 31325 12121 31352 12155
rect 31300 12112 31352 12121
rect 32772 12112 32824 12164
rect 34336 12112 34388 12164
rect 37464 12248 37516 12300
rect 35992 12180 36044 12232
rect 36544 12180 36596 12232
rect 31208 12044 31260 12096
rect 31668 12044 31720 12096
rect 35348 12044 35400 12096
rect 36360 12044 36412 12096
rect 36452 12087 36504 12096
rect 36452 12053 36461 12087
rect 36461 12053 36495 12087
rect 36495 12053 36504 12087
rect 36452 12044 36504 12053
rect 37096 12180 37148 12232
rect 36820 12112 36872 12164
rect 37004 12044 37056 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 4436 11883 4488 11892
rect 4436 11849 4445 11883
rect 4445 11849 4479 11883
rect 4479 11849 4488 11883
rect 4436 11840 4488 11849
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 3700 11704 3752 11756
rect 7748 11840 7800 11892
rect 8208 11840 8260 11892
rect 5448 11772 5500 11824
rect 7012 11772 7064 11824
rect 8392 11772 8444 11824
rect 9772 11840 9824 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 10048 11772 10100 11824
rect 4344 11679 4396 11688
rect 4344 11645 4353 11679
rect 4353 11645 4387 11679
rect 4387 11645 4396 11679
rect 4344 11636 4396 11645
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 6184 11679 6236 11688
rect 6184 11645 6193 11679
rect 6193 11645 6227 11679
rect 6227 11645 6236 11679
rect 6184 11636 6236 11645
rect 6552 11636 6604 11688
rect 7840 11679 7892 11688
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 12900 11840 12952 11892
rect 13084 11840 13136 11892
rect 11888 11772 11940 11824
rect 16948 11772 17000 11824
rect 17684 11840 17736 11892
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 20444 11840 20496 11892
rect 23940 11840 23992 11892
rect 33232 11883 33284 11892
rect 33232 11849 33241 11883
rect 33241 11849 33275 11883
rect 33275 11849 33284 11883
rect 33232 11840 33284 11849
rect 34796 11840 34848 11892
rect 23388 11772 23440 11824
rect 13728 11704 13780 11756
rect 13912 11704 13964 11756
rect 3424 11611 3476 11620
rect 3424 11577 3433 11611
rect 3433 11577 3467 11611
rect 3467 11577 3476 11611
rect 3424 11568 3476 11577
rect 4528 11568 4580 11620
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3608 11500 3660 11552
rect 4712 11500 4764 11552
rect 4804 11500 4856 11552
rect 12808 11636 12860 11688
rect 14096 11636 14148 11688
rect 20352 11704 20404 11756
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 23480 11704 23532 11756
rect 29736 11772 29788 11824
rect 35348 11772 35400 11824
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 17408 11636 17460 11688
rect 17500 11636 17552 11688
rect 18604 11679 18656 11688
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 19340 11636 19392 11688
rect 24676 11747 24728 11756
rect 24676 11713 24685 11747
rect 24685 11713 24719 11747
rect 24719 11713 24728 11747
rect 24676 11704 24728 11713
rect 13820 11611 13872 11620
rect 13820 11577 13829 11611
rect 13829 11577 13863 11611
rect 13863 11577 13872 11611
rect 13820 11568 13872 11577
rect 11612 11543 11664 11552
rect 11612 11509 11621 11543
rect 11621 11509 11655 11543
rect 11655 11509 11664 11543
rect 11612 11500 11664 11509
rect 12624 11500 12676 11552
rect 12900 11500 12952 11552
rect 21456 11568 21508 11620
rect 24308 11636 24360 11688
rect 25688 11704 25740 11756
rect 25964 11747 26016 11756
rect 25964 11713 25973 11747
rect 25973 11713 26007 11747
rect 26007 11713 26016 11747
rect 25964 11704 26016 11713
rect 26148 11747 26200 11756
rect 26148 11713 26157 11747
rect 26157 11713 26191 11747
rect 26191 11713 26200 11747
rect 26148 11704 26200 11713
rect 26240 11747 26292 11756
rect 26240 11713 26249 11747
rect 26249 11713 26283 11747
rect 26283 11713 26292 11747
rect 26240 11704 26292 11713
rect 26424 11704 26476 11756
rect 26608 11704 26660 11756
rect 26976 11747 27028 11756
rect 26976 11713 26985 11747
rect 26985 11713 27019 11747
rect 27019 11713 27028 11747
rect 26976 11704 27028 11713
rect 31024 11704 31076 11756
rect 31484 11704 31536 11756
rect 34796 11704 34848 11756
rect 36452 11772 36504 11824
rect 36728 11772 36780 11824
rect 31392 11636 31444 11688
rect 32772 11679 32824 11688
rect 32772 11645 32781 11679
rect 32781 11645 32815 11679
rect 32815 11645 32824 11679
rect 32772 11636 32824 11645
rect 23112 11568 23164 11620
rect 26608 11568 26660 11620
rect 26976 11568 27028 11620
rect 31576 11568 31628 11620
rect 33232 11636 33284 11688
rect 35716 11747 35768 11756
rect 35716 11713 35725 11747
rect 35725 11713 35759 11747
rect 35759 11713 35768 11747
rect 35716 11704 35768 11713
rect 36360 11704 36412 11756
rect 36176 11636 36228 11688
rect 36636 11679 36688 11688
rect 36636 11645 36645 11679
rect 36645 11645 36679 11679
rect 36679 11645 36688 11679
rect 36636 11636 36688 11645
rect 33600 11568 33652 11620
rect 35348 11611 35400 11620
rect 35348 11577 35357 11611
rect 35357 11577 35391 11611
rect 35391 11577 35400 11611
rect 35348 11568 35400 11577
rect 37832 11611 37884 11620
rect 37832 11577 37841 11611
rect 37841 11577 37875 11611
rect 37875 11577 37884 11611
rect 37832 11568 37884 11577
rect 21272 11500 21324 11552
rect 22284 11543 22336 11552
rect 22284 11509 22293 11543
rect 22293 11509 22327 11543
rect 22327 11509 22336 11543
rect 22284 11500 22336 11509
rect 24584 11500 24636 11552
rect 25044 11500 25096 11552
rect 28264 11500 28316 11552
rect 32680 11500 32732 11552
rect 34428 11500 34480 11552
rect 36544 11500 36596 11552
rect 36912 11500 36964 11552
rect 37372 11500 37424 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2504 11228 2556 11280
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 3608 11203 3660 11212
rect 3608 11169 3617 11203
rect 3617 11169 3651 11203
rect 3651 11169 3660 11203
rect 3608 11160 3660 11169
rect 1308 11092 1360 11144
rect 4620 11296 4672 11348
rect 5356 11296 5408 11348
rect 6460 11296 6512 11348
rect 5264 11228 5316 11280
rect 4160 11160 4212 11212
rect 4804 11160 4856 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 5908 11160 5960 11212
rect 7840 11228 7892 11280
rect 7380 11203 7432 11212
rect 7380 11169 7389 11203
rect 7389 11169 7423 11203
rect 7423 11169 7432 11203
rect 7380 11160 7432 11169
rect 8116 11160 8168 11212
rect 12624 11228 12676 11280
rect 17040 11296 17092 11348
rect 17132 11296 17184 11348
rect 17408 11339 17460 11348
rect 17408 11305 17417 11339
rect 17417 11305 17451 11339
rect 17451 11305 17460 11339
rect 17408 11296 17460 11305
rect 17684 11296 17736 11348
rect 3700 11024 3752 11076
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 8668 11092 8720 11144
rect 9036 11092 9088 11144
rect 11888 11092 11940 11144
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 12808 11160 12860 11169
rect 13176 11160 13228 11212
rect 14924 11160 14976 11212
rect 16672 11160 16724 11212
rect 17592 11160 17644 11212
rect 21824 11296 21876 11348
rect 13360 11092 13412 11144
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 15476 11092 15528 11144
rect 17776 11092 17828 11144
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 4068 11024 4120 11076
rect 14372 11067 14424 11076
rect 14372 11033 14381 11067
rect 14381 11033 14415 11067
rect 14415 11033 14424 11067
rect 14372 11024 14424 11033
rect 16212 11024 16264 11076
rect 16580 11024 16632 11076
rect 17040 11024 17092 11076
rect 18788 11135 18840 11144
rect 18788 11101 18797 11135
rect 18797 11101 18831 11135
rect 18831 11101 18840 11135
rect 18788 11092 18840 11101
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 24216 11092 24268 11144
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 24860 11135 24912 11144
rect 24860 11101 24869 11135
rect 24869 11101 24903 11135
rect 24903 11101 24912 11135
rect 24860 11092 24912 11101
rect 20996 11024 21048 11076
rect 24124 11024 24176 11076
rect 25964 11339 26016 11348
rect 25964 11305 25973 11339
rect 25973 11305 26007 11339
rect 26007 11305 26016 11339
rect 25964 11296 26016 11305
rect 30196 11296 30248 11348
rect 31760 11296 31812 11348
rect 28264 11203 28316 11212
rect 28264 11169 28273 11203
rect 28273 11169 28307 11203
rect 28307 11169 28316 11203
rect 28264 11160 28316 11169
rect 28540 11203 28592 11212
rect 28540 11169 28549 11203
rect 28549 11169 28583 11203
rect 28583 11169 28592 11203
rect 30932 11228 30984 11280
rect 28540 11160 28592 11169
rect 25964 11092 26016 11144
rect 26240 11135 26292 11144
rect 26240 11101 26249 11135
rect 26249 11101 26283 11135
rect 26283 11101 26292 11135
rect 26240 11092 26292 11101
rect 26332 11092 26384 11144
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 27804 11135 27856 11144
rect 27804 11101 27813 11135
rect 27813 11101 27847 11135
rect 27847 11101 27856 11135
rect 27804 11092 27856 11101
rect 27896 11135 27948 11144
rect 27896 11101 27905 11135
rect 27905 11101 27939 11135
rect 27939 11101 27948 11135
rect 27896 11092 27948 11101
rect 28816 11092 28868 11144
rect 32864 11296 32916 11348
rect 33600 11296 33652 11348
rect 36084 11339 36136 11348
rect 36084 11305 36093 11339
rect 36093 11305 36127 11339
rect 36127 11305 36136 11339
rect 36084 11296 36136 11305
rect 36176 11339 36228 11348
rect 36176 11305 36185 11339
rect 36185 11305 36219 11339
rect 36219 11305 36228 11339
rect 36176 11296 36228 11305
rect 36268 11339 36320 11348
rect 36268 11305 36277 11339
rect 36277 11305 36311 11339
rect 36311 11305 36320 11339
rect 36268 11296 36320 11305
rect 37096 11296 37148 11348
rect 30012 11135 30064 11144
rect 30012 11101 30021 11135
rect 30021 11101 30055 11135
rect 30055 11101 30064 11135
rect 30012 11092 30064 11101
rect 30104 11135 30156 11144
rect 30104 11101 30113 11135
rect 30113 11101 30147 11135
rect 30147 11101 30156 11135
rect 30104 11092 30156 11101
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 29092 11024 29144 11076
rect 29184 11067 29236 11076
rect 29184 11033 29193 11067
rect 29193 11033 29227 11067
rect 29227 11033 29236 11067
rect 29184 11024 29236 11033
rect 31024 11092 31076 11144
rect 32864 11135 32916 11144
rect 32864 11101 32873 11135
rect 32873 11101 32907 11135
rect 32907 11101 32916 11135
rect 32864 11092 32916 11101
rect 32956 11135 33008 11144
rect 32956 11101 32965 11135
rect 32965 11101 32999 11135
rect 32999 11101 33008 11135
rect 32956 11092 33008 11101
rect 33232 11135 33284 11144
rect 33232 11101 33241 11135
rect 33241 11101 33275 11135
rect 33275 11101 33284 11135
rect 33232 11092 33284 11101
rect 33876 11092 33928 11144
rect 36912 11203 36964 11212
rect 36912 11169 36921 11203
rect 36921 11169 36955 11203
rect 36955 11169 36964 11203
rect 36912 11160 36964 11169
rect 37004 11160 37056 11212
rect 30932 11024 30984 11076
rect 4804 10956 4856 11008
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 17776 10999 17828 11008
rect 17776 10965 17785 10999
rect 17785 10965 17819 10999
rect 17819 10965 17828 10999
rect 17776 10956 17828 10965
rect 17960 10956 18012 11008
rect 18420 10956 18472 11008
rect 22744 10956 22796 11008
rect 26332 10956 26384 11008
rect 28080 10956 28132 11008
rect 30104 10956 30156 11008
rect 30472 10956 30524 11008
rect 30656 10956 30708 11008
rect 32588 10999 32640 11008
rect 32588 10965 32597 10999
rect 32597 10965 32631 10999
rect 32631 10965 32640 10999
rect 32588 10956 32640 10965
rect 33324 10956 33376 11008
rect 34796 10956 34848 11008
rect 36268 11092 36320 11144
rect 36636 11135 36688 11144
rect 36636 11101 36645 11135
rect 36645 11101 36679 11135
rect 36679 11101 36688 11135
rect 36636 11092 36688 11101
rect 36084 11024 36136 11076
rect 37464 11024 37516 11076
rect 36176 10956 36228 11008
rect 36452 10956 36504 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 3700 10752 3752 10804
rect 1308 10616 1360 10668
rect 1584 10616 1636 10668
rect 2872 10684 2924 10736
rect 8484 10752 8536 10804
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 13636 10752 13688 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 14924 10752 14976 10804
rect 22284 10795 22336 10804
rect 22284 10761 22293 10795
rect 22293 10761 22327 10795
rect 22327 10761 22336 10795
rect 22284 10752 22336 10761
rect 22928 10752 22980 10804
rect 23296 10752 23348 10804
rect 8208 10684 8260 10736
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 3884 10616 3936 10668
rect 5356 10616 5408 10668
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 8300 10616 8352 10668
rect 8852 10616 8904 10668
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 11336 10684 11388 10736
rect 18328 10684 18380 10736
rect 20996 10684 21048 10736
rect 13360 10616 13412 10668
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 14648 10616 14700 10668
rect 17224 10616 17276 10668
rect 17592 10616 17644 10668
rect 4160 10548 4212 10600
rect 4712 10548 4764 10600
rect 8760 10548 8812 10600
rect 10968 10548 11020 10600
rect 15292 10548 15344 10600
rect 18144 10548 18196 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 20720 10548 20772 10600
rect 10324 10480 10376 10532
rect 22928 10659 22980 10668
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 24124 10684 24176 10736
rect 24860 10752 24912 10804
rect 29184 10795 29236 10804
rect 29184 10761 29193 10795
rect 29193 10761 29227 10795
rect 29227 10761 29236 10795
rect 29184 10752 29236 10761
rect 30196 10752 30248 10804
rect 33140 10752 33192 10804
rect 33968 10752 34020 10804
rect 34704 10752 34756 10804
rect 35348 10752 35400 10804
rect 36728 10752 36780 10804
rect 25688 10684 25740 10736
rect 23204 10659 23256 10668
rect 23204 10625 23213 10659
rect 23213 10625 23247 10659
rect 23247 10625 23256 10659
rect 23204 10616 23256 10625
rect 23480 10616 23532 10668
rect 23756 10616 23808 10668
rect 24308 10659 24360 10668
rect 24308 10625 24317 10659
rect 24317 10625 24351 10659
rect 24351 10625 24360 10659
rect 24308 10616 24360 10625
rect 25780 10659 25832 10668
rect 25780 10625 25789 10659
rect 25789 10625 25823 10659
rect 25823 10625 25832 10659
rect 25780 10616 25832 10625
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 26424 10659 26476 10668
rect 26424 10625 26433 10659
rect 26433 10625 26467 10659
rect 26467 10625 26476 10659
rect 26424 10616 26476 10625
rect 28540 10684 28592 10736
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 22468 10548 22520 10557
rect 22744 10523 22796 10532
rect 22744 10489 22753 10523
rect 22753 10489 22787 10523
rect 22787 10489 22796 10523
rect 22744 10480 22796 10489
rect 24584 10548 24636 10600
rect 26056 10548 26108 10600
rect 29000 10659 29052 10668
rect 29000 10625 29009 10659
rect 29009 10625 29043 10659
rect 29043 10625 29052 10659
rect 29000 10616 29052 10625
rect 30104 10616 30156 10668
rect 30472 10659 30524 10668
rect 30472 10625 30481 10659
rect 30481 10625 30515 10659
rect 30515 10625 30524 10659
rect 30472 10616 30524 10625
rect 30656 10659 30708 10668
rect 30656 10625 30665 10659
rect 30665 10625 30699 10659
rect 30699 10625 30708 10659
rect 30656 10616 30708 10625
rect 32956 10684 33008 10736
rect 30840 10659 30892 10668
rect 30840 10625 30849 10659
rect 30849 10625 30883 10659
rect 30883 10625 30892 10659
rect 30840 10616 30892 10625
rect 31024 10659 31076 10668
rect 31024 10625 31033 10659
rect 31033 10625 31067 10659
rect 31067 10625 31076 10659
rect 31024 10616 31076 10625
rect 29092 10548 29144 10600
rect 30012 10591 30064 10600
rect 30012 10557 30021 10591
rect 30021 10557 30055 10591
rect 30055 10557 30064 10591
rect 30012 10548 30064 10557
rect 30288 10548 30340 10600
rect 31116 10548 31168 10600
rect 32588 10548 32640 10600
rect 33140 10616 33192 10668
rect 33324 10659 33376 10668
rect 33324 10625 33333 10659
rect 33333 10625 33367 10659
rect 33367 10625 33376 10659
rect 33324 10616 33376 10625
rect 33600 10659 33652 10668
rect 33600 10625 33609 10659
rect 33609 10625 33643 10659
rect 33643 10625 33652 10659
rect 33600 10616 33652 10625
rect 33876 10659 33928 10668
rect 33876 10625 33885 10659
rect 33885 10625 33919 10659
rect 33919 10625 33928 10659
rect 33876 10616 33928 10625
rect 34520 10659 34572 10668
rect 34520 10625 34529 10659
rect 34529 10625 34563 10659
rect 34563 10625 34572 10659
rect 34520 10616 34572 10625
rect 36176 10684 36228 10736
rect 36912 10727 36964 10736
rect 34796 10616 34848 10668
rect 36544 10616 36596 10668
rect 36912 10693 36939 10727
rect 36939 10693 36964 10727
rect 36912 10684 36964 10693
rect 37004 10616 37056 10668
rect 37188 10616 37240 10668
rect 36176 10591 36228 10600
rect 36176 10557 36185 10591
rect 36185 10557 36219 10591
rect 36219 10557 36228 10591
rect 36176 10548 36228 10557
rect 8576 10412 8628 10464
rect 8668 10412 8720 10464
rect 11336 10412 11388 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 17868 10412 17920 10464
rect 18512 10412 18564 10464
rect 21456 10455 21508 10464
rect 21456 10421 21465 10455
rect 21465 10421 21499 10455
rect 21499 10421 21508 10455
rect 21456 10412 21508 10421
rect 21824 10455 21876 10464
rect 21824 10421 21833 10455
rect 21833 10421 21867 10455
rect 21867 10421 21876 10455
rect 21824 10412 21876 10421
rect 22376 10412 22428 10464
rect 24032 10480 24084 10532
rect 26148 10480 26200 10532
rect 27896 10480 27948 10532
rect 36084 10480 36136 10532
rect 36912 10548 36964 10600
rect 38384 10591 38436 10600
rect 38384 10557 38393 10591
rect 38393 10557 38427 10591
rect 38427 10557 38436 10591
rect 38384 10548 38436 10557
rect 24676 10412 24728 10464
rect 28264 10412 28316 10464
rect 30748 10412 30800 10464
rect 32312 10412 32364 10464
rect 32772 10455 32824 10464
rect 32772 10421 32781 10455
rect 32781 10421 32815 10455
rect 32815 10421 32824 10455
rect 32772 10412 32824 10421
rect 32956 10412 33008 10464
rect 33232 10412 33284 10464
rect 34612 10412 34664 10464
rect 35348 10412 35400 10464
rect 37832 10480 37884 10532
rect 36820 10412 36872 10464
rect 37280 10455 37332 10464
rect 37280 10421 37289 10455
rect 37289 10421 37323 10455
rect 37323 10421 37332 10455
rect 37280 10412 37332 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1308 10208 1360 10260
rect 8392 10208 8444 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 13820 10208 13872 10260
rect 14464 10208 14516 10260
rect 17960 10208 18012 10260
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 20720 10251 20772 10260
rect 20720 10217 20729 10251
rect 20729 10217 20763 10251
rect 20763 10217 20772 10251
rect 20720 10208 20772 10217
rect 23388 10208 23440 10260
rect 23664 10251 23716 10260
rect 23664 10217 23673 10251
rect 23673 10217 23707 10251
rect 23707 10217 23716 10251
rect 23664 10208 23716 10217
rect 14924 10140 14976 10192
rect 17132 10140 17184 10192
rect 4804 10072 4856 10124
rect 6552 10072 6604 10124
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 8576 10072 8628 10124
rect 11060 10072 11112 10124
rect 11612 10072 11664 10124
rect 12624 10072 12676 10124
rect 13176 10072 13228 10124
rect 15384 10072 15436 10124
rect 5264 9979 5316 9988
rect 5264 9945 5273 9979
rect 5273 9945 5307 9979
rect 5307 9945 5316 9979
rect 5264 9936 5316 9945
rect 940 9868 992 9920
rect 3884 9868 3936 9920
rect 8300 10004 8352 10056
rect 10324 10004 10376 10056
rect 10876 10004 10928 10056
rect 12900 10004 12952 10056
rect 13452 10004 13504 10056
rect 14188 10004 14240 10056
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 14648 10004 14700 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 11888 9936 11940 9988
rect 14004 9936 14056 9988
rect 16488 10047 16540 10056
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 17224 10072 17276 10124
rect 17776 10072 17828 10124
rect 18696 10115 18748 10124
rect 18696 10081 18705 10115
rect 18705 10081 18739 10115
rect 18739 10081 18748 10115
rect 18696 10072 18748 10081
rect 21824 10140 21876 10192
rect 21916 10140 21968 10192
rect 23940 10208 23992 10260
rect 24032 10251 24084 10260
rect 24032 10217 24041 10251
rect 24041 10217 24075 10251
rect 24075 10217 24084 10251
rect 24032 10208 24084 10217
rect 27160 10208 27212 10260
rect 28540 10208 28592 10260
rect 29000 10208 29052 10260
rect 30104 10251 30156 10260
rect 30104 10217 30113 10251
rect 30113 10217 30147 10251
rect 30147 10217 30156 10251
rect 30104 10208 30156 10217
rect 31024 10208 31076 10260
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 21456 10004 21508 10056
rect 6736 9911 6788 9920
rect 6736 9877 6745 9911
rect 6745 9877 6779 9911
rect 6779 9877 6788 9911
rect 6736 9868 6788 9877
rect 6828 9911 6880 9920
rect 6828 9877 6837 9911
rect 6837 9877 6871 9911
rect 6871 9877 6880 9911
rect 6828 9868 6880 9877
rect 9680 9868 9732 9920
rect 11244 9911 11296 9920
rect 11244 9877 11253 9911
rect 11253 9877 11287 9911
rect 11287 9877 11296 9911
rect 11244 9868 11296 9877
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 13176 9911 13228 9920
rect 13176 9877 13185 9911
rect 13185 9877 13219 9911
rect 13219 9877 13228 9911
rect 13176 9868 13228 9877
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 13544 9868 13596 9877
rect 16672 9868 16724 9920
rect 16856 9868 16908 9920
rect 17316 9868 17368 9920
rect 18328 9936 18380 9988
rect 19248 9936 19300 9988
rect 23112 10115 23164 10124
rect 23112 10081 23121 10115
rect 23121 10081 23155 10115
rect 23155 10081 23164 10115
rect 23112 10072 23164 10081
rect 27804 10140 27856 10192
rect 29092 10140 29144 10192
rect 23204 10004 23256 10056
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 24676 10115 24728 10124
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 24768 10115 24820 10124
rect 24768 10081 24777 10115
rect 24777 10081 24811 10115
rect 24811 10081 24820 10115
rect 24768 10072 24820 10081
rect 25688 10115 25740 10124
rect 25688 10081 25697 10115
rect 25697 10081 25731 10115
rect 25731 10081 25740 10115
rect 25688 10072 25740 10081
rect 26148 10115 26200 10124
rect 26148 10081 26157 10115
rect 26157 10081 26191 10115
rect 26191 10081 26200 10115
rect 26148 10072 26200 10081
rect 29644 10115 29696 10124
rect 29644 10081 29653 10115
rect 29653 10081 29687 10115
rect 29687 10081 29696 10115
rect 29644 10072 29696 10081
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 23848 10013 23851 10022
rect 23851 10013 23885 10022
rect 23885 10013 23900 10022
rect 23848 9970 23900 10013
rect 24124 10047 24176 10056
rect 24124 10013 24133 10047
rect 24133 10013 24167 10047
rect 24167 10013 24176 10047
rect 24124 10004 24176 10013
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 24492 10004 24544 10056
rect 25136 10004 25188 10056
rect 21548 9911 21600 9920
rect 21548 9877 21557 9911
rect 21557 9877 21591 9911
rect 21591 9877 21600 9911
rect 21548 9868 21600 9877
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 22192 9868 22244 9920
rect 22928 9868 22980 9920
rect 25780 9936 25832 9988
rect 25964 10004 26016 10056
rect 28264 10047 28316 10056
rect 28264 10013 28273 10047
rect 28273 10013 28307 10047
rect 28307 10013 28316 10047
rect 28264 10004 28316 10013
rect 27436 9936 27488 9988
rect 28448 9979 28500 9988
rect 28448 9945 28457 9979
rect 28457 9945 28491 9979
rect 28491 9945 28500 9979
rect 29736 10047 29788 10056
rect 29736 10013 29745 10047
rect 29745 10013 29779 10047
rect 29779 10013 29788 10047
rect 29736 10004 29788 10013
rect 30288 10140 30340 10192
rect 30748 10047 30800 10056
rect 30748 10013 30757 10047
rect 30757 10013 30791 10047
rect 30791 10013 30800 10047
rect 30748 10004 30800 10013
rect 28448 9936 28500 9945
rect 32404 10140 32456 10192
rect 34520 10208 34572 10260
rect 34980 10208 35032 10260
rect 34612 10140 34664 10192
rect 31116 10115 31168 10124
rect 31116 10081 31125 10115
rect 31125 10081 31159 10115
rect 31159 10081 31168 10115
rect 31116 10072 31168 10081
rect 31576 10047 31628 10056
rect 31576 10013 31585 10047
rect 31585 10013 31619 10047
rect 31619 10013 31628 10047
rect 31576 10004 31628 10013
rect 37280 10072 37332 10124
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 30932 9868 30984 9920
rect 31484 9979 31536 9988
rect 31484 9945 31493 9979
rect 31493 9945 31527 9979
rect 31527 9945 31536 9979
rect 34612 10004 34664 10056
rect 36636 10047 36688 10056
rect 36636 10013 36645 10047
rect 36645 10013 36679 10047
rect 36679 10013 36688 10047
rect 36636 10004 36688 10013
rect 31484 9936 31536 9945
rect 31668 9868 31720 9920
rect 32128 9868 32180 9920
rect 34336 9911 34388 9920
rect 34336 9877 34345 9911
rect 34345 9877 34379 9911
rect 34379 9877 34388 9911
rect 34336 9868 34388 9877
rect 35440 9936 35492 9988
rect 37372 9936 37424 9988
rect 36820 9868 36872 9920
rect 38384 9911 38436 9920
rect 38384 9877 38393 9911
rect 38393 9877 38427 9911
rect 38427 9877 38436 9911
rect 38384 9868 38436 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 10968 9664 11020 9716
rect 11888 9664 11940 9716
rect 13360 9664 13412 9716
rect 13544 9664 13596 9716
rect 9864 9596 9916 9648
rect 11244 9639 11296 9648
rect 11244 9605 11253 9639
rect 11253 9605 11287 9639
rect 11287 9605 11296 9639
rect 11244 9596 11296 9605
rect 13084 9596 13136 9648
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 16488 9664 16540 9716
rect 17316 9664 17368 9716
rect 18236 9664 18288 9716
rect 23020 9664 23072 9716
rect 23480 9664 23532 9716
rect 23664 9664 23716 9716
rect 24400 9664 24452 9716
rect 14280 9596 14332 9648
rect 14648 9596 14700 9648
rect 6828 9528 6880 9580
rect 7196 9528 7248 9580
rect 8484 9528 8536 9580
rect 10692 9528 10744 9580
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 8116 9460 8168 9512
rect 6644 9324 6696 9376
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 12624 9503 12676 9512
rect 12624 9469 12633 9503
rect 12633 9469 12667 9503
rect 12667 9469 12676 9503
rect 12624 9460 12676 9469
rect 11060 9392 11112 9444
rect 15660 9528 15712 9580
rect 16672 9596 16724 9648
rect 20996 9596 21048 9648
rect 21916 9596 21968 9648
rect 22192 9639 22244 9648
rect 22192 9605 22201 9639
rect 22201 9605 22235 9639
rect 22235 9605 22244 9639
rect 22192 9596 22244 9605
rect 14004 9460 14056 9512
rect 14188 9460 14240 9512
rect 14924 9460 14976 9512
rect 16396 9571 16448 9580
rect 16396 9537 16405 9571
rect 16405 9537 16439 9571
rect 16439 9537 16448 9571
rect 16396 9528 16448 9537
rect 16488 9528 16540 9580
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 22376 9571 22428 9580
rect 22376 9537 22385 9571
rect 22385 9537 22419 9571
rect 22419 9537 22428 9571
rect 22376 9528 22428 9537
rect 16948 9460 17000 9512
rect 17960 9460 18012 9512
rect 14280 9392 14332 9444
rect 15200 9435 15252 9444
rect 15200 9401 15209 9435
rect 15209 9401 15243 9435
rect 15243 9401 15252 9435
rect 15200 9392 15252 9401
rect 16396 9392 16448 9444
rect 10508 9324 10560 9376
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 12808 9324 12860 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 15292 9324 15344 9376
rect 17592 9324 17644 9376
rect 19708 9460 19760 9512
rect 21548 9460 21600 9512
rect 19248 9392 19300 9444
rect 22928 9528 22980 9580
rect 23204 9571 23256 9580
rect 23204 9537 23213 9571
rect 23213 9537 23247 9571
rect 23247 9537 23256 9571
rect 23204 9528 23256 9537
rect 23940 9596 23992 9648
rect 24860 9596 24912 9648
rect 25964 9664 26016 9716
rect 28448 9664 28500 9716
rect 29644 9664 29696 9716
rect 31484 9664 31536 9716
rect 31668 9707 31720 9716
rect 31668 9673 31677 9707
rect 31677 9673 31711 9707
rect 31711 9673 31720 9707
rect 31668 9664 31720 9673
rect 34336 9664 34388 9716
rect 34612 9664 34664 9716
rect 36912 9664 36964 9716
rect 23664 9571 23716 9580
rect 23664 9537 23673 9571
rect 23673 9537 23707 9571
rect 23707 9537 23716 9571
rect 23664 9528 23716 9537
rect 24952 9528 25004 9580
rect 25688 9639 25740 9648
rect 25688 9605 25697 9639
rect 25697 9605 25731 9639
rect 25731 9605 25740 9639
rect 25688 9596 25740 9605
rect 27804 9596 27856 9648
rect 25780 9528 25832 9580
rect 23020 9503 23072 9512
rect 23020 9469 23029 9503
rect 23029 9469 23063 9503
rect 23063 9469 23072 9503
rect 23020 9460 23072 9469
rect 26056 9460 26108 9512
rect 26240 9528 26292 9580
rect 28172 9528 28224 9580
rect 28356 9528 28408 9580
rect 29092 9528 29144 9580
rect 31024 9596 31076 9648
rect 29736 9571 29788 9580
rect 29736 9537 29745 9571
rect 29745 9537 29779 9571
rect 29779 9537 29788 9571
rect 29736 9528 29788 9537
rect 32128 9571 32180 9580
rect 32128 9537 32137 9571
rect 32137 9537 32171 9571
rect 32171 9537 32180 9571
rect 32128 9528 32180 9537
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 32404 9571 32456 9580
rect 32404 9537 32413 9571
rect 32413 9537 32447 9571
rect 32447 9537 32456 9571
rect 32404 9528 32456 9537
rect 32680 9571 32732 9580
rect 32680 9537 32689 9571
rect 32689 9537 32723 9571
rect 32723 9537 32732 9571
rect 32680 9528 32732 9537
rect 32772 9528 32824 9580
rect 24032 9392 24084 9444
rect 31024 9503 31076 9512
rect 31024 9469 31033 9503
rect 31033 9469 31067 9503
rect 31067 9469 31076 9503
rect 31024 9460 31076 9469
rect 34980 9528 35032 9580
rect 35440 9639 35492 9648
rect 35440 9605 35449 9639
rect 35449 9605 35483 9639
rect 35483 9605 35492 9639
rect 35440 9596 35492 9605
rect 35532 9571 35584 9580
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 32680 9392 32732 9444
rect 34428 9460 34480 9512
rect 34612 9503 34664 9512
rect 34612 9469 34621 9503
rect 34621 9469 34655 9503
rect 34655 9469 34664 9503
rect 34612 9460 34664 9469
rect 22928 9324 22980 9376
rect 24584 9324 24636 9376
rect 26424 9324 26476 9376
rect 29092 9324 29144 9376
rect 30932 9367 30984 9376
rect 30932 9333 30941 9367
rect 30941 9333 30975 9367
rect 30975 9333 30984 9367
rect 30932 9324 30984 9333
rect 33416 9367 33468 9376
rect 33416 9333 33425 9367
rect 33425 9333 33459 9367
rect 33459 9333 33468 9367
rect 33416 9324 33468 9333
rect 34704 9324 34756 9376
rect 35440 9460 35492 9512
rect 35624 9503 35676 9512
rect 35624 9469 35633 9503
rect 35633 9469 35667 9503
rect 35667 9469 35676 9503
rect 35624 9460 35676 9469
rect 35808 9503 35860 9512
rect 35808 9469 35817 9503
rect 35817 9469 35851 9503
rect 35851 9469 35860 9503
rect 35808 9460 35860 9469
rect 36544 9571 36596 9580
rect 36544 9537 36553 9571
rect 36553 9537 36587 9571
rect 36587 9537 36596 9571
rect 36544 9528 36596 9537
rect 36820 9571 36872 9580
rect 36820 9537 36829 9571
rect 36829 9537 36863 9571
rect 36863 9537 36872 9571
rect 36820 9528 36872 9537
rect 36912 9571 36964 9580
rect 36912 9537 36921 9571
rect 36921 9537 36955 9571
rect 36955 9537 36964 9571
rect 36912 9528 36964 9537
rect 37188 9596 37240 9648
rect 37280 9528 37332 9580
rect 36728 9503 36780 9512
rect 36728 9469 36737 9503
rect 36737 9469 36771 9503
rect 36771 9469 36780 9503
rect 36728 9460 36780 9469
rect 34980 9392 35032 9444
rect 34888 9324 34940 9376
rect 35900 9324 35952 9376
rect 36176 9392 36228 9444
rect 37004 9392 37056 9444
rect 37464 9460 37516 9512
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 8116 9163 8168 9172
rect 8116 9129 8125 9163
rect 8125 9129 8159 9163
rect 8159 9129 8168 9163
rect 8116 9120 8168 9129
rect 9404 9120 9456 9172
rect 10968 9120 11020 9172
rect 14556 9120 14608 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 16764 9163 16816 9172
rect 16764 9129 16773 9163
rect 16773 9129 16807 9163
rect 16807 9129 16816 9163
rect 16764 9120 16816 9129
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 26148 9120 26200 9172
rect 28172 9163 28224 9172
rect 28172 9129 28181 9163
rect 28181 9129 28215 9163
rect 28215 9129 28224 9163
rect 28172 9120 28224 9129
rect 28356 9163 28408 9172
rect 28356 9129 28365 9163
rect 28365 9129 28399 9163
rect 28399 9129 28408 9163
rect 28356 9120 28408 9129
rect 15384 9052 15436 9104
rect 21732 9052 21784 9104
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 13176 8984 13228 9036
rect 5448 8848 5500 8900
rect 9496 8916 9548 8968
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 9956 8959 10008 8968
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 10508 8916 10560 8968
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 14004 8984 14056 9036
rect 14188 8916 14240 8968
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 15844 8916 15896 8968
rect 18696 8984 18748 9036
rect 6552 8848 6604 8900
rect 8300 8891 8352 8900
rect 8300 8857 8309 8891
rect 8309 8857 8343 8891
rect 8343 8857 8352 8891
rect 8300 8848 8352 8857
rect 8576 8848 8628 8900
rect 7012 8780 7064 8832
rect 10876 8848 10928 8900
rect 13452 8848 13504 8900
rect 15016 8891 15068 8900
rect 15016 8857 15025 8891
rect 15025 8857 15059 8891
rect 15059 8857 15068 8891
rect 15016 8848 15068 8857
rect 18328 8959 18380 8968
rect 18328 8925 18337 8959
rect 18337 8925 18371 8959
rect 18371 8925 18380 8959
rect 18328 8916 18380 8925
rect 23204 8916 23256 8968
rect 25780 9052 25832 9104
rect 26056 8984 26108 9036
rect 25228 8959 25280 8968
rect 25228 8925 25237 8959
rect 25237 8925 25271 8959
rect 25271 8925 25280 8959
rect 25228 8916 25280 8925
rect 21640 8891 21692 8900
rect 21640 8857 21649 8891
rect 21649 8857 21683 8891
rect 21683 8857 21692 8891
rect 26332 8916 26384 8968
rect 31024 9120 31076 9172
rect 32680 9120 32732 9172
rect 35348 9120 35400 9172
rect 35808 9120 35860 9172
rect 36176 9120 36228 9172
rect 36728 9120 36780 9172
rect 33968 9052 34020 9104
rect 31300 8984 31352 9036
rect 34520 8984 34572 9036
rect 36636 9027 36688 9036
rect 36636 8993 36645 9027
rect 36645 8993 36679 9027
rect 36679 8993 36688 9027
rect 36636 8984 36688 8993
rect 21640 8848 21692 8857
rect 25596 8848 25648 8900
rect 10692 8780 10744 8832
rect 15108 8780 15160 8832
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 15660 8780 15712 8832
rect 16488 8780 16540 8832
rect 18696 8780 18748 8832
rect 21824 8823 21876 8832
rect 21824 8789 21833 8823
rect 21833 8789 21867 8823
rect 21867 8789 21876 8823
rect 21824 8780 21876 8789
rect 25412 8780 25464 8832
rect 25504 8823 25556 8832
rect 25504 8789 25513 8823
rect 25513 8789 25547 8823
rect 25547 8789 25556 8823
rect 25504 8780 25556 8789
rect 25964 8848 26016 8900
rect 27988 8891 28040 8900
rect 27988 8857 27997 8891
rect 27997 8857 28031 8891
rect 28031 8857 28040 8891
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 30104 8959 30156 8968
rect 30104 8925 30113 8959
rect 30113 8925 30147 8959
rect 30147 8925 30156 8959
rect 30104 8916 30156 8925
rect 27988 8848 28040 8857
rect 31760 8916 31812 8968
rect 31852 8959 31904 8968
rect 31852 8925 31861 8959
rect 31861 8925 31895 8959
rect 31895 8925 31904 8959
rect 31852 8916 31904 8925
rect 34704 8916 34756 8968
rect 34336 8848 34388 8900
rect 35532 8916 35584 8968
rect 36452 8959 36504 8968
rect 36452 8925 36461 8959
rect 36461 8925 36495 8959
rect 36495 8925 36504 8959
rect 36452 8916 36504 8925
rect 36912 8891 36964 8900
rect 36912 8857 36921 8891
rect 36921 8857 36955 8891
rect 36955 8857 36964 8891
rect 36912 8848 36964 8857
rect 37372 8848 37424 8900
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 36176 8780 36228 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 5356 8576 5408 8628
rect 3884 8440 3936 8492
rect 4804 8508 4856 8560
rect 4712 8440 4764 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 6828 8508 6880 8560
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 8300 8508 8352 8560
rect 9496 8508 9548 8560
rect 8576 8372 8628 8424
rect 11612 8576 11664 8628
rect 9772 8508 9824 8560
rect 14464 8576 14516 8628
rect 15568 8576 15620 8628
rect 17316 8576 17368 8628
rect 18696 8576 18748 8628
rect 22284 8576 22336 8628
rect 12808 8551 12860 8560
rect 12808 8517 12817 8551
rect 12817 8517 12851 8551
rect 12851 8517 12860 8551
rect 12808 8508 12860 8517
rect 13452 8508 13504 8560
rect 15108 8508 15160 8560
rect 16396 8508 16448 8560
rect 20996 8508 21048 8560
rect 21824 8508 21876 8560
rect 7472 8304 7524 8356
rect 2872 8236 2924 8288
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 5356 8236 5408 8245
rect 6000 8236 6052 8288
rect 6736 8236 6788 8288
rect 7748 8236 7800 8288
rect 9128 8236 9180 8288
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 9864 8372 9916 8381
rect 11704 8372 11756 8424
rect 14280 8415 14332 8424
rect 14280 8381 14289 8415
rect 14289 8381 14323 8415
rect 14323 8381 14332 8415
rect 14280 8372 14332 8381
rect 16212 8415 16264 8424
rect 16212 8381 16221 8415
rect 16221 8381 16255 8415
rect 16255 8381 16264 8415
rect 16212 8372 16264 8381
rect 17776 8415 17828 8424
rect 17776 8381 17785 8415
rect 17785 8381 17819 8415
rect 17819 8381 17828 8415
rect 17776 8372 17828 8381
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 23204 8440 23256 8492
rect 18604 8372 18656 8424
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 21456 8372 21508 8424
rect 23480 8483 23532 8492
rect 23480 8449 23489 8483
rect 23489 8449 23523 8483
rect 23523 8449 23532 8483
rect 23480 8440 23532 8449
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 24860 8576 24912 8628
rect 25228 8576 25280 8628
rect 26332 8576 26384 8628
rect 27988 8576 28040 8628
rect 29736 8576 29788 8628
rect 31300 8619 31352 8628
rect 31300 8585 31309 8619
rect 31309 8585 31343 8619
rect 31343 8585 31352 8619
rect 31300 8576 31352 8585
rect 31668 8619 31720 8628
rect 31668 8585 31693 8619
rect 31693 8585 31720 8619
rect 31668 8576 31720 8585
rect 31852 8619 31904 8628
rect 31852 8585 31861 8619
rect 31861 8585 31895 8619
rect 31895 8585 31904 8619
rect 31852 8576 31904 8585
rect 35256 8619 35308 8628
rect 35256 8585 35265 8619
rect 35265 8585 35299 8619
rect 35299 8585 35308 8619
rect 35256 8576 35308 8585
rect 36912 8576 36964 8628
rect 25596 8508 25648 8560
rect 24584 8440 24636 8492
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25504 8483 25556 8492
rect 25504 8449 25513 8483
rect 25513 8449 25547 8483
rect 25547 8449 25556 8483
rect 27436 8508 27488 8560
rect 28632 8508 28684 8560
rect 25504 8440 25556 8449
rect 26240 8440 26292 8492
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 28080 8483 28132 8492
rect 28080 8449 28089 8483
rect 28089 8449 28123 8483
rect 28123 8449 28132 8483
rect 28080 8440 28132 8449
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 31116 8483 31168 8492
rect 31116 8449 31125 8483
rect 31125 8449 31159 8483
rect 31159 8449 31168 8483
rect 31116 8440 31168 8449
rect 33968 8508 34020 8560
rect 34336 8483 34388 8492
rect 34336 8449 34345 8483
rect 34345 8449 34379 8483
rect 34379 8449 34388 8483
rect 34336 8440 34388 8449
rect 35992 8440 36044 8492
rect 37280 8440 37332 8492
rect 22376 8304 22428 8356
rect 27068 8415 27120 8424
rect 27068 8381 27077 8415
rect 27077 8381 27111 8415
rect 27111 8381 27120 8415
rect 27068 8372 27120 8381
rect 34612 8415 34664 8424
rect 34612 8381 34621 8415
rect 34621 8381 34655 8415
rect 34655 8381 34664 8415
rect 34612 8372 34664 8381
rect 34796 8415 34848 8424
rect 34796 8381 34805 8415
rect 34805 8381 34839 8415
rect 34839 8381 34848 8415
rect 34796 8372 34848 8381
rect 10508 8236 10560 8288
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 14372 8236 14424 8288
rect 15660 8279 15712 8288
rect 15660 8245 15669 8279
rect 15669 8245 15703 8279
rect 15703 8245 15712 8279
rect 15660 8236 15712 8245
rect 17224 8236 17276 8288
rect 24308 8279 24360 8288
rect 24308 8245 24317 8279
rect 24317 8245 24351 8279
rect 24351 8245 24360 8279
rect 24308 8236 24360 8245
rect 24860 8304 24912 8356
rect 31760 8304 31812 8356
rect 24952 8236 25004 8288
rect 26608 8236 26660 8288
rect 31300 8236 31352 8288
rect 34428 8279 34480 8288
rect 34428 8245 34437 8279
rect 34437 8245 34471 8279
rect 34471 8245 34480 8279
rect 34428 8236 34480 8245
rect 34796 8236 34848 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 6828 8075 6880 8084
rect 6828 8041 6837 8075
rect 6837 8041 6871 8075
rect 6871 8041 6880 8075
rect 6828 8032 6880 8041
rect 7196 8032 7248 8084
rect 7472 8032 7524 8084
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 9864 8032 9916 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 18696 8075 18748 8084
rect 18696 8041 18705 8075
rect 18705 8041 18739 8075
rect 18739 8041 18748 8075
rect 18696 8032 18748 8041
rect 23020 8032 23072 8084
rect 23296 8032 23348 8084
rect 9588 7964 9640 8016
rect 21180 7964 21232 8016
rect 21364 7964 21416 8016
rect 5448 7896 5500 7948
rect 8116 7896 8168 7948
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 6828 7828 6880 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 3424 7760 3476 7812
rect 3976 7760 4028 7812
rect 4804 7692 4856 7744
rect 5356 7803 5408 7812
rect 5356 7769 5365 7803
rect 5365 7769 5399 7803
rect 5399 7769 5408 7803
rect 5356 7760 5408 7769
rect 8852 7760 8904 7812
rect 7012 7692 7064 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 11520 7896 11572 7948
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 14372 7939 14424 7948
rect 14372 7905 14381 7939
rect 14381 7905 14415 7939
rect 14415 7905 14424 7939
rect 14372 7896 14424 7905
rect 16212 7939 16264 7948
rect 16212 7905 16221 7939
rect 16221 7905 16255 7939
rect 16255 7905 16264 7939
rect 16212 7896 16264 7905
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 17224 7939 17276 7948
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 16672 7828 16724 7880
rect 21364 7871 21416 7880
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 22468 7871 22520 7880
rect 22468 7837 22477 7871
rect 22477 7837 22511 7871
rect 22511 7837 22520 7871
rect 22468 7828 22520 7837
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 23296 7871 23348 7880
rect 23296 7837 23305 7871
rect 23305 7837 23339 7871
rect 23339 7837 23348 7871
rect 24676 7964 24728 8016
rect 24216 7896 24268 7948
rect 23296 7828 23348 7837
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 24308 7828 24360 7880
rect 24952 7964 25004 8016
rect 25228 7964 25280 8016
rect 27068 8032 27120 8084
rect 31116 8075 31168 8084
rect 31116 8041 31125 8075
rect 31125 8041 31159 8075
rect 31159 8041 31168 8075
rect 31116 8032 31168 8041
rect 28264 7964 28316 8016
rect 30104 8007 30156 8016
rect 30104 7973 30113 8007
rect 30113 7973 30147 8007
rect 30147 7973 30156 8007
rect 30104 7964 30156 7973
rect 34704 8032 34756 8084
rect 10324 7760 10376 7812
rect 11336 7760 11388 7812
rect 15384 7760 15436 7812
rect 18236 7760 18288 7812
rect 21824 7760 21876 7812
rect 22008 7760 22060 7812
rect 23664 7760 23716 7812
rect 24216 7760 24268 7812
rect 24860 7871 24912 7880
rect 24860 7837 24874 7871
rect 24874 7837 24908 7871
rect 24908 7837 24912 7871
rect 24860 7828 24912 7837
rect 25320 7871 25372 7880
rect 25320 7837 25329 7871
rect 25329 7837 25363 7871
rect 25363 7837 25372 7871
rect 25320 7828 25372 7837
rect 26792 7871 26844 7880
rect 26792 7837 26801 7871
rect 26801 7837 26835 7871
rect 26835 7837 26844 7871
rect 26792 7828 26844 7837
rect 24952 7760 25004 7812
rect 27344 7871 27396 7880
rect 27344 7837 27353 7871
rect 27353 7837 27387 7871
rect 27387 7837 27396 7871
rect 27344 7828 27396 7837
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 28632 7828 28684 7880
rect 33784 7896 33836 7948
rect 27160 7760 27212 7812
rect 29184 7760 29236 7812
rect 31392 7828 31444 7880
rect 31760 7871 31812 7880
rect 31760 7837 31769 7871
rect 31769 7837 31803 7871
rect 31803 7837 31812 7871
rect 31760 7828 31812 7837
rect 36544 7964 36596 8016
rect 36820 7964 36872 8016
rect 34428 7896 34480 7948
rect 34796 7828 34848 7880
rect 35256 7828 35308 7880
rect 30380 7803 30432 7812
rect 30380 7769 30389 7803
rect 30389 7769 30423 7803
rect 30423 7769 30432 7803
rect 30380 7760 30432 7769
rect 36268 7828 36320 7880
rect 37280 8032 37332 8084
rect 37004 7760 37056 7812
rect 37280 7871 37332 7880
rect 37280 7837 37289 7871
rect 37289 7837 37323 7871
rect 37323 7837 37332 7871
rect 37280 7828 37332 7837
rect 38476 7896 38528 7948
rect 37924 7871 37976 7880
rect 37924 7837 37933 7871
rect 37933 7837 37967 7871
rect 37967 7837 37976 7871
rect 37924 7828 37976 7837
rect 7288 7692 7340 7701
rect 11520 7692 11572 7744
rect 16488 7735 16540 7744
rect 16488 7701 16497 7735
rect 16497 7701 16531 7735
rect 16531 7701 16540 7735
rect 16488 7692 16540 7701
rect 16948 7692 17000 7744
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22100 7692 22152 7701
rect 22376 7692 22428 7744
rect 23296 7692 23348 7744
rect 24584 7692 24636 7744
rect 31944 7735 31996 7744
rect 31944 7701 31953 7735
rect 31953 7701 31987 7735
rect 31987 7701 31996 7735
rect 31944 7692 31996 7701
rect 33508 7692 33560 7744
rect 35348 7735 35400 7744
rect 35348 7701 35357 7735
rect 35357 7701 35391 7735
rect 35391 7701 35400 7735
rect 35348 7692 35400 7701
rect 35992 7692 36044 7744
rect 36084 7692 36136 7744
rect 37372 7735 37424 7744
rect 37372 7701 37381 7735
rect 37381 7701 37415 7735
rect 37415 7701 37424 7735
rect 37372 7692 37424 7701
rect 38384 7735 38436 7744
rect 38384 7701 38393 7735
rect 38393 7701 38427 7735
rect 38427 7701 38436 7735
rect 38384 7692 38436 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 10324 7531 10376 7540
rect 10324 7497 10333 7531
rect 10333 7497 10367 7531
rect 10367 7497 10376 7531
rect 10324 7488 10376 7497
rect 11152 7488 11204 7540
rect 2872 7463 2924 7472
rect 2872 7429 2881 7463
rect 2881 7429 2915 7463
rect 2915 7429 2924 7463
rect 2872 7420 2924 7429
rect 3976 7352 4028 7404
rect 848 7284 900 7336
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 4068 7284 4120 7336
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5264 7352 5316 7404
rect 7564 7352 7616 7404
rect 10140 7463 10192 7472
rect 10140 7429 10165 7463
rect 10165 7429 10192 7463
rect 10140 7420 10192 7429
rect 10416 7463 10468 7472
rect 10416 7429 10425 7463
rect 10425 7429 10459 7463
rect 10459 7429 10468 7463
rect 10416 7420 10468 7429
rect 15660 7488 15712 7540
rect 16396 7488 16448 7540
rect 16488 7488 16540 7540
rect 17776 7488 17828 7540
rect 21364 7488 21416 7540
rect 22744 7488 22796 7540
rect 15200 7420 15252 7472
rect 16948 7463 17000 7472
rect 16948 7429 16957 7463
rect 16957 7429 16991 7463
rect 16991 7429 17000 7463
rect 16948 7420 17000 7429
rect 18236 7420 18288 7472
rect 19984 7420 20036 7472
rect 11336 7352 11388 7404
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 22100 7352 22152 7404
rect 24216 7488 24268 7540
rect 22928 7395 22980 7404
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 23296 7420 23348 7472
rect 25044 7488 25096 7540
rect 25136 7488 25188 7540
rect 26792 7488 26844 7540
rect 27344 7488 27396 7540
rect 37924 7488 37976 7540
rect 8576 7284 8628 7336
rect 10508 7284 10560 7336
rect 11060 7284 11112 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 21456 7284 21508 7336
rect 21640 7284 21692 7336
rect 21732 7216 21784 7268
rect 23296 7216 23348 7268
rect 4436 7148 4488 7200
rect 4804 7148 4856 7200
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 7748 7148 7800 7200
rect 10784 7148 10836 7200
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 23848 7191 23900 7200
rect 23848 7157 23857 7191
rect 23857 7157 23891 7191
rect 23891 7157 23900 7191
rect 23848 7148 23900 7157
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 24768 7395 24820 7404
rect 24768 7361 24778 7395
rect 24778 7361 24812 7395
rect 24812 7361 24820 7395
rect 24768 7352 24820 7361
rect 24952 7395 25004 7404
rect 24952 7361 24961 7395
rect 24961 7361 24995 7395
rect 24995 7361 25004 7395
rect 24952 7352 25004 7361
rect 25044 7395 25096 7404
rect 25044 7361 25053 7395
rect 25053 7361 25087 7395
rect 25087 7361 25096 7395
rect 25044 7352 25096 7361
rect 25136 7395 25188 7404
rect 25136 7361 25150 7395
rect 25150 7361 25184 7395
rect 25184 7361 25188 7395
rect 25136 7352 25188 7361
rect 27528 7352 27580 7404
rect 32312 7395 32364 7404
rect 32312 7361 32321 7395
rect 32321 7361 32355 7395
rect 32355 7361 32364 7395
rect 32312 7352 32364 7361
rect 31944 7284 31996 7336
rect 32956 7395 33008 7404
rect 32956 7361 32965 7395
rect 32965 7361 32999 7395
rect 32999 7361 33008 7395
rect 32956 7352 33008 7361
rect 33140 7395 33192 7404
rect 33140 7361 33149 7395
rect 33149 7361 33183 7395
rect 33183 7361 33192 7395
rect 33140 7352 33192 7361
rect 33416 7395 33468 7404
rect 33416 7361 33425 7395
rect 33425 7361 33459 7395
rect 33459 7361 33468 7395
rect 33416 7352 33468 7361
rect 33508 7395 33560 7404
rect 33508 7361 33517 7395
rect 33517 7361 33551 7395
rect 33551 7361 33560 7395
rect 33508 7352 33560 7361
rect 33692 7395 33744 7404
rect 33692 7361 33701 7395
rect 33701 7361 33735 7395
rect 33735 7361 33744 7395
rect 33692 7352 33744 7361
rect 36084 7352 36136 7404
rect 36176 7395 36228 7404
rect 36176 7361 36185 7395
rect 36185 7361 36219 7395
rect 36219 7361 36228 7395
rect 36176 7352 36228 7361
rect 37004 7420 37056 7472
rect 36452 7395 36504 7404
rect 36452 7361 36461 7395
rect 36461 7361 36495 7395
rect 36495 7361 36504 7395
rect 36452 7352 36504 7361
rect 36544 7395 36596 7404
rect 36544 7361 36553 7395
rect 36553 7361 36587 7395
rect 36587 7361 36596 7395
rect 36544 7352 36596 7361
rect 35808 7327 35860 7336
rect 35808 7293 35817 7327
rect 35817 7293 35851 7327
rect 35851 7293 35860 7327
rect 35808 7284 35860 7293
rect 24676 7216 24728 7268
rect 27436 7216 27488 7268
rect 32680 7259 32732 7268
rect 32680 7225 32689 7259
rect 32689 7225 32723 7259
rect 32723 7225 32732 7259
rect 32680 7216 32732 7225
rect 24952 7148 25004 7200
rect 25504 7148 25556 7200
rect 33416 7148 33468 7200
rect 35716 7148 35768 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3976 6987 4028 6996
rect 3976 6953 3985 6987
rect 3985 6953 4019 6987
rect 4019 6953 4028 6987
rect 3976 6944 4028 6953
rect 4896 6944 4948 6996
rect 7196 6944 7248 6996
rect 20720 6944 20772 6996
rect 21456 6987 21508 6996
rect 21456 6953 21465 6987
rect 21465 6953 21499 6987
rect 21499 6953 21508 6987
rect 21456 6944 21508 6953
rect 27804 6987 27856 6996
rect 27804 6953 27813 6987
rect 27813 6953 27847 6987
rect 27847 6953 27856 6987
rect 27804 6944 27856 6953
rect 30380 6987 30432 6996
rect 30380 6953 30389 6987
rect 30389 6953 30423 6987
rect 30423 6953 30432 6987
rect 30380 6944 30432 6953
rect 37372 6944 37424 6996
rect 4068 6876 4120 6928
rect 2688 6808 2740 6860
rect 4160 6808 4212 6860
rect 3148 6740 3200 6792
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 1676 6715 1728 6724
rect 1676 6681 1685 6715
rect 1685 6681 1719 6715
rect 1719 6681 1728 6715
rect 1676 6672 1728 6681
rect 3240 6715 3292 6724
rect 3240 6681 3249 6715
rect 3249 6681 3283 6715
rect 3283 6681 3292 6715
rect 3240 6672 3292 6681
rect 3792 6672 3844 6724
rect 7840 6672 7892 6724
rect 3332 6604 3384 6656
rect 5540 6604 5592 6656
rect 9220 6715 9272 6724
rect 9220 6681 9229 6715
rect 9229 6681 9263 6715
rect 9263 6681 9272 6715
rect 9220 6672 9272 6681
rect 9772 6672 9824 6724
rect 12900 6808 12952 6860
rect 13452 6808 13504 6860
rect 15200 6876 15252 6928
rect 20996 6808 21048 6860
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 11060 6672 11112 6724
rect 12072 6672 12124 6724
rect 12440 6715 12492 6724
rect 12440 6681 12449 6715
rect 12449 6681 12483 6715
rect 12483 6681 12492 6715
rect 12440 6672 12492 6681
rect 12716 6672 12768 6724
rect 12900 6672 12952 6724
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 10508 6604 10560 6656
rect 12164 6604 12216 6656
rect 16580 6740 16632 6792
rect 18512 6715 18564 6724
rect 18512 6681 18521 6715
rect 18521 6681 18555 6715
rect 18555 6681 18564 6715
rect 18512 6672 18564 6681
rect 19616 6672 19668 6724
rect 23480 6740 23532 6792
rect 25136 6740 25188 6792
rect 27252 6808 27304 6860
rect 26056 6783 26108 6792
rect 26056 6749 26065 6783
rect 26065 6749 26099 6783
rect 26099 6749 26108 6783
rect 26056 6740 26108 6749
rect 26148 6783 26200 6792
rect 26148 6749 26157 6783
rect 26157 6749 26191 6783
rect 26191 6749 26200 6783
rect 26148 6740 26200 6749
rect 21364 6672 21416 6724
rect 25412 6672 25464 6724
rect 27436 6672 27488 6724
rect 29092 6783 29144 6792
rect 29092 6749 29101 6783
rect 29101 6749 29135 6783
rect 29135 6749 29144 6783
rect 29092 6740 29144 6749
rect 29276 6783 29328 6792
rect 29276 6749 29285 6783
rect 29285 6749 29319 6783
rect 29319 6749 29328 6783
rect 29276 6740 29328 6749
rect 33140 6808 33192 6860
rect 35808 6851 35860 6860
rect 35808 6817 35817 6851
rect 35817 6817 35851 6851
rect 35851 6817 35860 6851
rect 35808 6808 35860 6817
rect 36360 6851 36412 6860
rect 36360 6817 36369 6851
rect 36369 6817 36403 6851
rect 36403 6817 36412 6851
rect 36360 6808 36412 6817
rect 38476 6851 38528 6860
rect 38476 6817 38485 6851
rect 38485 6817 38519 6851
rect 38519 6817 38528 6851
rect 38476 6808 38528 6817
rect 31944 6740 31996 6792
rect 32680 6783 32732 6792
rect 32680 6749 32689 6783
rect 32689 6749 32723 6783
rect 32723 6749 32732 6783
rect 32680 6740 32732 6749
rect 32956 6740 33008 6792
rect 33416 6783 33468 6792
rect 33416 6749 33425 6783
rect 33425 6749 33459 6783
rect 33459 6749 33468 6783
rect 33416 6740 33468 6749
rect 33508 6783 33560 6792
rect 33508 6749 33518 6783
rect 33518 6749 33552 6783
rect 33552 6749 33560 6783
rect 33508 6740 33560 6749
rect 33784 6783 33836 6792
rect 33784 6749 33793 6783
rect 33793 6749 33827 6783
rect 33827 6749 33836 6783
rect 33784 6740 33836 6749
rect 33876 6740 33928 6792
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 22560 6604 22612 6656
rect 24400 6604 24452 6656
rect 29368 6604 29420 6656
rect 32312 6715 32364 6724
rect 32312 6681 32321 6715
rect 32321 6681 32355 6715
rect 32355 6681 32364 6715
rect 32312 6672 32364 6681
rect 33324 6672 33376 6724
rect 33692 6715 33744 6724
rect 33692 6681 33701 6715
rect 33701 6681 33735 6715
rect 33735 6681 33744 6715
rect 33692 6672 33744 6681
rect 35348 6740 35400 6792
rect 32404 6604 32456 6656
rect 37464 6672 37516 6724
rect 34796 6604 34848 6656
rect 35440 6647 35492 6656
rect 35440 6613 35449 6647
rect 35449 6613 35483 6647
rect 35483 6613 35492 6647
rect 35440 6604 35492 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 7748 6400 7800 6452
rect 848 6264 900 6316
rect 1676 6196 1728 6248
rect 2872 6196 2924 6248
rect 3332 6264 3384 6316
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 3240 6196 3292 6248
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 9220 6400 9272 6452
rect 9956 6400 10008 6452
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 8116 6264 8168 6316
rect 10140 6332 10192 6384
rect 10876 6400 10928 6452
rect 11704 6400 11756 6452
rect 8024 6196 8076 6248
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 5264 6171 5316 6180
rect 5264 6137 5273 6171
rect 5273 6137 5307 6171
rect 5307 6137 5316 6171
rect 5264 6128 5316 6137
rect 4712 6103 4764 6112
rect 4712 6069 4721 6103
rect 4721 6069 4755 6103
rect 4755 6069 4764 6103
rect 4712 6060 4764 6069
rect 8300 6128 8352 6180
rect 9128 6196 9180 6248
rect 10508 6264 10560 6316
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 11796 6332 11848 6384
rect 11520 6264 11572 6316
rect 12072 6332 12124 6384
rect 23020 6400 23072 6452
rect 23480 6400 23532 6452
rect 24400 6443 24452 6452
rect 24400 6409 24409 6443
rect 24409 6409 24443 6443
rect 24443 6409 24452 6443
rect 24400 6400 24452 6409
rect 24492 6400 24544 6452
rect 12532 6332 12584 6384
rect 24676 6332 24728 6384
rect 26056 6400 26108 6452
rect 27252 6443 27304 6452
rect 27252 6409 27261 6443
rect 27261 6409 27295 6443
rect 27295 6409 27304 6443
rect 27252 6400 27304 6409
rect 29276 6400 29328 6452
rect 25412 6332 25464 6384
rect 9312 6128 9364 6180
rect 10784 6171 10836 6180
rect 10784 6137 10793 6171
rect 10793 6137 10827 6171
rect 10827 6137 10836 6171
rect 10784 6128 10836 6137
rect 12256 6128 12308 6180
rect 12808 6264 12860 6316
rect 12992 6264 13044 6316
rect 14096 6264 14148 6316
rect 16672 6264 16724 6316
rect 18512 6264 18564 6316
rect 22008 6264 22060 6316
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 23204 6196 23256 6248
rect 24216 6264 24268 6316
rect 24860 6264 24912 6316
rect 25044 6264 25096 6316
rect 25136 6307 25188 6316
rect 25136 6273 25145 6307
rect 25145 6273 25179 6307
rect 25179 6273 25188 6307
rect 25136 6264 25188 6273
rect 25228 6307 25280 6316
rect 25228 6273 25237 6307
rect 25237 6273 25271 6307
rect 25271 6273 25280 6307
rect 25228 6264 25280 6273
rect 25320 6307 25372 6316
rect 25320 6273 25329 6307
rect 25329 6273 25363 6307
rect 25363 6273 25372 6307
rect 25320 6264 25372 6273
rect 25504 6307 25556 6316
rect 25504 6273 25513 6307
rect 25513 6273 25547 6307
rect 25547 6273 25556 6307
rect 25504 6264 25556 6273
rect 25964 6307 26016 6316
rect 25964 6273 25973 6307
rect 25973 6273 26007 6307
rect 26007 6273 26016 6307
rect 25964 6264 26016 6273
rect 26148 6264 26200 6316
rect 27436 6332 27488 6384
rect 26792 6307 26844 6316
rect 26792 6273 26801 6307
rect 26801 6273 26835 6307
rect 26835 6273 26844 6307
rect 26792 6264 26844 6273
rect 24768 6196 24820 6248
rect 12440 6128 12492 6180
rect 22652 6128 22704 6180
rect 26792 6128 26844 6180
rect 27712 6239 27764 6248
rect 27712 6205 27721 6239
rect 27721 6205 27755 6239
rect 27755 6205 27764 6239
rect 29000 6264 29052 6316
rect 27712 6196 27764 6205
rect 29368 6307 29420 6316
rect 29368 6273 29377 6307
rect 29377 6273 29411 6307
rect 29411 6273 29420 6307
rect 29368 6264 29420 6273
rect 30656 6307 30708 6316
rect 30656 6273 30665 6307
rect 30665 6273 30699 6307
rect 30699 6273 30708 6307
rect 30656 6264 30708 6273
rect 31300 6375 31352 6384
rect 31300 6341 31309 6375
rect 31309 6341 31343 6375
rect 31343 6341 31352 6375
rect 31300 6332 31352 6341
rect 33324 6443 33376 6452
rect 33324 6409 33333 6443
rect 33333 6409 33367 6443
rect 33367 6409 33376 6443
rect 33324 6400 33376 6409
rect 36452 6400 36504 6452
rect 31852 6332 31904 6384
rect 31576 6307 31628 6316
rect 31576 6273 31585 6307
rect 31585 6273 31619 6307
rect 31619 6273 31628 6307
rect 31576 6264 31628 6273
rect 31576 6128 31628 6180
rect 32404 6307 32456 6316
rect 32404 6273 32413 6307
rect 32413 6273 32447 6307
rect 32447 6273 32456 6307
rect 32404 6264 32456 6273
rect 32772 6264 32824 6316
rect 33140 6307 33192 6316
rect 33140 6273 33149 6307
rect 33149 6273 33183 6307
rect 33183 6273 33192 6307
rect 33140 6264 33192 6273
rect 34612 6307 34664 6316
rect 34612 6273 34621 6307
rect 34621 6273 34655 6307
rect 34655 6273 34664 6307
rect 34612 6264 34664 6273
rect 34796 6307 34848 6316
rect 34796 6273 34803 6307
rect 34803 6273 34848 6307
rect 34796 6264 34848 6273
rect 35440 6332 35492 6384
rect 33324 6196 33376 6248
rect 34428 6196 34480 6248
rect 34796 6128 34848 6180
rect 35624 6264 35676 6316
rect 35348 6196 35400 6248
rect 35992 6264 36044 6316
rect 8208 6060 8260 6112
rect 8760 6060 8812 6112
rect 10692 6060 10744 6112
rect 10968 6060 11020 6112
rect 11244 6060 11296 6112
rect 11980 6103 12032 6112
rect 11980 6069 11989 6103
rect 11989 6069 12023 6103
rect 12023 6069 12032 6103
rect 11980 6060 12032 6069
rect 22744 6060 22796 6112
rect 25044 6060 25096 6112
rect 26424 6060 26476 6112
rect 32036 6060 32088 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5540 5856 5592 5908
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 2596 5720 2648 5772
rect 4712 5720 4764 5772
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 9128 5856 9180 5908
rect 848 5652 900 5704
rect 3148 5584 3200 5636
rect 3884 5652 3936 5704
rect 5632 5695 5684 5704
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 6000 5652 6052 5704
rect 6552 5652 6604 5704
rect 7564 5652 7616 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8116 5652 8168 5704
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 8576 5627 8628 5636
rect 8576 5593 8585 5627
rect 8585 5593 8619 5627
rect 8619 5593 8628 5627
rect 8576 5584 8628 5593
rect 9220 5627 9272 5636
rect 9220 5593 9229 5627
rect 9229 5593 9263 5627
rect 9263 5593 9272 5627
rect 9220 5584 9272 5593
rect 9312 5627 9364 5636
rect 9312 5593 9321 5627
rect 9321 5593 9355 5627
rect 9355 5593 9364 5627
rect 9312 5584 9364 5593
rect 2964 5516 3016 5568
rect 3700 5516 3752 5568
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 6092 5559 6144 5568
rect 6092 5525 6101 5559
rect 6101 5525 6135 5559
rect 6135 5525 6144 5559
rect 6092 5516 6144 5525
rect 7104 5516 7156 5568
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 9588 5627 9640 5636
rect 9588 5593 9597 5627
rect 9597 5593 9631 5627
rect 9631 5593 9640 5627
rect 9588 5584 9640 5593
rect 11152 5788 11204 5840
rect 11428 5899 11480 5908
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 22836 5856 22888 5908
rect 26792 5899 26844 5908
rect 26792 5865 26801 5899
rect 26801 5865 26835 5899
rect 26835 5865 26844 5899
rect 26792 5856 26844 5865
rect 27712 5856 27764 5908
rect 30656 5856 30708 5908
rect 32312 5856 32364 5908
rect 33140 5856 33192 5908
rect 33876 5856 33928 5908
rect 34428 5899 34480 5908
rect 34428 5865 34437 5899
rect 34437 5865 34471 5899
rect 34471 5865 34480 5899
rect 34428 5856 34480 5865
rect 34612 5856 34664 5908
rect 35440 5856 35492 5908
rect 35624 5899 35676 5908
rect 35624 5865 35633 5899
rect 35633 5865 35667 5899
rect 35667 5865 35676 5899
rect 35624 5856 35676 5865
rect 22376 5788 22428 5840
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 12900 5720 12952 5729
rect 21732 5763 21784 5772
rect 21732 5729 21741 5763
rect 21741 5729 21775 5763
rect 21775 5729 21784 5763
rect 21732 5720 21784 5729
rect 22560 5763 22612 5772
rect 22560 5729 22569 5763
rect 22569 5729 22603 5763
rect 22603 5729 22612 5763
rect 22560 5720 22612 5729
rect 22836 5720 22888 5772
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 10692 5652 10744 5704
rect 11152 5652 11204 5704
rect 11888 5652 11940 5704
rect 11428 5584 11480 5636
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 12532 5652 12584 5704
rect 13360 5652 13412 5704
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 16672 5652 16724 5704
rect 22652 5652 22704 5704
rect 23020 5652 23072 5704
rect 12716 5584 12768 5636
rect 22008 5584 22060 5636
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 23204 5695 23256 5704
rect 23204 5661 23213 5695
rect 23213 5661 23247 5695
rect 23247 5661 23256 5695
rect 23204 5652 23256 5661
rect 23480 5652 23532 5704
rect 24308 5720 24360 5772
rect 25136 5831 25188 5840
rect 25136 5797 25145 5831
rect 25145 5797 25179 5831
rect 25179 5797 25188 5831
rect 25136 5788 25188 5797
rect 23848 5652 23900 5704
rect 25320 5720 25372 5772
rect 11888 5516 11940 5568
rect 13360 5516 13412 5568
rect 21180 5559 21232 5568
rect 21180 5525 21189 5559
rect 21189 5525 21223 5559
rect 21223 5525 21232 5559
rect 21180 5516 21232 5525
rect 23296 5559 23348 5568
rect 23296 5525 23305 5559
rect 23305 5525 23339 5559
rect 23339 5525 23348 5559
rect 23296 5516 23348 5525
rect 25044 5652 25096 5704
rect 24676 5627 24728 5636
rect 24676 5593 24685 5627
rect 24685 5593 24719 5627
rect 24719 5593 24728 5627
rect 24676 5584 24728 5593
rect 25228 5584 25280 5636
rect 25596 5584 25648 5636
rect 26056 5652 26108 5704
rect 26424 5695 26476 5704
rect 26424 5661 26433 5695
rect 26433 5661 26467 5695
rect 26467 5661 26476 5695
rect 26424 5652 26476 5661
rect 27344 5652 27396 5704
rect 31852 5695 31904 5704
rect 31852 5661 31861 5695
rect 31861 5661 31895 5695
rect 31895 5661 31904 5695
rect 31852 5652 31904 5661
rect 32036 5695 32088 5704
rect 32036 5661 32045 5695
rect 32045 5661 32079 5695
rect 32079 5661 32088 5695
rect 32036 5652 32088 5661
rect 32404 5652 32456 5704
rect 32772 5695 32824 5704
rect 32772 5661 32781 5695
rect 32781 5661 32815 5695
rect 32815 5661 32824 5695
rect 32772 5652 32824 5661
rect 33784 5695 33836 5704
rect 33784 5661 33793 5695
rect 33793 5661 33827 5695
rect 33827 5661 33836 5695
rect 33784 5652 33836 5661
rect 33876 5652 33928 5704
rect 34796 5720 34848 5772
rect 34520 5695 34572 5704
rect 34520 5661 34529 5695
rect 34529 5661 34563 5695
rect 34563 5661 34572 5695
rect 34520 5652 34572 5661
rect 34704 5695 34756 5704
rect 34704 5661 34713 5695
rect 34713 5661 34747 5695
rect 34747 5661 34756 5695
rect 34704 5652 34756 5661
rect 24860 5516 24912 5568
rect 25044 5559 25096 5568
rect 25044 5525 25053 5559
rect 25053 5525 25087 5559
rect 25087 5525 25096 5559
rect 25044 5516 25096 5525
rect 25964 5516 26016 5568
rect 27160 5627 27212 5636
rect 27160 5593 27169 5627
rect 27169 5593 27203 5627
rect 27203 5593 27212 5627
rect 27160 5584 27212 5593
rect 29736 5627 29788 5636
rect 29736 5593 29745 5627
rect 29745 5593 29779 5627
rect 29779 5593 29788 5627
rect 29736 5584 29788 5593
rect 29828 5584 29880 5636
rect 35072 5695 35124 5704
rect 35072 5661 35081 5695
rect 35081 5661 35115 5695
rect 35115 5661 35124 5695
rect 35072 5652 35124 5661
rect 35348 5695 35400 5704
rect 35348 5661 35357 5695
rect 35357 5661 35391 5695
rect 35391 5661 35400 5695
rect 35348 5652 35400 5661
rect 35808 5652 35860 5704
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 3792 5312 3844 5364
rect 4160 5244 4212 5296
rect 5632 5312 5684 5364
rect 6920 5312 6972 5364
rect 7380 5312 7432 5364
rect 10508 5312 10560 5364
rect 13360 5355 13412 5364
rect 13360 5321 13369 5355
rect 13369 5321 13403 5355
rect 13403 5321 13412 5355
rect 13360 5312 13412 5321
rect 22008 5355 22060 5364
rect 22008 5321 22017 5355
rect 22017 5321 22051 5355
rect 22051 5321 22060 5355
rect 22008 5312 22060 5321
rect 4804 5244 4856 5296
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 3700 5176 3752 5228
rect 6184 5176 6236 5228
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 7380 5219 7432 5228
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 11980 5287 12032 5296
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 12900 5244 12952 5296
rect 7932 5176 7984 5228
rect 8300 5176 8352 5228
rect 848 5108 900 5160
rect 5724 5108 5776 5160
rect 8208 5108 8260 5160
rect 8392 5108 8444 5160
rect 9496 5176 9548 5228
rect 9864 5176 9916 5228
rect 11244 5176 11296 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 9680 5108 9732 5160
rect 12808 5176 12860 5228
rect 21364 5244 21416 5296
rect 22652 5312 22704 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 24308 5312 24360 5364
rect 9588 5040 9640 5092
rect 18512 5176 18564 5228
rect 13728 5108 13780 5160
rect 21180 5108 21232 5160
rect 22376 5219 22428 5228
rect 22376 5185 22385 5219
rect 22385 5185 22419 5219
rect 22419 5185 22428 5219
rect 22376 5176 22428 5185
rect 23296 5244 23348 5296
rect 24860 5287 24912 5296
rect 24860 5253 24869 5287
rect 24869 5253 24903 5287
rect 24903 5253 24912 5287
rect 24860 5244 24912 5253
rect 25136 5244 25188 5296
rect 29736 5312 29788 5364
rect 29828 5312 29880 5364
rect 31576 5312 31628 5364
rect 25596 5287 25648 5296
rect 25596 5253 25605 5287
rect 25605 5253 25639 5287
rect 25639 5253 25648 5287
rect 25596 5244 25648 5253
rect 22744 5219 22796 5228
rect 22744 5185 22753 5219
rect 22753 5185 22787 5219
rect 22787 5185 22796 5219
rect 22744 5176 22796 5185
rect 22836 5176 22888 5228
rect 23940 5176 23992 5228
rect 25228 5219 25280 5228
rect 25228 5185 25237 5219
rect 25237 5185 25271 5219
rect 25271 5185 25280 5219
rect 25228 5176 25280 5185
rect 29368 5219 29420 5228
rect 29368 5185 29377 5219
rect 29377 5185 29411 5219
rect 29411 5185 29420 5219
rect 29368 5176 29420 5185
rect 21732 5040 21784 5092
rect 24492 5040 24544 5092
rect 25412 5108 25464 5160
rect 28172 5108 28224 5160
rect 29184 5151 29236 5160
rect 29184 5117 29193 5151
rect 29193 5117 29227 5151
rect 29227 5117 29236 5151
rect 30840 5219 30892 5228
rect 30840 5185 30849 5219
rect 30849 5185 30883 5219
rect 30883 5185 30892 5219
rect 30840 5176 30892 5185
rect 29184 5108 29236 5117
rect 25964 5040 26016 5092
rect 31576 5219 31628 5228
rect 31576 5185 31585 5219
rect 31585 5185 31619 5219
rect 31619 5185 31628 5219
rect 31576 5176 31628 5185
rect 32772 5312 32824 5364
rect 33324 5355 33376 5364
rect 33324 5321 33349 5355
rect 33349 5321 33376 5355
rect 33324 5312 33376 5321
rect 33784 5312 33836 5364
rect 34704 5312 34756 5364
rect 35072 5312 35124 5364
rect 33140 5287 33192 5296
rect 33140 5253 33149 5287
rect 33149 5253 33183 5287
rect 33183 5253 33192 5287
rect 33140 5244 33192 5253
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 6828 4972 6880 5024
rect 9404 5015 9456 5024
rect 9404 4981 9413 5015
rect 9413 4981 9447 5015
rect 9447 4981 9456 5015
rect 9404 4972 9456 4981
rect 11244 4972 11296 5024
rect 12164 5015 12216 5024
rect 12164 4981 12173 5015
rect 12173 4981 12207 5015
rect 12207 4981 12216 5015
rect 12164 4972 12216 4981
rect 12348 5015 12400 5024
rect 12348 4981 12357 5015
rect 12357 4981 12391 5015
rect 12391 4981 12400 5015
rect 12348 4972 12400 4981
rect 12624 4972 12676 5024
rect 22192 5015 22244 5024
rect 22192 4981 22201 5015
rect 22201 4981 22235 5015
rect 22235 4981 22244 5015
rect 22192 4972 22244 4981
rect 25780 5015 25832 5024
rect 25780 4981 25789 5015
rect 25789 4981 25823 5015
rect 25823 4981 25832 5015
rect 25780 4972 25832 4981
rect 28632 4972 28684 5024
rect 29828 5083 29880 5092
rect 29828 5049 29837 5083
rect 29837 5049 29871 5083
rect 29871 5049 29880 5083
rect 29828 5040 29880 5049
rect 33324 5176 33376 5228
rect 34152 5176 34204 5228
rect 34060 5108 34112 5160
rect 34796 5176 34848 5228
rect 35348 5176 35400 5228
rect 33876 5083 33928 5092
rect 33876 5049 33885 5083
rect 33885 5049 33919 5083
rect 33919 5049 33928 5083
rect 33876 5040 33928 5049
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 8300 4811 8352 4820
rect 8300 4777 8309 4811
rect 8309 4777 8343 4811
rect 8343 4777 8352 4811
rect 8300 4768 8352 4777
rect 8484 4768 8536 4820
rect 9036 4768 9088 4820
rect 9680 4811 9732 4820
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 3976 4700 4028 4752
rect 4068 4632 4120 4684
rect 5356 4632 5408 4684
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 23480 4768 23532 4820
rect 25228 4768 25280 4820
rect 9220 4632 9272 4684
rect 12164 4675 12216 4684
rect 12164 4641 12173 4675
rect 12173 4641 12207 4675
rect 12207 4641 12216 4675
rect 12164 4632 12216 4641
rect 15844 4632 15896 4684
rect 18512 4632 18564 4684
rect 21732 4632 21784 4684
rect 3792 4564 3844 4616
rect 5540 4564 5592 4616
rect 6092 4564 6144 4616
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 4252 4539 4304 4548
rect 4252 4505 4261 4539
rect 4261 4505 4295 4539
rect 4295 4505 4304 4539
rect 4252 4496 4304 4505
rect 7932 4564 7984 4616
rect 6920 4496 6972 4548
rect 8576 4496 8628 4548
rect 9588 4564 9640 4616
rect 11336 4564 11388 4616
rect 12532 4564 12584 4616
rect 22284 4564 22336 4616
rect 26240 4700 26292 4752
rect 23756 4632 23808 4684
rect 27620 4768 27672 4820
rect 27804 4700 27856 4752
rect 29368 4768 29420 4820
rect 33876 4768 33928 4820
rect 34060 4811 34112 4820
rect 34060 4777 34069 4811
rect 34069 4777 34103 4811
rect 34103 4777 34112 4811
rect 34060 4768 34112 4777
rect 34152 4811 34204 4820
rect 34152 4777 34161 4811
rect 34161 4777 34195 4811
rect 34195 4777 34204 4811
rect 34152 4768 34204 4777
rect 35348 4811 35400 4820
rect 35348 4777 35357 4811
rect 35357 4777 35391 4811
rect 35391 4777 35400 4811
rect 35348 4768 35400 4777
rect 30840 4700 30892 4752
rect 26424 4675 26476 4684
rect 26424 4641 26433 4675
rect 26433 4641 26467 4675
rect 26467 4641 26476 4675
rect 26424 4632 26476 4641
rect 11428 4496 11480 4548
rect 13636 4539 13688 4548
rect 13636 4505 13645 4539
rect 13645 4505 13679 4539
rect 13679 4505 13688 4539
rect 13636 4496 13688 4505
rect 13728 4496 13780 4548
rect 19984 4496 20036 4548
rect 22008 4496 22060 4548
rect 848 4428 900 4480
rect 4620 4428 4672 4480
rect 22376 4496 22428 4548
rect 22744 4539 22796 4548
rect 22744 4505 22753 4539
rect 22753 4505 22787 4539
rect 22787 4505 22796 4539
rect 23388 4607 23440 4616
rect 23388 4573 23397 4607
rect 23397 4573 23431 4607
rect 23431 4573 23440 4607
rect 23388 4564 23440 4573
rect 22744 4496 22796 4505
rect 23112 4539 23164 4548
rect 23112 4505 23121 4539
rect 23121 4505 23155 4539
rect 23155 4505 23164 4539
rect 23112 4496 23164 4505
rect 23940 4607 23992 4616
rect 23940 4573 23949 4607
rect 23949 4573 23983 4607
rect 23983 4573 23992 4607
rect 23940 4564 23992 4573
rect 24860 4564 24912 4616
rect 25320 4564 25372 4616
rect 26700 4564 26752 4616
rect 26884 4564 26936 4616
rect 26976 4496 27028 4548
rect 27896 4632 27948 4684
rect 28632 4675 28684 4684
rect 28632 4641 28641 4675
rect 28641 4641 28675 4675
rect 28675 4641 28684 4675
rect 28632 4632 28684 4641
rect 33508 4632 33560 4684
rect 27436 4607 27488 4616
rect 27436 4573 27445 4607
rect 27445 4573 27479 4607
rect 27479 4573 27488 4607
rect 27436 4564 27488 4573
rect 28172 4564 28224 4616
rect 33416 4564 33468 4616
rect 34796 4564 34848 4616
rect 23756 4428 23808 4480
rect 23848 4428 23900 4480
rect 26240 4471 26292 4480
rect 26240 4437 26249 4471
rect 26249 4437 26283 4471
rect 26283 4437 26292 4471
rect 26240 4428 26292 4437
rect 26608 4428 26660 4480
rect 27528 4496 27580 4548
rect 27620 4496 27672 4548
rect 28724 4496 28776 4548
rect 34060 4496 34112 4548
rect 27252 4428 27304 4480
rect 28080 4428 28132 4480
rect 34704 4471 34756 4480
rect 34704 4437 34713 4471
rect 34713 4437 34747 4471
rect 34747 4437 34756 4471
rect 34704 4428 34756 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4160 4224 4212 4276
rect 4252 4224 4304 4276
rect 10416 4224 10468 4276
rect 12348 4224 12400 4276
rect 13636 4224 13688 4276
rect 22284 4224 22336 4276
rect 23112 4224 23164 4276
rect 24308 4224 24360 4276
rect 25412 4224 25464 4276
rect 4804 4156 4856 4208
rect 11428 4156 11480 4208
rect 12164 4156 12216 4208
rect 22008 4156 22060 4208
rect 5816 4088 5868 4140
rect 6000 4088 6052 4140
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 7104 4088 7156 4140
rect 7564 4088 7616 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 3516 4063 3568 4072
rect 3516 4029 3525 4063
rect 3525 4029 3559 4063
rect 3559 4029 3568 4063
rect 3516 4020 3568 4029
rect 5540 4020 5592 4072
rect 9496 3952 9548 4004
rect 9680 3952 9732 4004
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 11888 4088 11940 4140
rect 12348 4088 12400 4140
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 21732 4088 21784 4140
rect 21824 4020 21876 4072
rect 23848 4199 23900 4208
rect 23848 4165 23857 4199
rect 23857 4165 23891 4199
rect 23891 4165 23900 4199
rect 23848 4156 23900 4165
rect 23940 4156 23992 4208
rect 24032 4131 24084 4140
rect 24032 4097 24041 4131
rect 24041 4097 24075 4131
rect 24075 4097 24084 4131
rect 24032 4088 24084 4097
rect 24400 4088 24452 4140
rect 23756 3952 23808 4004
rect 24124 3995 24176 4004
rect 24124 3961 24133 3995
rect 24133 3961 24167 3995
rect 24167 3961 24176 3995
rect 24124 3952 24176 3961
rect 25780 4156 25832 4208
rect 26240 4224 26292 4276
rect 26332 4224 26384 4276
rect 27252 4224 27304 4276
rect 24676 3952 24728 4004
rect 25320 4131 25372 4140
rect 25320 4097 25329 4131
rect 25329 4097 25363 4131
rect 25363 4097 25372 4131
rect 25320 4088 25372 4097
rect 25688 4088 25740 4140
rect 24860 4063 24912 4072
rect 24860 4029 24869 4063
rect 24869 4029 24903 4063
rect 24903 4029 24912 4063
rect 24860 4020 24912 4029
rect 25044 4063 25096 4072
rect 25044 4029 25053 4063
rect 25053 4029 25087 4063
rect 25087 4029 25096 4063
rect 25044 4020 25096 4029
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5540 3884 5592 3936
rect 5632 3884 5684 3936
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 7288 3884 7340 3936
rect 9956 3884 10008 3936
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 10968 3927 11020 3936
rect 10968 3893 10977 3927
rect 10977 3893 11011 3927
rect 11011 3893 11020 3927
rect 10968 3884 11020 3893
rect 22376 3927 22428 3936
rect 22376 3893 22385 3927
rect 22385 3893 22419 3927
rect 22419 3893 22428 3927
rect 22376 3884 22428 3893
rect 22744 3884 22796 3936
rect 26884 4156 26936 4208
rect 27804 4199 27856 4208
rect 27804 4165 27813 4199
rect 27813 4165 27847 4199
rect 27847 4165 27856 4199
rect 27804 4156 27856 4165
rect 28172 4267 28224 4276
rect 28172 4233 28181 4267
rect 28181 4233 28215 4267
rect 28215 4233 28224 4267
rect 28172 4224 28224 4233
rect 28632 4224 28684 4276
rect 31576 4224 31628 4276
rect 30840 4156 30892 4208
rect 33416 4224 33468 4276
rect 33508 4267 33560 4276
rect 33508 4233 33517 4267
rect 33517 4233 33551 4267
rect 33551 4233 33560 4267
rect 33508 4224 33560 4233
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 27528 4063 27580 4072
rect 27528 4029 27537 4063
rect 27537 4029 27571 4063
rect 27571 4029 27580 4063
rect 27528 4020 27580 4029
rect 27712 3952 27764 4004
rect 27620 3884 27672 3936
rect 29552 4131 29604 4140
rect 29552 4097 29561 4131
rect 29561 4097 29595 4131
rect 29595 4097 29604 4131
rect 29552 4088 29604 4097
rect 29828 4131 29880 4140
rect 29828 4097 29837 4131
rect 29837 4097 29871 4131
rect 29871 4097 29880 4131
rect 29828 4088 29880 4097
rect 29092 4063 29144 4072
rect 29092 4029 29101 4063
rect 29101 4029 29135 4063
rect 29135 4029 29144 4063
rect 29092 4020 29144 4029
rect 29184 4063 29236 4072
rect 29184 4029 29193 4063
rect 29193 4029 29227 4063
rect 29227 4029 29236 4063
rect 29184 4020 29236 4029
rect 30932 4020 30984 4072
rect 29000 3952 29052 4004
rect 31116 4088 31168 4140
rect 31484 4131 31536 4140
rect 31484 4097 31493 4131
rect 31493 4097 31527 4131
rect 31527 4097 31536 4131
rect 31484 4088 31536 4097
rect 31576 4131 31628 4140
rect 31576 4097 31585 4131
rect 31585 4097 31619 4131
rect 31619 4097 31628 4131
rect 31576 4088 31628 4097
rect 32036 4088 32088 4140
rect 32312 4020 32364 4072
rect 33140 4020 33192 4072
rect 28172 3884 28224 3936
rect 30656 3884 30708 3936
rect 31116 3884 31168 3936
rect 34704 3884 34756 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3516 3680 3568 3732
rect 3884 3680 3936 3732
rect 4620 3680 4672 3732
rect 4804 3680 4856 3732
rect 6092 3680 6144 3732
rect 7104 3723 7156 3732
rect 7104 3689 7113 3723
rect 7113 3689 7147 3723
rect 7147 3689 7156 3723
rect 7104 3680 7156 3689
rect 7840 3680 7892 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 11520 3680 11572 3732
rect 23388 3680 23440 3732
rect 23572 3680 23624 3732
rect 848 3612 900 3664
rect 7564 3612 7616 3664
rect 9588 3612 9640 3664
rect 4160 3544 4212 3596
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 5632 3587 5684 3596
rect 5632 3553 5641 3587
rect 5641 3553 5675 3587
rect 5675 3553 5684 3587
rect 5632 3544 5684 3553
rect 3884 3476 3936 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 4620 3476 4672 3528
rect 4988 3408 5040 3460
rect 7104 3476 7156 3528
rect 8300 3476 8352 3528
rect 5632 3408 5684 3460
rect 6092 3408 6144 3460
rect 8576 3408 8628 3460
rect 8668 3451 8720 3460
rect 8668 3417 8677 3451
rect 8677 3417 8711 3451
rect 8711 3417 8720 3451
rect 8668 3408 8720 3417
rect 3792 3340 3844 3392
rect 3976 3340 4028 3392
rect 4528 3383 4580 3392
rect 4528 3349 4537 3383
rect 4537 3349 4571 3383
rect 4571 3349 4580 3383
rect 4528 3340 4580 3349
rect 6368 3340 6420 3392
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 8300 3340 8352 3392
rect 8852 3476 8904 3528
rect 9220 3544 9272 3596
rect 10968 3612 11020 3664
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 11244 3612 11296 3664
rect 11888 3451 11940 3460
rect 11888 3417 11897 3451
rect 11897 3417 11931 3451
rect 11931 3417 11940 3451
rect 11888 3408 11940 3417
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 13268 3476 13320 3528
rect 12348 3408 12400 3460
rect 11796 3340 11848 3392
rect 22652 3408 22704 3460
rect 23020 3408 23072 3460
rect 24032 3680 24084 3732
rect 25412 3723 25464 3732
rect 25412 3689 25421 3723
rect 25421 3689 25455 3723
rect 25455 3689 25464 3723
rect 25412 3680 25464 3689
rect 27896 3723 27948 3732
rect 27896 3689 27905 3723
rect 27905 3689 27939 3723
rect 27939 3689 27948 3723
rect 27896 3680 27948 3689
rect 29828 3680 29880 3732
rect 30288 3723 30340 3732
rect 24860 3612 24912 3664
rect 24308 3544 24360 3596
rect 24768 3587 24820 3596
rect 24768 3553 24777 3587
rect 24777 3553 24811 3587
rect 24811 3553 24820 3587
rect 24768 3544 24820 3553
rect 24492 3476 24544 3528
rect 25320 3544 25372 3596
rect 26884 3587 26936 3596
rect 26884 3553 26893 3587
rect 26893 3553 26927 3587
rect 26927 3553 26936 3587
rect 29552 3612 29604 3664
rect 29736 3612 29788 3664
rect 30288 3689 30297 3723
rect 30297 3689 30331 3723
rect 30331 3689 30340 3723
rect 30288 3680 30340 3689
rect 30656 3680 30708 3732
rect 30748 3612 30800 3664
rect 26884 3544 26936 3553
rect 23756 3408 23808 3460
rect 25044 3408 25096 3460
rect 25688 3476 25740 3528
rect 26240 3519 26292 3528
rect 26240 3485 26249 3519
rect 26249 3485 26283 3519
rect 26283 3485 26292 3519
rect 26240 3476 26292 3485
rect 26424 3519 26476 3528
rect 26424 3485 26433 3519
rect 26433 3485 26467 3519
rect 26467 3485 26476 3519
rect 26424 3476 26476 3485
rect 25596 3451 25648 3460
rect 25596 3417 25605 3451
rect 25605 3417 25639 3451
rect 25639 3417 25648 3451
rect 25596 3408 25648 3417
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 30564 3544 30616 3596
rect 31024 3680 31076 3732
rect 31116 3723 31168 3732
rect 31116 3689 31125 3723
rect 31125 3689 31159 3723
rect 31159 3689 31168 3723
rect 31116 3680 31168 3689
rect 31300 3680 31352 3732
rect 32036 3723 32088 3732
rect 32036 3689 32045 3723
rect 32045 3689 32079 3723
rect 32079 3689 32088 3723
rect 32036 3680 32088 3689
rect 32312 3723 32364 3732
rect 32312 3689 32321 3723
rect 32321 3689 32355 3723
rect 32355 3689 32364 3723
rect 32312 3680 32364 3689
rect 27436 3519 27488 3528
rect 27436 3485 27445 3519
rect 27445 3485 27479 3519
rect 27479 3485 27488 3519
rect 27436 3476 27488 3485
rect 27620 3519 27672 3528
rect 27620 3485 27629 3519
rect 27629 3485 27663 3519
rect 27663 3485 27672 3519
rect 27620 3476 27672 3485
rect 27712 3519 27764 3528
rect 27712 3485 27721 3519
rect 27721 3485 27755 3519
rect 27755 3485 27764 3519
rect 27712 3476 27764 3485
rect 22192 3340 22244 3392
rect 24768 3340 24820 3392
rect 27068 3408 27120 3460
rect 28540 3519 28592 3528
rect 28540 3485 28549 3519
rect 28549 3485 28583 3519
rect 28583 3485 28592 3519
rect 28540 3476 28592 3485
rect 28724 3519 28776 3528
rect 28724 3485 28733 3519
rect 28733 3485 28767 3519
rect 28767 3485 28776 3519
rect 28724 3476 28776 3485
rect 26792 3340 26844 3392
rect 27160 3383 27212 3392
rect 27160 3349 27169 3383
rect 27169 3349 27203 3383
rect 27203 3349 27212 3383
rect 27160 3340 27212 3349
rect 29736 3519 29788 3528
rect 29736 3485 29745 3519
rect 29745 3485 29779 3519
rect 29779 3485 29788 3519
rect 29736 3476 29788 3485
rect 29184 3340 29236 3392
rect 30104 3451 30156 3460
rect 30104 3417 30113 3451
rect 30113 3417 30147 3451
rect 30147 3417 30156 3451
rect 30840 3476 30892 3528
rect 31024 3476 31076 3528
rect 31392 3519 31444 3528
rect 31392 3485 31401 3519
rect 31401 3485 31435 3519
rect 31435 3485 31444 3519
rect 31392 3476 31444 3485
rect 31484 3476 31536 3528
rect 31668 3519 31720 3528
rect 31668 3485 31677 3519
rect 31677 3485 31711 3519
rect 31711 3485 31720 3519
rect 31668 3476 31720 3485
rect 30104 3408 30156 3417
rect 31300 3408 31352 3460
rect 32312 3519 32364 3528
rect 32312 3485 32321 3519
rect 32321 3485 32355 3519
rect 32355 3485 32364 3519
rect 32312 3476 32364 3485
rect 38476 3519 38528 3528
rect 38476 3485 38485 3519
rect 38485 3485 38519 3519
rect 38519 3485 38528 3519
rect 38476 3476 38528 3485
rect 30748 3340 30800 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 4528 3136 4580 3188
rect 5632 3179 5684 3188
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 8300 3136 8352 3188
rect 4160 3068 4212 3120
rect 4804 3068 4856 3120
rect 5724 3000 5776 3052
rect 7196 3068 7248 3120
rect 8760 3068 8812 3120
rect 9220 3111 9272 3120
rect 9220 3077 9229 3111
rect 9229 3077 9263 3111
rect 9263 3077 9272 3111
rect 9220 3068 9272 3077
rect 13268 3179 13320 3188
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 9772 3068 9824 3120
rect 11796 3111 11848 3120
rect 11796 3077 11805 3111
rect 11805 3077 11839 3111
rect 11839 3077 11848 3111
rect 11796 3068 11848 3077
rect 12532 3068 12584 3120
rect 25596 3136 25648 3188
rect 26608 3136 26660 3188
rect 27712 3136 27764 3188
rect 30104 3179 30156 3188
rect 30104 3145 30113 3179
rect 30113 3145 30147 3179
rect 30147 3145 30156 3179
rect 30104 3136 30156 3145
rect 848 2932 900 2984
rect 7104 3000 7156 3052
rect 22744 3068 22796 3120
rect 23756 3068 23808 3120
rect 7932 2932 7984 2984
rect 8760 2932 8812 2984
rect 5816 2864 5868 2916
rect 3976 2796 4028 2848
rect 7104 2796 7156 2848
rect 9588 2975 9640 2984
rect 9588 2941 9597 2975
rect 9597 2941 9631 2975
rect 9631 2941 9640 2975
rect 9588 2932 9640 2941
rect 10508 2932 10560 2984
rect 11060 2796 11112 2848
rect 23020 2932 23072 2984
rect 24124 3043 24176 3052
rect 24124 3009 24133 3043
rect 24133 3009 24167 3043
rect 24167 3009 24176 3043
rect 24124 3000 24176 3009
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 24768 3000 24820 3052
rect 26792 3000 26844 3052
rect 27068 3000 27120 3052
rect 27160 3043 27212 3052
rect 27160 3009 27181 3043
rect 27181 3009 27212 3043
rect 30288 3068 30340 3120
rect 27160 3000 27212 3009
rect 24400 2796 24452 2848
rect 28172 2975 28224 2984
rect 28172 2941 28181 2975
rect 28181 2941 28215 2975
rect 28215 2941 28224 2975
rect 28172 2932 28224 2941
rect 28540 2932 28592 2984
rect 29092 2932 29144 2984
rect 32312 3136 32364 3188
rect 31576 3068 31628 3120
rect 30748 3043 30800 3052
rect 30748 3009 30757 3043
rect 30757 3009 30791 3043
rect 30791 3009 30800 3043
rect 30748 3000 30800 3009
rect 30932 3000 30984 3052
rect 31300 3043 31352 3052
rect 31300 3009 31309 3043
rect 31309 3009 31343 3043
rect 31343 3009 31352 3043
rect 31300 3000 31352 3009
rect 31484 3000 31536 3052
rect 30564 2932 30616 2984
rect 31668 2932 31720 2984
rect 38476 2975 38528 2984
rect 38476 2941 38485 2975
rect 38485 2941 38519 2975
rect 38519 2941 38528 2975
rect 38476 2932 38528 2941
rect 26976 2864 27028 2916
rect 31392 2864 31444 2916
rect 30288 2796 30340 2848
rect 34796 2796 34848 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8576 2592 8628 2644
rect 14924 2592 14976 2644
rect 5448 2456 5500 2508
rect 7288 2456 7340 2508
rect 8484 2456 8536 2508
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 7932 2320 7984 2372
rect 21364 2431 21416 2440
rect 21364 2397 21373 2431
rect 21373 2397 21407 2431
rect 21407 2397 21416 2431
rect 21364 2388 21416 2397
rect 23848 2388 23900 2440
rect 29644 2388 29696 2440
rect 30288 2388 30340 2440
rect 35440 2388 35492 2440
rect 36084 2388 36136 2440
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 21272 2252 21324 2304
rect 24492 2252 24544 2304
rect 27068 2252 27120 2304
rect 27712 2252 27764 2304
rect 29000 2252 29052 2304
rect 38476 2295 38528 2304
rect 38476 2261 38485 2295
rect 38485 2261 38519 2295
rect 38519 2261 38528 2295
rect 38476 2252 38528 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 3238 39200 3294 40000
rect 5170 39200 5226 40000
rect 23846 39200 23902 40000
rect 25778 39200 25834 40000
rect 26422 39200 26478 40000
rect 27066 39200 27122 40000
rect 27710 39200 27766 40000
rect 28354 39200 28410 40000
rect 28998 39200 29054 40000
rect 29642 39200 29698 40000
rect 30286 39200 30342 40000
rect 30930 39200 30986 40000
rect 31574 39200 31630 40000
rect 32218 39200 32274 40000
rect 32862 39200 32918 40000
rect 33506 39200 33562 40000
rect 34150 39200 34206 40000
rect 34794 39200 34850 40000
rect 35438 39200 35494 40000
rect 36082 39200 36138 40000
rect 36726 39200 36782 40000
rect 38566 39536 38622 39545
rect 38566 39471 38622 39480
rect 1306 37496 1362 37505
rect 3252 37466 3280 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 1306 37431 1308 37440
rect 1360 37431 1362 37440
rect 3240 37460 3292 37466
rect 1308 37402 1360 37408
rect 3240 37402 3292 37408
rect 848 37324 900 37330
rect 848 37266 900 37272
rect 860 36961 888 37266
rect 5184 37262 5212 39200
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 6828 37120 6880 37126
rect 6828 37062 6880 37068
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 846 36952 902 36961
rect 4874 36955 5182 36964
rect 846 36887 902 36896
rect 5724 36848 5776 36854
rect 5724 36790 5776 36796
rect 5172 36712 5224 36718
rect 5172 36654 5224 36660
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 5184 36378 5212 36654
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 848 36304 900 36310
rect 846 36272 848 36281
rect 5264 36304 5316 36310
rect 900 36272 902 36281
rect 5264 36246 5316 36252
rect 846 36207 902 36216
rect 3332 36236 3384 36242
rect 3332 36178 3384 36184
rect 848 35624 900 35630
rect 846 35592 848 35601
rect 900 35592 902 35601
rect 846 35527 902 35536
rect 3240 35488 3292 35494
rect 3240 35430 3292 35436
rect 2872 35148 2924 35154
rect 2872 35090 2924 35096
rect 848 35080 900 35086
rect 848 35022 900 35028
rect 860 34921 888 35022
rect 846 34912 902 34921
rect 846 34847 902 34856
rect 2884 34678 2912 35090
rect 3252 35086 3280 35430
rect 3344 35154 3372 36178
rect 4436 36168 4488 36174
rect 4436 36110 4488 36116
rect 4448 35834 4476 36110
rect 4712 36032 4764 36038
rect 4712 35974 4764 35980
rect 4436 35828 4488 35834
rect 4436 35770 4488 35776
rect 4724 35630 4752 35974
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 5276 35698 5304 36246
rect 5460 36230 5672 36258
rect 5460 35834 5488 36230
rect 5644 36174 5672 36230
rect 5632 36168 5684 36174
rect 5632 36110 5684 36116
rect 5540 36100 5592 36106
rect 5540 36042 5592 36048
rect 5552 35834 5580 36042
rect 5448 35828 5500 35834
rect 5448 35770 5500 35776
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5264 35692 5316 35698
rect 5264 35634 5316 35640
rect 4712 35624 4764 35630
rect 5460 35578 5488 35770
rect 4712 35566 4764 35572
rect 4620 35488 4672 35494
rect 4620 35430 4672 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3976 35284 4028 35290
rect 3976 35226 4028 35232
rect 3332 35148 3384 35154
rect 3332 35090 3384 35096
rect 3240 35080 3292 35086
rect 3240 35022 3292 35028
rect 2872 34672 2924 34678
rect 2872 34614 2924 34620
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 110 33824 166 33833
rect 110 33759 166 33768
rect 124 19446 152 33759
rect 2240 33454 2268 34478
rect 3240 33992 3292 33998
rect 3344 33980 3372 35090
rect 3884 34740 3936 34746
rect 3884 34682 3936 34688
rect 3292 33952 3372 33980
rect 3424 33992 3476 33998
rect 3240 33934 3292 33940
rect 3424 33934 3476 33940
rect 2504 33856 2556 33862
rect 2504 33798 2556 33804
rect 2516 33590 2544 33798
rect 2504 33584 2556 33590
rect 2504 33526 2556 33532
rect 2228 33448 2280 33454
rect 2228 33390 2280 33396
rect 2240 32026 2268 33390
rect 3252 33318 3280 33934
rect 3436 33658 3464 33934
rect 3424 33652 3476 33658
rect 3424 33594 3476 33600
rect 3240 33312 3292 33318
rect 3240 33254 3292 33260
rect 3436 32910 3464 33594
rect 3792 33584 3844 33590
rect 3792 33526 3844 33532
rect 3424 32904 3476 32910
rect 3424 32846 3476 32852
rect 3436 32298 3464 32846
rect 3700 32768 3752 32774
rect 3700 32710 3752 32716
rect 3712 32450 3740 32710
rect 3804 32586 3832 33526
rect 3896 32978 3924 34682
rect 3988 34610 4016 35226
rect 4632 35154 4660 35430
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 4344 35080 4396 35086
rect 4344 35022 4396 35028
rect 4356 34678 4384 35022
rect 4344 34672 4396 34678
rect 4344 34614 4396 34620
rect 3976 34604 4028 34610
rect 3976 34546 4028 34552
rect 3884 32972 3936 32978
rect 3884 32914 3936 32920
rect 3988 32774 4016 34546
rect 4724 34406 4752 35566
rect 5276 35550 5488 35578
rect 5276 34950 5304 35550
rect 5736 35290 5764 36790
rect 6552 36712 6604 36718
rect 6552 36654 6604 36660
rect 6184 36576 6236 36582
rect 6184 36518 6236 36524
rect 6196 36174 6224 36518
rect 6184 36168 6236 36174
rect 6184 36110 6236 36116
rect 6564 35698 6592 36654
rect 6840 36174 6868 37062
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 7208 36378 7236 36654
rect 8128 36582 8156 37198
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 21180 37188 21232 37194
rect 21180 37130 21232 37136
rect 19616 37120 19668 37126
rect 19616 37062 19668 37068
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 8392 36780 8444 36786
rect 8392 36722 8444 36728
rect 8944 36780 8996 36786
rect 8944 36722 8996 36728
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 8116 36576 8168 36582
rect 8116 36518 8168 36524
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7300 36258 7328 36518
rect 7472 36372 7524 36378
rect 7472 36314 7524 36320
rect 8116 36372 8168 36378
rect 8116 36314 8168 36320
rect 7208 36230 7328 36258
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 6828 36168 6880 36174
rect 6828 36110 6880 36116
rect 6552 35692 6604 35698
rect 6552 35634 6604 35640
rect 6092 35624 6144 35630
rect 6092 35566 6144 35572
rect 6104 35290 6132 35566
rect 5724 35284 5776 35290
rect 5724 35226 5776 35232
rect 6092 35284 6144 35290
rect 6092 35226 6144 35232
rect 5736 35086 5764 35226
rect 5724 35080 5776 35086
rect 5724 35022 5776 35028
rect 5264 34944 5316 34950
rect 5264 34886 5316 34892
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4712 34400 4764 34406
rect 4712 34342 4764 34348
rect 5080 34400 5132 34406
rect 5080 34342 5132 34348
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5092 34066 5120 34342
rect 5080 34060 5132 34066
rect 5080 34002 5132 34008
rect 4528 33992 4580 33998
rect 4528 33934 4580 33940
rect 4540 33454 4568 33934
rect 5276 33844 5304 34886
rect 5632 34400 5684 34406
rect 5632 34342 5684 34348
rect 5644 34202 5672 34342
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 6104 34134 6132 35226
rect 6564 34610 6592 35634
rect 6656 35086 6684 36110
rect 7208 36106 7236 36230
rect 7196 36100 7248 36106
rect 7196 36042 7248 36048
rect 7208 35086 7236 36042
rect 7288 35760 7340 35766
rect 7288 35702 7340 35708
rect 6644 35080 6696 35086
rect 6644 35022 6696 35028
rect 7196 35080 7248 35086
rect 7196 35022 7248 35028
rect 6552 34604 6604 34610
rect 6552 34546 6604 34552
rect 6368 34536 6420 34542
rect 6368 34478 6420 34484
rect 6092 34128 6144 34134
rect 6092 34070 6144 34076
rect 5356 33992 5408 33998
rect 5408 33940 5672 33946
rect 5356 33934 5672 33940
rect 5368 33918 5672 33934
rect 6104 33930 6132 34070
rect 5448 33856 5500 33862
rect 5276 33816 5448 33844
rect 5448 33798 5500 33804
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4620 33516 4672 33522
rect 4620 33458 4672 33464
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 4528 33448 4580 33454
rect 4528 33390 4580 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 32994 4660 33458
rect 4540 32966 4660 32994
rect 3976 32768 4028 32774
rect 3976 32710 4028 32716
rect 3804 32558 3924 32586
rect 4540 32570 4568 32966
rect 4724 32570 4752 33458
rect 5644 33454 5672 33918
rect 6092 33924 6144 33930
rect 6092 33866 6144 33872
rect 5724 33856 5776 33862
rect 5724 33798 5776 33804
rect 5632 33448 5684 33454
rect 5632 33390 5684 33396
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 4908 33114 4936 33254
rect 4896 33108 4948 33114
rect 4896 33050 4948 33056
rect 5644 32774 5672 33390
rect 5736 33318 5764 33798
rect 5724 33312 5776 33318
rect 5724 33254 5776 33260
rect 6000 33312 6052 33318
rect 6000 33254 6052 33260
rect 6012 32978 6040 33254
rect 6000 32972 6052 32978
rect 6000 32914 6052 32920
rect 5632 32768 5684 32774
rect 5632 32710 5684 32716
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 3712 32422 3832 32450
rect 3424 32292 3476 32298
rect 3424 32234 3476 32240
rect 2228 32020 2280 32026
rect 2228 31962 2280 31968
rect 2504 32020 2556 32026
rect 2504 31962 2556 31968
rect 2240 31346 2268 31962
rect 2516 31890 2544 31962
rect 2504 31884 2556 31890
rect 2504 31826 2556 31832
rect 3804 31822 3832 32422
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3804 31482 3832 31758
rect 3792 31476 3844 31482
rect 3792 31418 3844 31424
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 3608 31272 3660 31278
rect 3608 31214 3660 31220
rect 3620 30938 3648 31214
rect 3608 30932 3660 30938
rect 3608 30874 3660 30880
rect 3792 30252 3844 30258
rect 3792 30194 3844 30200
rect 846 30152 902 30161
rect 846 30087 848 30096
rect 900 30087 902 30096
rect 848 30058 900 30064
rect 848 29640 900 29646
rect 848 29582 900 29588
rect 3332 29640 3384 29646
rect 3332 29582 3384 29588
rect 860 29481 888 29582
rect 846 29472 902 29481
rect 846 29407 902 29416
rect 3344 29102 3372 29582
rect 3424 29504 3476 29510
rect 3424 29446 3476 29452
rect 3436 29238 3464 29446
rect 3424 29232 3476 29238
rect 3424 29174 3476 29180
rect 848 29096 900 29102
rect 848 29038 900 29044
rect 3332 29096 3384 29102
rect 3332 29038 3384 29044
rect 3700 29096 3752 29102
rect 3700 29038 3752 29044
rect 860 28801 888 29038
rect 2964 28960 3016 28966
rect 2964 28902 3016 28908
rect 846 28792 902 28801
rect 846 28727 902 28736
rect 2976 28558 3004 28902
rect 3344 28558 3372 29038
rect 3712 28762 3740 29038
rect 3700 28756 3752 28762
rect 3700 28698 3752 28704
rect 3804 28642 3832 30194
rect 3896 30122 3924 32558
rect 3976 32564 4028 32570
rect 3976 32506 4028 32512
rect 4528 32564 4580 32570
rect 4528 32506 4580 32512
rect 4712 32564 4764 32570
rect 4712 32506 4764 32512
rect 3988 31754 4016 32506
rect 5644 32366 5672 32710
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4804 32360 4856 32366
rect 4804 32302 4856 32308
rect 5632 32360 5684 32366
rect 5632 32302 5684 32308
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 31958 4660 32302
rect 4620 31952 4672 31958
rect 4620 31894 4672 31900
rect 3988 31748 4120 31754
rect 3988 31726 4068 31748
rect 4068 31690 4120 31696
rect 4080 30734 4108 31690
rect 4620 31204 4672 31210
rect 4620 31146 4672 31152
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30734 4660 31146
rect 4816 31142 4844 32302
rect 6276 32292 6328 32298
rect 6276 32234 6328 32240
rect 5356 32224 5408 32230
rect 5356 32166 5408 32172
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4804 31136 4856 31142
rect 4804 31078 4856 31084
rect 4816 30870 4844 31078
rect 4804 30864 4856 30870
rect 4804 30806 4856 30812
rect 5368 30802 5396 32166
rect 6288 31958 6316 32234
rect 6276 31952 6328 31958
rect 6276 31894 6328 31900
rect 5816 31680 5868 31686
rect 5816 31622 5868 31628
rect 5724 31408 5776 31414
rect 5724 31350 5776 31356
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5356 30796 5408 30802
rect 5356 30738 5408 30744
rect 4068 30728 4120 30734
rect 4068 30670 4120 30676
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 4080 30394 4108 30670
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 3884 30116 3936 30122
rect 3884 30058 3936 30064
rect 3896 29578 3924 30058
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 3884 29572 3936 29578
rect 3884 29514 3936 29520
rect 4252 29504 4304 29510
rect 4252 29446 4304 29452
rect 4264 29170 4292 29446
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 4252 29164 4304 29170
rect 4252 29106 4304 29112
rect 4080 28694 4108 29106
rect 4724 29102 4752 29650
rect 4816 29238 4844 30670
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5460 30258 5488 31078
rect 5736 30666 5764 31350
rect 5828 31346 5856 31622
rect 5816 31340 5868 31346
rect 5816 31282 5868 31288
rect 5724 30660 5776 30666
rect 5724 30602 5776 30608
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 5736 30002 5764 30602
rect 5828 30258 5856 31282
rect 5816 30252 5868 30258
rect 5816 30194 5868 30200
rect 5736 29974 5856 30002
rect 5264 29708 5316 29714
rect 5264 29650 5316 29656
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4816 29102 4844 29174
rect 4712 29096 4764 29102
rect 4712 29038 4764 29044
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3712 28614 3832 28642
rect 4068 28688 4120 28694
rect 4068 28630 4120 28636
rect 4816 28626 4844 29038
rect 4804 28620 4856 28626
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 3332 28552 3384 28558
rect 3332 28494 3384 28500
rect 3608 28552 3660 28558
rect 3608 28494 3660 28500
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 1412 27470 1440 27950
rect 2792 27470 2820 28086
rect 3148 27940 3200 27946
rect 3148 27882 3200 27888
rect 2872 27872 2924 27878
rect 2872 27814 2924 27820
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 2780 27464 2832 27470
rect 2780 27406 2832 27412
rect 1412 25362 1440 27406
rect 1676 27396 1728 27402
rect 1676 27338 1728 27344
rect 1688 26926 1716 27338
rect 2884 27146 2912 27814
rect 3160 27470 3188 27882
rect 3344 27538 3372 28494
rect 3620 28150 3648 28494
rect 3608 28144 3660 28150
rect 3608 28086 3660 28092
rect 3424 28008 3476 28014
rect 3424 27950 3476 27956
rect 3436 27674 3464 27950
rect 3620 27674 3648 28086
rect 3424 27668 3476 27674
rect 3424 27610 3476 27616
rect 3608 27668 3660 27674
rect 3608 27610 3660 27616
rect 3436 27554 3464 27610
rect 3332 27532 3384 27538
rect 3436 27526 3648 27554
rect 3332 27474 3384 27480
rect 3620 27470 3648 27526
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3608 27464 3660 27470
rect 3608 27406 3660 27412
rect 2792 27118 2912 27146
rect 1676 26920 1728 26926
rect 1676 26862 1728 26868
rect 2792 26382 2820 27118
rect 2780 26376 2832 26382
rect 2780 26318 2832 26324
rect 2688 26308 2740 26314
rect 2688 26250 2740 26256
rect 2700 25362 2728 26250
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 2688 25356 2740 25362
rect 2688 25298 2740 25304
rect 3068 25294 3096 27406
rect 3160 26926 3188 27406
rect 3332 27328 3384 27334
rect 3332 27270 3384 27276
rect 3344 26994 3372 27270
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 3148 26920 3200 26926
rect 3148 26862 3200 26868
rect 3160 26586 3188 26862
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 3436 26382 3464 27066
rect 3332 26376 3384 26382
rect 3332 26318 3384 26324
rect 3424 26376 3476 26382
rect 3424 26318 3476 26324
rect 3344 25906 3372 26318
rect 3240 25900 3292 25906
rect 3240 25842 3292 25848
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 3148 25424 3200 25430
rect 3148 25366 3200 25372
rect 3056 25288 3108 25294
rect 1306 25256 1362 25265
rect 3056 25230 3108 25236
rect 1306 25191 1362 25200
rect 1768 25220 1820 25226
rect 1320 24682 1348 25191
rect 1768 25162 1820 25168
rect 2964 25220 3016 25226
rect 2964 25162 3016 25168
rect 1780 24750 1808 25162
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 1768 24744 1820 24750
rect 1768 24686 1820 24692
rect 2044 24744 2096 24750
rect 2044 24686 2096 24692
rect 1308 24676 1360 24682
rect 1308 24618 1360 24624
rect 2056 24614 2084 24686
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1676 23656 1728 23662
rect 1676 23598 1728 23604
rect 1412 22574 1440 23598
rect 1688 23322 1716 23598
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 2056 23118 2084 24550
rect 2044 23112 2096 23118
rect 2044 23054 2096 23060
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22710 2360 22918
rect 2320 22704 2372 22710
rect 2320 22646 2372 22652
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 2056 20466 2084 22510
rect 2884 21894 2912 24754
rect 2976 24614 3004 25162
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2976 24206 3004 24550
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2976 23866 3004 24142
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 3068 23798 3096 25230
rect 3160 25158 3188 25366
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3160 24750 3188 25094
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3160 24138 3188 24686
rect 3252 24410 3280 25842
rect 3344 25498 3372 25842
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 3436 24274 3464 24550
rect 3424 24268 3476 24274
rect 3424 24210 3476 24216
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3148 24132 3200 24138
rect 3148 24074 3200 24080
rect 3056 23792 3108 23798
rect 3056 23734 3108 23740
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 2976 23118 3004 23666
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 3068 22964 3096 23734
rect 3344 23730 3372 24142
rect 3608 24132 3660 24138
rect 3608 24074 3660 24080
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 3436 23254 3464 24006
rect 3620 23662 3648 24074
rect 3608 23656 3660 23662
rect 3608 23598 3660 23604
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 3148 22976 3200 22982
rect 3068 22936 3148 22964
rect 3068 22710 3096 22936
rect 3148 22918 3200 22924
rect 3056 22704 3108 22710
rect 3056 22646 3108 22652
rect 3712 21894 3740 28614
rect 4804 28562 4856 28568
rect 3792 28552 3844 28558
rect 3792 28494 3844 28500
rect 4068 28552 4120 28558
rect 4068 28494 4120 28500
rect 4712 28552 4764 28558
rect 5276 28506 5304 29650
rect 5828 29170 5856 29974
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 5816 29164 5868 29170
rect 5816 29106 5868 29112
rect 4712 28494 4764 28500
rect 3804 27878 3832 28494
rect 3976 28076 4028 28082
rect 3976 28018 4028 28024
rect 3792 27872 3844 27878
rect 3792 27814 3844 27820
rect 3988 27674 4016 28018
rect 4080 28014 4108 28494
rect 4724 28082 4752 28494
rect 5184 28490 5304 28506
rect 5828 28490 5856 29106
rect 6196 28966 6224 29582
rect 6380 29578 6408 34478
rect 6920 33992 6972 33998
rect 7300 33946 7328 35702
rect 7484 35290 7512 36314
rect 8128 36174 8156 36314
rect 8116 36168 8168 36174
rect 8116 36110 8168 36116
rect 7748 36032 7800 36038
rect 7748 35974 7800 35980
rect 7840 36032 7892 36038
rect 7840 35974 7892 35980
rect 7472 35284 7524 35290
rect 7472 35226 7524 35232
rect 7760 35154 7788 35974
rect 7852 35630 7880 35974
rect 8128 35834 8156 36110
rect 8116 35828 8168 35834
rect 8116 35770 8168 35776
rect 7840 35624 7892 35630
rect 7840 35566 7892 35572
rect 8024 35624 8076 35630
rect 8024 35566 8076 35572
rect 8036 35290 8064 35566
rect 8024 35284 8076 35290
rect 8024 35226 8076 35232
rect 7748 35148 7800 35154
rect 7748 35090 7800 35096
rect 7380 34944 7432 34950
rect 7380 34886 7432 34892
rect 7392 34202 7420 34886
rect 7380 34196 7432 34202
rect 7380 34138 7432 34144
rect 6920 33934 6972 33940
rect 6932 32570 6960 33934
rect 7208 33918 7328 33946
rect 7012 33856 7064 33862
rect 7012 33798 7064 33804
rect 7024 33590 7052 33798
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 7012 33584 7064 33590
rect 7012 33526 7064 33532
rect 7012 32836 7064 32842
rect 7012 32778 7064 32784
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 7024 32450 7052 32778
rect 7116 32570 7144 33594
rect 7104 32564 7156 32570
rect 7104 32506 7156 32512
rect 7208 32450 7236 33918
rect 8024 33856 8076 33862
rect 8024 33798 8076 33804
rect 7288 33516 7340 33522
rect 7288 33458 7340 33464
rect 7300 32978 7328 33458
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 7288 32972 7340 32978
rect 7288 32914 7340 32920
rect 7484 32774 7512 33390
rect 8036 32910 8064 33798
rect 8220 33538 8248 36722
rect 8404 36242 8432 36722
rect 8668 36576 8720 36582
rect 8668 36518 8720 36524
rect 8680 36242 8708 36518
rect 8956 36378 8984 36722
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 8944 36372 8996 36378
rect 8944 36314 8996 36320
rect 8392 36236 8444 36242
rect 8392 36178 8444 36184
rect 8668 36236 8720 36242
rect 8668 36178 8720 36184
rect 19260 36174 19288 36654
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 13084 35692 13136 35698
rect 13084 35634 13136 35640
rect 8392 35488 8444 35494
rect 8392 35430 8444 35436
rect 8404 35222 8432 35430
rect 8392 35216 8444 35222
rect 8392 35158 8444 35164
rect 8772 33930 8800 35634
rect 11060 35624 11112 35630
rect 11060 35566 11112 35572
rect 10876 35556 10928 35562
rect 10876 35498 10928 35504
rect 10784 35284 10836 35290
rect 10784 35226 10836 35232
rect 10796 34610 10824 35226
rect 10888 34610 10916 35498
rect 11072 35154 11100 35566
rect 12440 35488 12492 35494
rect 12440 35430 12492 35436
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 10968 35012 11020 35018
rect 10968 34954 11020 34960
rect 10980 34746 11008 34954
rect 10968 34740 11020 34746
rect 10968 34682 11020 34688
rect 9772 34604 9824 34610
rect 9772 34546 9824 34552
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 10876 34604 10928 34610
rect 10876 34546 10928 34552
rect 9220 34536 9272 34542
rect 9220 34478 9272 34484
rect 8760 33924 8812 33930
rect 8760 33866 8812 33872
rect 9232 33862 9260 34478
rect 9220 33856 9272 33862
rect 9220 33798 9272 33804
rect 8128 33522 8248 33538
rect 8116 33516 8248 33522
rect 8168 33510 8248 33516
rect 8116 33458 8168 33464
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 7472 32768 7524 32774
rect 7472 32710 7524 32716
rect 7564 32768 7616 32774
rect 7564 32710 7616 32716
rect 7484 32502 7512 32710
rect 6644 32428 6696 32434
rect 6644 32370 6696 32376
rect 6920 32428 6972 32434
rect 7024 32422 7236 32450
rect 7472 32496 7524 32502
rect 7472 32438 7524 32444
rect 7576 32434 7604 32710
rect 7564 32428 7616 32434
rect 6920 32370 6972 32376
rect 6656 32026 6684 32370
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6932 31890 6960 32370
rect 6552 31884 6604 31890
rect 6552 31826 6604 31832
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 6564 31754 6592 31826
rect 6736 31816 6788 31822
rect 6736 31758 6788 31764
rect 6564 31726 6684 31754
rect 6656 31346 6684 31726
rect 6748 31686 6776 31758
rect 6736 31680 6788 31686
rect 6736 31622 6788 31628
rect 6748 31482 6776 31622
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 6644 31340 6696 31346
rect 6644 31282 6696 31288
rect 6748 30938 6776 31418
rect 6840 31346 6868 31418
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 6736 30932 6788 30938
rect 6736 30874 6788 30880
rect 6828 30252 6880 30258
rect 6828 30194 6880 30200
rect 6840 29578 6868 30194
rect 7116 30122 7144 32422
rect 7564 32370 7616 32376
rect 7288 31884 7340 31890
rect 7288 31826 7340 31832
rect 7300 31754 7328 31826
rect 7576 31822 7604 32370
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7748 31816 7800 31822
rect 7748 31758 7800 31764
rect 7196 31748 7248 31754
rect 7196 31690 7248 31696
rect 7288 31748 7340 31754
rect 7288 31690 7340 31696
rect 7656 31748 7708 31754
rect 7656 31690 7708 31696
rect 7208 31414 7236 31690
rect 7196 31408 7248 31414
rect 7196 31350 7248 31356
rect 7208 30734 7236 31350
rect 7300 31210 7328 31690
rect 7564 31680 7616 31686
rect 7564 31622 7616 31628
rect 7576 31346 7604 31622
rect 7564 31340 7616 31346
rect 7564 31282 7616 31288
rect 7380 31272 7432 31278
rect 7380 31214 7432 31220
rect 7288 31204 7340 31210
rect 7288 31146 7340 31152
rect 7196 30728 7248 30734
rect 7300 30716 7328 31146
rect 7392 30938 7420 31214
rect 7380 30932 7432 30938
rect 7380 30874 7432 30880
rect 7668 30734 7696 31690
rect 7760 31482 7788 31758
rect 7748 31476 7800 31482
rect 7748 31418 7800 31424
rect 8128 31346 8156 33458
rect 9232 33454 9260 33798
rect 9784 33590 9812 34546
rect 9956 34536 10008 34542
rect 9956 34478 10008 34484
rect 9680 33584 9732 33590
rect 9680 33526 9732 33532
rect 9772 33584 9824 33590
rect 9772 33526 9824 33532
rect 8852 33448 8904 33454
rect 8852 33390 8904 33396
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 9496 33448 9548 33454
rect 9496 33390 9548 33396
rect 8576 33312 8628 33318
rect 8576 33254 8628 33260
rect 8588 32910 8616 33254
rect 8864 32978 8892 33390
rect 8852 32972 8904 32978
rect 8852 32914 8904 32920
rect 8576 32904 8628 32910
rect 8576 32846 8628 32852
rect 9508 32434 9536 33390
rect 9692 33114 9720 33526
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9968 32910 9996 34478
rect 10232 34400 10284 34406
rect 10232 34342 10284 34348
rect 10324 34400 10376 34406
rect 10324 34342 10376 34348
rect 10244 33658 10272 34342
rect 10336 34066 10364 34342
rect 10324 34060 10376 34066
rect 10324 34002 10376 34008
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9772 32496 9824 32502
rect 9772 32438 9824 32444
rect 9496 32428 9548 32434
rect 9496 32370 9548 32376
rect 8116 31340 8168 31346
rect 8116 31282 8168 31288
rect 7380 30728 7432 30734
rect 7300 30688 7380 30716
rect 7196 30670 7248 30676
rect 7380 30670 7432 30676
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7392 30394 7420 30670
rect 8128 30410 8156 31282
rect 9508 31278 9536 32370
rect 9496 31272 9548 31278
rect 9496 31214 9548 31220
rect 9508 30802 9536 31214
rect 9496 30796 9548 30802
rect 9496 30738 9548 30744
rect 9036 30592 9088 30598
rect 9036 30534 9088 30540
rect 7380 30388 7432 30394
rect 7380 30330 7432 30336
rect 8036 30382 8156 30410
rect 8036 30326 8064 30382
rect 9048 30326 9076 30534
rect 8024 30320 8076 30326
rect 8024 30262 8076 30268
rect 9036 30320 9088 30326
rect 9036 30262 9088 30268
rect 7104 30116 7156 30122
rect 7104 30058 7156 30064
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6828 29572 6880 29578
rect 6828 29514 6880 29520
rect 6184 28960 6236 28966
rect 6184 28902 6236 28908
rect 5172 28484 5304 28490
rect 5224 28478 5304 28484
rect 5172 28426 5224 28432
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5276 28150 5304 28478
rect 5816 28484 5868 28490
rect 5816 28426 5868 28432
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5264 28144 5316 28150
rect 5264 28086 5316 28092
rect 4620 28076 4672 28082
rect 4620 28018 4672 28024
rect 4712 28076 4764 28082
rect 4712 28018 4764 28024
rect 4068 28008 4120 28014
rect 4068 27950 4120 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 3988 27130 4016 27610
rect 4632 27470 4660 28018
rect 5460 27878 5488 28358
rect 6196 27946 6224 28902
rect 6184 27940 6236 27946
rect 6184 27882 6236 27888
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 5264 27396 5316 27402
rect 5264 27338 5316 27344
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 3976 27124 4028 27130
rect 3976 27066 4028 27072
rect 5276 26926 5304 27338
rect 6380 27334 6408 29514
rect 6840 29170 6868 29514
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 7116 29102 7144 30058
rect 7472 29640 7524 29646
rect 7656 29640 7708 29646
rect 7472 29582 7524 29588
rect 7576 29600 7656 29628
rect 7380 29504 7432 29510
rect 7380 29446 7432 29452
rect 7392 29238 7420 29446
rect 7380 29232 7432 29238
rect 7380 29174 7432 29180
rect 7104 29096 7156 29102
rect 7104 29038 7156 29044
rect 7484 28762 7512 29582
rect 7472 28756 7524 28762
rect 7472 28698 7524 28704
rect 7012 28688 7064 28694
rect 7012 28630 7064 28636
rect 6736 28620 6788 28626
rect 6736 28562 6788 28568
rect 6644 28416 6696 28422
rect 6644 28358 6696 28364
rect 6656 28218 6684 28358
rect 6644 28212 6696 28218
rect 6644 28154 6696 28160
rect 6748 28082 6776 28562
rect 6920 28552 6972 28558
rect 6920 28494 6972 28500
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6932 28014 6960 28494
rect 7024 28150 7052 28630
rect 7380 28620 7432 28626
rect 7380 28562 7432 28568
rect 7012 28144 7064 28150
rect 7012 28086 7064 28092
rect 6920 28008 6972 28014
rect 6920 27950 6972 27956
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 6368 27328 6420 27334
rect 6368 27270 6420 27276
rect 3976 26920 4028 26926
rect 3976 26862 4028 26868
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 3988 26586 4016 26862
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5276 26586 5304 26862
rect 3976 26580 4028 26586
rect 3976 26522 4028 26528
rect 5264 26580 5316 26586
rect 5264 26522 5316 26528
rect 5276 26450 5304 26522
rect 5264 26444 5316 26450
rect 5264 26386 5316 26392
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 4080 25362 4108 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4724 24886 4752 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3896 22574 3924 24686
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3988 23526 4016 24346
rect 4724 24274 4752 24822
rect 4988 24336 5040 24342
rect 4986 24304 4988 24313
rect 5040 24304 5042 24313
rect 4712 24268 4764 24274
rect 4986 24239 5042 24248
rect 4712 24210 4764 24216
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 3976 23520 4028 23526
rect 3976 23462 4028 23468
rect 3988 23118 4016 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5184 23322 5212 23802
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5172 23316 5224 23322
rect 5172 23258 5224 23264
rect 5184 23118 5212 23258
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 5172 23112 5224 23118
rect 5172 23054 5224 23060
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 3896 22098 3924 22510
rect 3988 22438 4016 23054
rect 4068 22976 4120 22982
rect 4908 22964 4936 23054
rect 4068 22918 4120 22924
rect 4816 22936 4936 22964
rect 5172 22976 5224 22982
rect 4080 22710 4108 22918
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3884 22092 3936 22098
rect 4080 22094 4108 22646
rect 4816 22574 4844 22936
rect 5368 22964 5396 23598
rect 5224 22936 5396 22964
rect 5172 22918 5224 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4080 22066 4200 22094
rect 3884 22034 3936 22040
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 2792 20534 2820 20742
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2056 19922 2084 20402
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 1676 19780 1728 19786
rect 1676 19722 1728 19728
rect 112 19440 164 19446
rect 112 19382 164 19388
rect 1688 19310 1716 19722
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 2792 18272 2820 19790
rect 2884 19446 2912 20878
rect 3712 20874 3740 21830
rect 3700 20868 3752 20874
rect 3700 20810 3752 20816
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3436 20602 3464 20742
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3712 20058 3740 20198
rect 3804 20058 3832 21966
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 21622 4016 21830
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 4172 21350 4200 22066
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4632 21622 4660 22034
rect 4724 21690 4752 22510
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 4816 21554 4844 22510
rect 5368 22438 5396 22936
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5184 22030 5212 22170
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5368 21554 5396 22374
rect 5460 22234 5488 27270
rect 6276 27056 6328 27062
rect 6276 26998 6328 27004
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 5816 26784 5868 26790
rect 5816 26726 5868 26732
rect 5632 26240 5684 26246
rect 5632 26182 5684 26188
rect 5644 25974 5672 26182
rect 5632 25968 5684 25974
rect 5632 25910 5684 25916
rect 5828 25906 5856 26726
rect 6104 25906 6132 26930
rect 6288 26314 6316 26998
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6276 26308 6328 26314
rect 6276 26250 6328 26256
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 6092 25900 6144 25906
rect 6092 25842 6144 25848
rect 6000 25832 6052 25838
rect 6000 25774 6052 25780
rect 6012 25430 6040 25774
rect 6092 25492 6144 25498
rect 6092 25434 6144 25440
rect 6000 25424 6052 25430
rect 6000 25366 6052 25372
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5644 24410 5672 25230
rect 5724 25152 5776 25158
rect 5724 25094 5776 25100
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5736 24750 5764 25094
rect 5724 24744 5776 24750
rect 5724 24686 5776 24692
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5724 23112 5776 23118
rect 5920 23066 5948 25094
rect 6012 24426 6040 25366
rect 6104 24954 6132 25434
rect 6184 25220 6236 25226
rect 6184 25162 6236 25168
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 6104 24614 6132 24890
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 6012 24398 6132 24426
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 6012 23118 6040 23598
rect 6104 23118 6132 24398
rect 6196 24206 6224 25162
rect 6288 24886 6316 26250
rect 6380 26246 6408 26930
rect 6368 26240 6420 26246
rect 6368 26182 6420 26188
rect 6380 25838 6408 26182
rect 6368 25832 6420 25838
rect 6368 25774 6420 25780
rect 6380 25226 6408 25774
rect 6828 25764 6880 25770
rect 6828 25706 6880 25712
rect 6840 25294 6868 25706
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6276 24880 6328 24886
rect 6276 24822 6328 24828
rect 6380 24818 6408 25162
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 6380 24070 6408 24754
rect 6932 24614 6960 27814
rect 7024 27470 7052 28086
rect 7392 28014 7420 28562
rect 7472 28484 7524 28490
rect 7472 28426 7524 28432
rect 7380 28008 7432 28014
rect 7380 27950 7432 27956
rect 7288 27600 7340 27606
rect 7288 27542 7340 27548
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 7012 26308 7064 26314
rect 7012 26250 7064 26256
rect 7024 25498 7052 26250
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 7116 25294 7144 25638
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7300 24750 7328 27542
rect 7484 27470 7512 28426
rect 7576 28218 7604 29600
rect 7656 29582 7708 29588
rect 8036 29306 8064 30262
rect 9508 30258 9536 30738
rect 9784 30598 9812 32438
rect 10232 32360 10284 32366
rect 10232 32302 10284 32308
rect 10244 32026 10272 32302
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10428 31822 10456 33526
rect 10796 33114 10824 34546
rect 10784 33108 10836 33114
rect 10784 33050 10836 33056
rect 10888 32026 10916 34546
rect 11072 34066 11100 35090
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11716 34678 11744 34886
rect 12452 34678 12480 35430
rect 13096 35290 13124 35634
rect 13636 35624 13688 35630
rect 13636 35566 13688 35572
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 13084 35284 13136 35290
rect 13084 35226 13136 35232
rect 12728 35086 12756 35226
rect 13544 35148 13596 35154
rect 13544 35090 13596 35096
rect 12716 35080 12768 35086
rect 12636 35040 12716 35068
rect 12636 34746 12664 35040
rect 12716 35022 12768 35028
rect 13452 35080 13504 35086
rect 13452 35022 13504 35028
rect 13084 34944 13136 34950
rect 13084 34886 13136 34892
rect 12624 34740 12676 34746
rect 12624 34682 12676 34688
rect 11704 34672 11756 34678
rect 11704 34614 11756 34620
rect 12440 34672 12492 34678
rect 12440 34614 12492 34620
rect 13096 34542 13124 34886
rect 12164 34536 12216 34542
rect 12164 34478 12216 34484
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 11612 34400 11664 34406
rect 11612 34342 11664 34348
rect 11060 34060 11112 34066
rect 11060 34002 11112 34008
rect 11624 33930 11652 34342
rect 12176 34066 12204 34478
rect 13096 34202 13124 34478
rect 13464 34202 13492 35022
rect 13556 34610 13584 35090
rect 13648 34660 13676 35566
rect 17040 35284 17092 35290
rect 17040 35226 17092 35232
rect 16304 35216 16356 35222
rect 16304 35158 16356 35164
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 15660 35080 15712 35086
rect 15660 35022 15712 35028
rect 13924 34746 13952 35022
rect 15016 35012 15068 35018
rect 15016 34954 15068 34960
rect 15292 35012 15344 35018
rect 15292 34954 15344 34960
rect 13912 34740 13964 34746
rect 13912 34682 13964 34688
rect 13728 34672 13780 34678
rect 13648 34632 13728 34660
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 13084 34196 13136 34202
rect 13084 34138 13136 34144
rect 13452 34196 13504 34202
rect 13452 34138 13504 34144
rect 12164 34060 12216 34066
rect 12164 34002 12216 34008
rect 11612 33924 11664 33930
rect 11612 33866 11664 33872
rect 11060 33584 11112 33590
rect 11060 33526 11112 33532
rect 10968 33516 11020 33522
rect 10968 33458 11020 33464
rect 10980 33114 11008 33458
rect 10968 33108 11020 33114
rect 10968 33050 11020 33056
rect 11072 33046 11100 33526
rect 11796 33108 11848 33114
rect 11796 33050 11848 33056
rect 11060 33040 11112 33046
rect 11060 32982 11112 32988
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 10508 32020 10560 32026
rect 10508 31962 10560 31968
rect 10876 32020 10928 32026
rect 10876 31962 10928 31968
rect 10520 31890 10548 31962
rect 10508 31884 10560 31890
rect 10508 31826 10560 31832
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10520 31362 10548 31826
rect 10692 31748 10744 31754
rect 10968 31748 11020 31754
rect 10744 31708 10968 31736
rect 10692 31690 10744 31696
rect 10968 31690 11020 31696
rect 10428 31334 10548 31362
rect 10428 31278 10456 31334
rect 10416 31272 10468 31278
rect 10416 31214 10468 31220
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10152 30666 10180 31078
rect 10140 30660 10192 30666
rect 10140 30602 10192 30608
rect 10232 30660 10284 30666
rect 10232 30602 10284 30608
rect 9772 30592 9824 30598
rect 9772 30534 9824 30540
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 9232 29714 9260 29990
rect 9220 29708 9272 29714
rect 9220 29650 9272 29656
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 8944 29640 8996 29646
rect 8944 29582 8996 29588
rect 8024 29300 8076 29306
rect 8024 29242 8076 29248
rect 8128 29034 8156 29582
rect 8116 29028 8168 29034
rect 8116 28970 8168 28976
rect 8128 28558 8156 28970
rect 8208 28756 8260 28762
rect 8208 28698 8260 28704
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8220 28490 8248 28698
rect 8956 28626 8984 29582
rect 10244 29578 10272 30602
rect 10428 30258 10456 31214
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10428 29714 10456 30194
rect 10876 30184 10928 30190
rect 10876 30126 10928 30132
rect 10416 29708 10468 29714
rect 10416 29650 10468 29656
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9416 29170 9444 29446
rect 10244 29306 10272 29514
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 8944 28620 8996 28626
rect 8944 28562 8996 28568
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 7564 28212 7616 28218
rect 7564 28154 7616 28160
rect 7576 27674 7604 28154
rect 8220 28014 8248 28426
rect 8956 28234 8984 28562
rect 10244 28490 10272 29242
rect 9588 28484 9640 28490
rect 9588 28426 9640 28432
rect 10232 28484 10284 28490
rect 10232 28426 10284 28432
rect 8864 28218 8984 28234
rect 9600 28218 9628 28426
rect 8852 28212 8984 28218
rect 8904 28206 8984 28212
rect 9588 28212 9640 28218
rect 8852 28154 8904 28160
rect 9588 28154 9640 28160
rect 10244 28150 10272 28426
rect 10232 28144 10284 28150
rect 10232 28086 10284 28092
rect 10428 28082 10456 29650
rect 10888 29510 10916 30126
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 10888 29238 10916 29446
rect 10876 29232 10928 29238
rect 10876 29174 10928 29180
rect 10508 28960 10560 28966
rect 10508 28902 10560 28908
rect 10520 28082 10548 28902
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 7564 27668 7616 27674
rect 7564 27610 7616 27616
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 8312 26586 8340 26862
rect 9404 26784 9456 26790
rect 9456 26732 9536 26738
rect 9404 26726 9536 26732
rect 9416 26710 9536 26726
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8116 26444 8168 26450
rect 8116 26386 8168 26392
rect 8128 25770 8156 26386
rect 9508 26382 9536 26710
rect 9692 26586 9720 26862
rect 10244 26790 10272 27406
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 10244 26450 10272 26726
rect 10232 26444 10284 26450
rect 10232 26386 10284 26392
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 9772 26376 9824 26382
rect 9772 26318 9824 26324
rect 10048 26376 10100 26382
rect 10048 26318 10100 26324
rect 8496 26042 8524 26318
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 8588 25974 8616 26318
rect 9508 26042 9536 26318
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 9600 26042 9628 26182
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 8576 25968 8628 25974
rect 8576 25910 8628 25916
rect 8852 25900 8904 25906
rect 8852 25842 8904 25848
rect 8392 25832 8444 25838
rect 8392 25774 8444 25780
rect 8116 25764 8168 25770
rect 8116 25706 8168 25712
rect 8128 25498 8156 25706
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 8024 24948 8076 24954
rect 8024 24890 8076 24896
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6564 24274 6592 24550
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6920 24200 6972 24206
rect 6840 24160 6920 24188
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6840 23322 6868 24160
rect 6920 24142 6972 24148
rect 7024 24138 7052 24686
rect 7300 24410 7328 24686
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7392 24290 7420 24346
rect 7300 24274 7420 24290
rect 7484 24274 7512 24550
rect 7668 24313 7696 24754
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7852 24410 7880 24686
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7654 24304 7710 24313
rect 7288 24268 7420 24274
rect 7340 24262 7420 24268
rect 7472 24268 7524 24274
rect 7288 24210 7340 24216
rect 7654 24239 7710 24248
rect 7472 24210 7524 24216
rect 7668 24206 7696 24239
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7024 23662 7052 24074
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6460 23248 6512 23254
rect 6460 23190 6512 23196
rect 6472 23118 6500 23190
rect 6840 23118 6868 23258
rect 5776 23060 5948 23066
rect 5724 23054 5948 23060
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 5736 23038 5948 23054
rect 5632 22976 5684 22982
rect 5552 22936 5632 22964
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5552 21486 5580 22936
rect 5632 22918 5684 22924
rect 5724 22976 5776 22982
rect 5724 22918 5776 22924
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5644 22030 5672 22714
rect 5736 22574 5764 22918
rect 5920 22642 5948 23038
rect 6184 23044 6236 23050
rect 6184 22986 6236 22992
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5724 22568 5776 22574
rect 5920 22522 5948 22578
rect 5724 22510 5776 22516
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3896 20330 3924 20878
rect 4816 20874 4844 21286
rect 4804 20868 4856 20874
rect 4804 20810 4856 20816
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4724 20398 4752 20742
rect 4816 20534 4844 20810
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5368 20602 5396 20810
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 4804 20528 4856 20534
rect 4856 20476 5028 20482
rect 4804 20470 5028 20476
rect 4816 20454 5028 20470
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 3884 20324 3936 20330
rect 3884 20266 3936 20272
rect 3700 20052 3752 20058
rect 3700 19994 3752 20000
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 3436 19378 3464 19654
rect 3528 19378 3556 19722
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 2872 18284 2924 18290
rect 2792 18244 2872 18272
rect 2872 18226 2924 18232
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1412 16658 1440 18158
rect 1780 17882 1808 18158
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 15026 1440 16594
rect 1676 16516 1728 16522
rect 1676 16458 1728 16464
rect 1688 16182 1716 16458
rect 1676 16176 1728 16182
rect 1676 16118 1728 16124
rect 2424 16114 2452 16934
rect 2516 16454 2544 17138
rect 2884 17082 2912 18226
rect 3252 18222 3280 18702
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3436 18154 3464 19314
rect 3528 18970 3556 19314
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3712 18766 3740 19994
rect 3896 19990 3924 20266
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 3896 19786 3924 19926
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3988 18970 4016 19790
rect 4080 19446 4108 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4724 19854 4752 20334
rect 5000 20262 5028 20454
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4712 19848 4764 19854
rect 4632 19796 4712 19802
rect 4632 19790 4764 19796
rect 4632 19774 4752 19790
rect 5000 19786 5028 20198
rect 4988 19780 5040 19786
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 4528 18896 4580 18902
rect 4448 18844 4528 18850
rect 4632 18850 4660 19774
rect 4988 19722 5040 19728
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 4580 18844 4660 18850
rect 4448 18822 4660 18844
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 2976 17678 3004 18090
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3160 17218 3188 17614
rect 3068 17190 3188 17218
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 2700 17066 3004 17082
rect 2700 17060 3016 17066
rect 2700 17054 2964 17060
rect 2700 16522 2728 17054
rect 2964 17002 3016 17008
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2872 16992 2924 16998
rect 3068 16946 3096 17190
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 2872 16934 2924 16940
rect 2688 16516 2740 16522
rect 2688 16458 2740 16464
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 16182 2544 16390
rect 2504 16176 2556 16182
rect 2504 16118 2556 16124
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2516 15706 2544 16118
rect 2700 15994 2728 16458
rect 2792 16114 2820 16934
rect 2884 16250 2912 16934
rect 2976 16918 3096 16946
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2976 16046 3004 16918
rect 3160 16794 3188 17070
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3160 16454 3188 16730
rect 3252 16522 3280 17206
rect 3804 17134 3832 18226
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3896 17270 3924 18158
rect 3988 18086 4016 18702
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 4080 17864 4108 18090
rect 4356 18086 4384 18702
rect 4448 18290 4476 18822
rect 4724 18766 4752 19654
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5276 19310 5304 19654
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4540 18426 4568 18702
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4080 17836 4200 17864
rect 4172 17678 4200 17836
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4448 17270 4476 17614
rect 4528 17604 4580 17610
rect 4528 17546 4580 17552
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 4080 16658 4108 17138
rect 4540 16998 4568 17546
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3240 16516 3292 16522
rect 3240 16458 3292 16464
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 2964 16040 3016 16046
rect 2700 15966 2820 15994
rect 2964 15982 3016 15988
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2516 15502 2544 15642
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 13938 1440 14962
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2424 14414 2452 15302
rect 2792 15026 2820 15966
rect 2976 15502 3004 15982
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2976 15026 3004 15438
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1872 13394 1900 14350
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 13546 2728 14214
rect 2792 14006 2820 14962
rect 3068 14414 3096 15438
rect 3160 15434 3188 16390
rect 3252 15910 3280 16458
rect 4080 16182 4108 16594
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16250 4200 16390
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15706 4660 18566
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4724 17882 4752 18294
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3252 14482 3280 14758
rect 3620 14482 3648 15098
rect 4080 14958 4108 15506
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2792 13870 2820 13942
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 3344 13734 3372 14214
rect 3620 14074 3648 14418
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3712 14006 3740 14758
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 2700 13530 2820 13546
rect 2700 13524 2832 13530
rect 2700 13518 2780 13524
rect 2780 13466 2832 13472
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2516 12782 2544 13194
rect 2792 12918 2820 13330
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2516 11286 2544 12718
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 1308 11144 1360 11150
rect 1308 11086 1360 11092
rect 1320 10985 1348 11086
rect 1584 11008 1636 11014
rect 1306 10976 1362 10985
rect 1584 10950 1636 10956
rect 1306 10911 1362 10920
rect 1596 10674 1624 10950
rect 2516 10674 2544 11222
rect 2884 10742 2912 11494
rect 2976 11218 3004 11698
rect 3436 11626 3464 12106
rect 3712 11762 3740 13942
rect 3896 13530 3924 14350
rect 4080 14346 4108 14894
rect 4264 14822 4292 15574
rect 4724 15178 4752 16934
rect 4540 15150 4752 15178
rect 4540 14958 4568 15150
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4632 14906 4660 15030
rect 4816 15008 4844 18566
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4908 17542 4936 18226
rect 5000 17882 5028 18226
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 5092 17814 5120 18022
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5080 17808 5132 17814
rect 5080 17750 5132 17756
rect 5092 17610 5120 17750
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17338 5304 17478
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5368 17134 5396 17818
rect 5460 17490 5488 21354
rect 5644 21010 5672 21966
rect 5736 21554 5764 22510
rect 5828 22494 5948 22522
rect 5828 21554 5856 22494
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5920 22234 5948 22374
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 6012 21418 6040 22578
rect 6196 21690 6224 22986
rect 6380 22094 6408 23054
rect 6656 22710 6684 23054
rect 6840 22778 6868 23054
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 7024 22710 7052 22918
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 7484 22574 7512 24074
rect 8036 22710 8064 24890
rect 8128 24886 8156 25434
rect 8404 25362 8432 25774
rect 8864 25430 8892 25842
rect 9220 25492 9272 25498
rect 9220 25434 9272 25440
rect 8852 25424 8904 25430
rect 8852 25366 8904 25372
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 9232 25294 9260 25434
rect 9508 25294 9536 25978
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 8116 24880 8168 24886
rect 8116 24822 8168 24828
rect 8496 24818 8524 25094
rect 9048 24886 9076 25162
rect 9036 24880 9088 24886
rect 9036 24822 9088 24828
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 24206 8156 24550
rect 8220 24274 8248 24754
rect 8772 24342 8800 24754
rect 8760 24336 8812 24342
rect 8760 24278 8812 24284
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8220 23866 8248 24210
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 8312 23866 8340 24074
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8404 22778 8432 23666
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8496 23118 8524 23462
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7484 22234 7512 22510
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 6380 22066 6500 22094
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6472 21554 6500 22066
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5552 20058 5580 20402
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5644 19922 5672 20946
rect 7944 20942 7972 21286
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7668 20398 7696 20878
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7760 20466 7788 20742
rect 8036 20534 8064 22646
rect 8496 22098 8524 23054
rect 8588 22982 8616 23802
rect 8772 23254 8800 24006
rect 9048 23866 9076 24074
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 8852 23792 8904 23798
rect 8852 23734 8904 23740
rect 8760 23248 8812 23254
rect 8760 23190 8812 23196
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8680 22710 8708 22918
rect 8772 22778 8800 23190
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8864 22166 8892 23734
rect 9048 23730 9076 23802
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 8956 23526 8984 23666
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8496 21010 8524 22034
rect 9048 22030 9076 23666
rect 9140 23594 9168 24754
rect 9232 24614 9260 25230
rect 9600 24970 9628 25978
rect 9784 25770 9812 26318
rect 9772 25764 9824 25770
rect 9772 25706 9824 25712
rect 10060 25702 10088 26318
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 10152 25838 10180 25910
rect 10140 25832 10192 25838
rect 10140 25774 10192 25780
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 9508 24954 9628 24970
rect 9508 24948 9640 24954
rect 9508 24942 9588 24948
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9324 24410 9352 24550
rect 9508 24410 9536 24942
rect 9588 24890 9640 24896
rect 9680 24812 9732 24818
rect 9600 24772 9680 24800
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 9232 23730 9260 24142
rect 9600 23866 9628 24772
rect 9680 24754 9732 24760
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9876 24274 9904 24618
rect 9864 24268 9916 24274
rect 9864 24210 9916 24216
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9600 23730 9628 23802
rect 9876 23746 9904 24210
rect 9784 23730 9904 23746
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9772 23724 9904 23730
rect 9824 23718 9904 23724
rect 9772 23666 9824 23672
rect 9128 23588 9180 23594
rect 9128 23530 9180 23536
rect 9232 23322 9260 23666
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9220 23044 9272 23050
rect 9220 22986 9272 22992
rect 9232 22778 9260 22986
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9600 22438 9628 23666
rect 10152 23662 10180 25774
rect 10244 24818 10272 26386
rect 10508 26308 10560 26314
rect 10508 26250 10560 26256
rect 10520 25838 10548 26250
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 11072 25158 11100 32846
rect 11336 32836 11388 32842
rect 11336 32778 11388 32784
rect 11152 32768 11204 32774
rect 11152 32710 11204 32716
rect 11164 31958 11192 32710
rect 11348 32230 11376 32778
rect 11808 32570 11836 33050
rect 12176 32842 12204 34002
rect 13096 33930 13124 34138
rect 13556 33998 13584 34546
rect 13648 34202 13676 34632
rect 13728 34614 13780 34620
rect 13636 34196 13688 34202
rect 13636 34138 13688 34144
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13924 33930 13952 34682
rect 14924 34672 14976 34678
rect 14476 34620 14924 34626
rect 14476 34614 14976 34620
rect 14476 34610 14964 34614
rect 14464 34604 14964 34610
rect 14516 34598 14964 34604
rect 14464 34546 14516 34552
rect 13084 33924 13136 33930
rect 13084 33866 13136 33872
rect 13912 33924 13964 33930
rect 13912 33866 13964 33872
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 12164 32836 12216 32842
rect 12164 32778 12216 32784
rect 13084 32836 13136 32842
rect 13084 32778 13136 32784
rect 13544 32836 13596 32842
rect 13544 32778 13596 32784
rect 13636 32836 13688 32842
rect 13636 32778 13688 32784
rect 11796 32564 11848 32570
rect 11796 32506 11848 32512
rect 12624 32564 12676 32570
rect 12624 32506 12676 32512
rect 11336 32224 11388 32230
rect 11336 32166 11388 32172
rect 11152 31952 11204 31958
rect 11152 31894 11204 31900
rect 11164 31278 11192 31894
rect 11348 31890 11376 32166
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 11808 31754 11836 32506
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12544 32026 12572 32302
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 11796 31748 11848 31754
rect 11796 31690 11848 31696
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 11716 31346 11744 31622
rect 12452 31482 12480 31758
rect 12440 31476 12492 31482
rect 12440 31418 12492 31424
rect 12636 31414 12664 32506
rect 12624 31408 12676 31414
rect 12624 31350 12676 31356
rect 13096 31346 13124 32778
rect 13556 32434 13584 32778
rect 13648 32502 13676 32778
rect 14200 32570 14228 32846
rect 14936 32842 14964 34598
rect 15028 34542 15056 34954
rect 15016 34536 15068 34542
rect 15016 34478 15068 34484
rect 15028 33998 15056 34478
rect 15304 34202 15332 34954
rect 15476 34944 15528 34950
rect 15476 34886 15528 34892
rect 15488 34678 15516 34886
rect 15672 34746 15700 35022
rect 16120 35012 16172 35018
rect 16120 34954 16172 34960
rect 16028 34944 16080 34950
rect 16028 34886 16080 34892
rect 15660 34740 15712 34746
rect 15660 34682 15712 34688
rect 15476 34672 15528 34678
rect 15476 34614 15528 34620
rect 16040 34610 16068 34886
rect 16132 34678 16160 34954
rect 16120 34672 16172 34678
rect 16120 34614 16172 34620
rect 16316 34610 16344 35158
rect 17052 34610 17080 35226
rect 17500 35080 17552 35086
rect 17500 35022 17552 35028
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 17408 35012 17460 35018
rect 17408 34954 17460 34960
rect 17420 34746 17448 34954
rect 17512 34950 17540 35022
rect 17500 34944 17552 34950
rect 17500 34886 17552 34892
rect 17868 34944 17920 34950
rect 17868 34886 17920 34892
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 16028 34604 16080 34610
rect 16028 34546 16080 34552
rect 16304 34604 16356 34610
rect 16304 34546 16356 34552
rect 17040 34604 17092 34610
rect 17040 34546 17092 34552
rect 15752 34536 15804 34542
rect 15752 34478 15804 34484
rect 15292 34196 15344 34202
rect 15292 34138 15344 34144
rect 15764 34066 15792 34478
rect 16212 34400 16264 34406
rect 16212 34342 16264 34348
rect 16224 34066 16252 34342
rect 15752 34060 15804 34066
rect 15672 34020 15752 34048
rect 15016 33992 15068 33998
rect 15016 33934 15068 33940
rect 15568 33516 15620 33522
rect 15568 33458 15620 33464
rect 15384 33312 15436 33318
rect 15384 33254 15436 33260
rect 14924 32836 14976 32842
rect 14924 32778 14976 32784
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14188 32564 14240 32570
rect 14188 32506 14240 32512
rect 14660 32502 14688 32710
rect 14936 32502 14964 32778
rect 13636 32496 13688 32502
rect 13636 32438 13688 32444
rect 14648 32496 14700 32502
rect 14648 32438 14700 32444
rect 14924 32496 14976 32502
rect 14924 32438 14976 32444
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14108 31482 14136 32370
rect 15396 32366 15424 33254
rect 15580 33046 15608 33458
rect 15568 33040 15620 33046
rect 15568 32982 15620 32988
rect 15672 32570 15700 34020
rect 15752 34002 15804 34008
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16316 33946 16344 34546
rect 16224 33918 16344 33946
rect 15936 33040 15988 33046
rect 15936 32982 15988 32988
rect 15660 32564 15712 32570
rect 15660 32506 15712 32512
rect 15384 32360 15436 32366
rect 15384 32302 15436 32308
rect 15396 32026 15424 32302
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15292 31884 15344 31890
rect 15292 31826 15344 31832
rect 15200 31816 15252 31822
rect 15200 31758 15252 31764
rect 14372 31680 14424 31686
rect 14372 31622 14424 31628
rect 14096 31476 14148 31482
rect 14096 31418 14148 31424
rect 13360 31408 13412 31414
rect 13360 31350 13412 31356
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 11796 31272 11848 31278
rect 11796 31214 11848 31220
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11164 30326 11192 30738
rect 11152 30320 11204 30326
rect 11152 30262 11204 30268
rect 11256 30122 11284 31078
rect 11808 30938 11836 31214
rect 11796 30932 11848 30938
rect 11796 30874 11848 30880
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11716 30258 11744 30534
rect 12360 30258 12388 31282
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 11244 30116 11296 30122
rect 11244 30058 11296 30064
rect 12636 30054 12664 30670
rect 13372 30326 13400 31350
rect 13912 31136 13964 31142
rect 13912 31078 13964 31084
rect 13636 30728 13688 30734
rect 13688 30676 13860 30682
rect 13636 30670 13860 30676
rect 13648 30654 13860 30670
rect 13924 30666 13952 31078
rect 14108 30938 14136 31418
rect 14384 31278 14412 31622
rect 15212 31482 15240 31758
rect 15304 31482 15332 31826
rect 15948 31754 15976 32982
rect 15936 31748 15988 31754
rect 15936 31690 15988 31696
rect 16120 31680 16172 31686
rect 16120 31622 16172 31628
rect 15200 31476 15252 31482
rect 15200 31418 15252 31424
rect 15292 31476 15344 31482
rect 15292 31418 15344 31424
rect 14372 31272 14424 31278
rect 14372 31214 14424 31220
rect 14096 30932 14148 30938
rect 14096 30874 14148 30880
rect 15212 30802 15240 31418
rect 16132 31414 16160 31622
rect 16224 31482 16252 33918
rect 17052 33862 17080 34546
rect 17420 34066 17448 34682
rect 17408 34060 17460 34066
rect 17408 34002 17460 34008
rect 17040 33856 17092 33862
rect 17040 33798 17092 33804
rect 16304 33448 16356 33454
rect 16304 33390 16356 33396
rect 16316 32910 16344 33390
rect 17040 33108 17092 33114
rect 17040 33050 17092 33056
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16316 32570 16344 32846
rect 16948 32768 17000 32774
rect 16948 32710 17000 32716
rect 16304 32564 16356 32570
rect 16304 32506 16356 32512
rect 16316 31754 16344 32506
rect 16960 32502 16988 32710
rect 16948 32496 17000 32502
rect 16948 32438 17000 32444
rect 16396 32360 16448 32366
rect 16396 32302 16448 32308
rect 16408 31754 16436 32302
rect 17052 32026 17080 33050
rect 17512 32910 17540 34886
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17604 33930 17632 34682
rect 17880 34542 17908 34886
rect 17868 34536 17920 34542
rect 17868 34478 17920 34484
rect 17880 33998 17908 34478
rect 18340 34202 18368 35022
rect 18880 34944 18932 34950
rect 18880 34886 18932 34892
rect 18892 34678 18920 34886
rect 18880 34672 18932 34678
rect 18880 34614 18932 34620
rect 19260 34542 19288 36110
rect 19444 35698 19472 36790
rect 19628 36582 19656 37062
rect 20824 36922 20852 37130
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20076 36848 20128 36854
rect 20076 36790 20128 36796
rect 19616 36576 19668 36582
rect 19616 36518 19668 36524
rect 20088 36378 20116 36790
rect 20076 36372 20128 36378
rect 20076 36314 20128 36320
rect 19524 36100 19576 36106
rect 19524 36042 19576 36048
rect 19984 36100 20036 36106
rect 19984 36042 20036 36048
rect 19536 35834 19564 36042
rect 19524 35828 19576 35834
rect 19524 35770 19576 35776
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19996 34746 20024 36042
rect 20088 35698 20116 36314
rect 20824 36174 20852 36858
rect 20812 36168 20864 36174
rect 21192 36156 21220 37130
rect 23860 37126 23888 39200
rect 24216 37256 24268 37262
rect 24216 37198 24268 37204
rect 25504 37256 25556 37262
rect 25504 37198 25556 37204
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 24228 36922 24256 37198
rect 21732 36916 21784 36922
rect 21732 36858 21784 36864
rect 24216 36916 24268 36922
rect 24216 36858 24268 36864
rect 21364 36712 21416 36718
rect 21364 36654 21416 36660
rect 21272 36168 21324 36174
rect 21192 36128 21272 36156
rect 20812 36110 20864 36116
rect 21272 36110 21324 36116
rect 20996 36032 21048 36038
rect 20996 35974 21048 35980
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 21008 35630 21036 35974
rect 20996 35624 21048 35630
rect 20996 35566 21048 35572
rect 21284 35562 21312 36110
rect 20444 35556 20496 35562
rect 20444 35498 20496 35504
rect 21272 35556 21324 35562
rect 21272 35498 21324 35504
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 19248 34536 19300 34542
rect 19248 34478 19300 34484
rect 18328 34196 18380 34202
rect 18328 34138 18380 34144
rect 19260 34066 19288 34478
rect 19248 34060 19300 34066
rect 19300 34020 19380 34048
rect 19248 34002 19300 34008
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 17592 33924 17644 33930
rect 17592 33866 17644 33872
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 18708 33318 18736 33458
rect 19352 33454 19380 34020
rect 19996 33930 20024 34682
rect 20352 34536 20404 34542
rect 20456 34524 20484 35498
rect 20536 35488 20588 35494
rect 20536 35430 20588 35436
rect 20548 35290 20576 35430
rect 20536 35284 20588 35290
rect 20536 35226 20588 35232
rect 21376 35018 21404 36654
rect 21744 36378 21772 36858
rect 23940 36848 23992 36854
rect 23940 36790 23992 36796
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22664 36378 22692 36654
rect 21732 36372 21784 36378
rect 21732 36314 21784 36320
rect 22652 36372 22704 36378
rect 22652 36314 22704 36320
rect 23664 36236 23716 36242
rect 23664 36178 23716 36184
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 22376 36168 22428 36174
rect 22376 36110 22428 36116
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 21468 35698 21496 35974
rect 21824 35760 21876 35766
rect 21824 35702 21876 35708
rect 21456 35692 21508 35698
rect 21456 35634 21508 35640
rect 21364 35012 21416 35018
rect 21364 34954 21416 34960
rect 20404 34496 20484 34524
rect 20352 34478 20404 34484
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 19524 33924 19576 33930
rect 19524 33866 19576 33872
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 19340 33448 19392 33454
rect 19340 33390 19392 33396
rect 18696 33312 18748 33318
rect 18696 33254 18748 33260
rect 18144 33108 18196 33114
rect 18144 33050 18196 33056
rect 18156 32910 18184 33050
rect 18708 32978 18736 33254
rect 18696 32972 18748 32978
rect 18696 32914 18748 32920
rect 19352 32910 19380 33390
rect 19536 33114 19564 33866
rect 19524 33108 19576 33114
rect 19524 33050 19576 33056
rect 17500 32904 17552 32910
rect 17500 32846 17552 32852
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 19340 32904 19392 32910
rect 19340 32846 19392 32852
rect 17512 32230 17540 32846
rect 17500 32224 17552 32230
rect 17500 32166 17552 32172
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 16304 31748 16356 31754
rect 16408 31726 16528 31754
rect 16304 31690 16356 31696
rect 16212 31476 16264 31482
rect 16264 31436 16436 31464
rect 16212 31418 16264 31424
rect 16120 31408 16172 31414
rect 16040 31356 16120 31362
rect 16040 31350 16172 31356
rect 16040 31334 16160 31350
rect 16212 31340 16264 31346
rect 15752 31136 15804 31142
rect 15752 31078 15804 31084
rect 14648 30796 14700 30802
rect 14648 30738 14700 30744
rect 15200 30796 15252 30802
rect 15200 30738 15252 30744
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 13360 30320 13412 30326
rect 13832 30308 13860 30654
rect 13912 30660 13964 30666
rect 13912 30602 13964 30608
rect 14004 30660 14056 30666
rect 14004 30602 14056 30608
rect 13912 30320 13964 30326
rect 13832 30280 13912 30308
rect 13360 30262 13412 30268
rect 13912 30262 13964 30268
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12636 29646 12664 29990
rect 13372 29850 13400 30262
rect 13360 29844 13412 29850
rect 13360 29786 13412 29792
rect 11152 29640 11204 29646
rect 12624 29640 12676 29646
rect 11204 29600 11284 29628
rect 11152 29582 11204 29588
rect 11256 29102 11284 29600
rect 12624 29582 12676 29588
rect 11520 29572 11572 29578
rect 11520 29514 11572 29520
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 11244 29096 11296 29102
rect 11244 29038 11296 29044
rect 11256 28762 11284 29038
rect 11244 28756 11296 28762
rect 11244 28698 11296 28704
rect 11440 28626 11468 29446
rect 11532 29306 11560 29514
rect 12636 29306 12664 29582
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 13372 29238 13400 29786
rect 13360 29232 13412 29238
rect 13360 29174 13412 29180
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11152 28552 11204 28558
rect 11152 28494 11204 28500
rect 11164 28082 11192 28494
rect 12636 28150 12664 29038
rect 12912 28762 12940 29106
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 13372 28558 13400 29174
rect 14016 29102 14044 30602
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14108 30258 14136 30534
rect 14568 30326 14596 30670
rect 14660 30394 14688 30738
rect 15764 30734 15792 31078
rect 16040 30938 16068 31334
rect 16212 31282 16264 31288
rect 16120 31272 16172 31278
rect 16120 31214 16172 31220
rect 16132 30938 16160 31214
rect 16028 30932 16080 30938
rect 16028 30874 16080 30880
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 15752 30728 15804 30734
rect 15752 30670 15804 30676
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14556 30320 14608 30326
rect 14556 30262 14608 30268
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14648 30184 14700 30190
rect 14648 30126 14700 30132
rect 14832 30184 14884 30190
rect 14832 30126 14884 30132
rect 14660 29850 14688 30126
rect 14648 29844 14700 29850
rect 14648 29786 14700 29792
rect 14844 29306 14872 30126
rect 15028 30122 15056 30670
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 15304 30190 15332 30602
rect 15752 30592 15804 30598
rect 15752 30534 15804 30540
rect 15292 30184 15344 30190
rect 15292 30126 15344 30132
rect 15016 30116 15068 30122
rect 15016 30058 15068 30064
rect 15028 29714 15056 30058
rect 15764 29714 15792 30534
rect 16040 30258 16068 30874
rect 16224 30870 16252 31282
rect 16408 31278 16436 31436
rect 16396 31272 16448 31278
rect 16396 31214 16448 31220
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16212 30864 16264 30870
rect 16212 30806 16264 30812
rect 16224 30394 16252 30806
rect 16316 30666 16344 30874
rect 16408 30666 16436 31214
rect 16500 30682 16528 31726
rect 17052 31482 17080 31962
rect 17696 31958 17724 32846
rect 17776 32768 17828 32774
rect 17776 32710 17828 32716
rect 17788 31958 17816 32710
rect 18156 32230 18184 32846
rect 18236 32768 18288 32774
rect 18236 32710 18288 32716
rect 18248 32434 18276 32710
rect 19352 32570 19380 32846
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 18512 32496 18564 32502
rect 18512 32438 18564 32444
rect 18880 32496 18932 32502
rect 18880 32438 18932 32444
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 18144 32224 18196 32230
rect 18144 32166 18196 32172
rect 17684 31952 17736 31958
rect 17604 31900 17684 31906
rect 17604 31894 17736 31900
rect 17776 31952 17828 31958
rect 17776 31894 17828 31900
rect 17500 31884 17552 31890
rect 17500 31826 17552 31832
rect 17604 31878 17724 31894
rect 17040 31476 17092 31482
rect 17040 31418 17092 31424
rect 16948 31340 17000 31346
rect 16948 31282 17000 31288
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16500 30666 16620 30682
rect 16304 30660 16356 30666
rect 16304 30602 16356 30608
rect 16396 30660 16448 30666
rect 16396 30602 16448 30608
rect 16500 30660 16632 30666
rect 16500 30654 16580 30660
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 15016 29708 15068 29714
rect 15016 29650 15068 29656
rect 15752 29708 15804 29714
rect 15752 29650 15804 29656
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 14004 29096 14056 29102
rect 14004 29038 14056 29044
rect 13544 28620 13596 28626
rect 13544 28562 13596 28568
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 13452 28484 13504 28490
rect 13452 28426 13504 28432
rect 12992 28416 13044 28422
rect 12992 28358 13044 28364
rect 12624 28144 12676 28150
rect 12624 28086 12676 28092
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 13004 28014 13032 28358
rect 12992 28008 13044 28014
rect 12992 27950 13044 27956
rect 13464 27418 13492 28426
rect 13556 27538 13584 28562
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 14188 28416 14240 28422
rect 14188 28358 14240 28364
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13544 27532 13596 27538
rect 13544 27474 13596 27480
rect 12624 27396 12676 27402
rect 13464 27390 13584 27418
rect 13648 27402 13676 28086
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 12624 27338 12676 27344
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11164 25702 11192 26862
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11532 26042 11560 26726
rect 12636 26314 12664 27338
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 11164 25498 11192 25638
rect 11152 25492 11204 25498
rect 11152 25434 11204 25440
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10244 24274 10272 24754
rect 10336 24750 10364 25094
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 10508 24608 10560 24614
rect 10508 24550 10560 24556
rect 10520 24274 10548 24550
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10244 23798 10272 24210
rect 10796 23798 10824 24754
rect 10232 23792 10284 23798
rect 10232 23734 10284 23740
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10244 23186 10272 23734
rect 11164 23730 11192 25162
rect 11808 24138 11836 26250
rect 13096 26246 13124 27270
rect 13464 27130 13492 27270
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13268 27056 13320 27062
rect 13268 26998 13320 27004
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 13188 26586 13216 26930
rect 13280 26586 13308 26998
rect 13452 26852 13504 26858
rect 13452 26794 13504 26800
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 11980 26240 12032 26246
rect 11980 26182 12032 26188
rect 13084 26240 13136 26246
rect 13084 26182 13136 26188
rect 11992 25906 12020 26182
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 12084 24818 12112 25230
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 12084 24410 12112 24754
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11164 23526 11192 23666
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 8944 21684 8996 21690
rect 9048 21672 9076 21966
rect 9692 21962 9720 22986
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 8996 21644 9076 21672
rect 8944 21626 8996 21632
rect 9692 21622 9720 21898
rect 9968 21622 9996 22034
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5736 19378 5764 20334
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6656 19922 6684 20198
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 6012 19242 6040 19722
rect 7484 19718 7512 20334
rect 7760 20058 7788 20402
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7932 19780 7984 19786
rect 8036 19768 8064 20470
rect 8496 20058 8524 20946
rect 8588 20602 8616 21422
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8588 19854 8616 20538
rect 9416 20534 9444 21082
rect 9692 21026 9720 21558
rect 10520 21486 10548 23122
rect 11808 22778 11836 24074
rect 12636 23662 12664 25094
rect 12728 24818 12756 25842
rect 13096 25838 13124 26182
rect 13188 26042 13216 26522
rect 13176 26036 13228 26042
rect 13176 25978 13228 25984
rect 13084 25832 13136 25838
rect 13280 25786 13308 26522
rect 13464 26382 13492 26794
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13084 25774 13136 25780
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11256 21962 11284 22034
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21690 11100 21830
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 10600 21480 10652 21486
rect 10600 21422 10652 21428
rect 10520 21162 10548 21422
rect 9600 20998 9720 21026
rect 10428 21134 10548 21162
rect 9600 20602 9628 20998
rect 10428 20942 10456 21134
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9692 20466 9720 20878
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 10612 19922 10640 21422
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10704 21010 10732 21286
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 11256 20874 11284 21898
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 7984 19740 8064 19768
rect 7932 19722 7984 19728
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7484 19378 7512 19654
rect 7944 19446 7972 19722
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6932 18834 6960 19110
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6564 17746 6592 18022
rect 6840 17746 6868 18634
rect 7484 18222 7512 19314
rect 8496 18970 8524 19314
rect 9784 19310 9812 19654
rect 10336 19310 10364 19654
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8024 18760 8076 18766
rect 8484 18760 8536 18766
rect 8076 18720 8156 18748
rect 8024 18702 8076 18708
rect 7564 18352 7616 18358
rect 7932 18352 7984 18358
rect 7616 18300 7696 18306
rect 7564 18294 7696 18300
rect 7932 18294 7984 18300
rect 7576 18278 7696 18294
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5460 17462 5580 17490
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5368 16726 5396 17070
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5080 16108 5132 16114
rect 5080 16050 5132 16056
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4908 15366 4936 15846
rect 5092 15638 5120 16050
rect 5276 15706 5304 16458
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5080 15632 5132 15638
rect 5080 15574 5132 15580
rect 5368 15570 5396 16662
rect 5460 16250 5488 17274
rect 5552 17082 5580 17462
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5552 17054 5672 17082
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5552 16114 5580 16934
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5644 15994 5672 17054
rect 5460 15966 5672 15994
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5080 15020 5132 15026
rect 4816 14980 5080 15008
rect 5080 14962 5132 14968
rect 4632 14878 4752 14906
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14550 4660 14758
rect 4724 14634 4752 14878
rect 4724 14618 4844 14634
rect 5276 14618 5304 15438
rect 5460 15178 5488 15966
rect 5460 15150 5580 15178
rect 5736 15162 5764 17138
rect 5920 17134 5948 17546
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5920 16522 5948 17070
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6380 16046 6408 16458
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6748 15994 6776 16934
rect 6840 16674 6868 17682
rect 7576 17678 7604 18022
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7024 16794 7052 17478
rect 7576 17134 7604 17614
rect 7668 17542 7696 18278
rect 7944 17746 7972 18294
rect 7932 17740 7984 17746
rect 7852 17700 7932 17728
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 17134 7696 17478
rect 7852 17338 7880 17700
rect 7932 17682 7984 17688
rect 8128 17542 8156 18720
rect 8484 18702 8536 18708
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 9128 18760 9180 18766
rect 9232 18748 9260 19246
rect 9180 18720 9260 18748
rect 9128 18702 9180 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18290 8340 18566
rect 8496 18426 8524 18702
rect 8680 18426 8708 18702
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8772 17882 8800 18226
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8128 17270 8156 17478
rect 9140 17270 9168 18158
rect 9232 17610 9260 18720
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9416 18426 9444 18634
rect 10336 18426 10364 19246
rect 10612 19224 10640 19858
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10784 19236 10836 19242
rect 10612 19196 10784 19224
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10428 17678 10456 18634
rect 10704 18222 10732 19196
rect 10784 19178 10836 19184
rect 10980 18902 11008 19246
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 18290 10916 18566
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9232 17270 9260 17546
rect 9324 17338 9352 17546
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 8116 17264 8168 17270
rect 8036 17212 8116 17218
rect 8036 17206 8168 17212
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 8036 17190 8156 17206
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6840 16658 6960 16674
rect 6840 16652 6972 16658
rect 6840 16646 6920 16652
rect 6840 16182 6868 16646
rect 6920 16594 6972 16600
rect 7576 16250 7604 17070
rect 8036 16522 8064 17190
rect 9232 16590 9260 17206
rect 10704 17134 10732 18158
rect 10888 17542 10916 18226
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10888 17338 10916 17478
rect 11164 17338 11192 17546
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11348 17218 11376 22578
rect 11704 22094 11756 22098
rect 11808 22094 11836 22714
rect 12084 22642 12112 22918
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 11704 22092 11836 22094
rect 11756 22066 11836 22092
rect 12532 22092 12584 22098
rect 11704 22034 11756 22040
rect 12532 22034 12584 22040
rect 11716 21894 11744 22034
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11808 21690 11836 21898
rect 12452 21690 12480 21898
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11624 20602 11652 21490
rect 12176 20942 12204 21558
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12176 20602 12204 20742
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12544 20466 12572 22034
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12728 20806 12756 21490
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12544 19922 12572 20402
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 11808 17610 11836 19722
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11900 19378 11928 19654
rect 12268 19378 12296 19722
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12452 19242 12480 19654
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12452 18766 12480 19178
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 11900 17882 11928 18158
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11256 17190 11376 17218
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 9692 16658 9720 17070
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16658 9812 16934
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 7932 16108 7984 16114
rect 8036 16096 8064 16458
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 16182 9168 16390
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 7984 16068 8064 16096
rect 7932 16050 7984 16056
rect 9232 16046 9260 16526
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9416 16250 9444 16390
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 6828 16040 6880 16046
rect 6748 15988 6828 15994
rect 6748 15982 6880 15988
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 6748 15966 6868 15982
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 4724 14612 4856 14618
rect 4724 14606 4804 14612
rect 4804 14554 4856 14560
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3988 13530 4016 14010
rect 4356 14006 4384 14350
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13716 4200 13806
rect 4080 13688 4200 13716
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4080 13410 4108 13688
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4080 13382 4200 13410
rect 4172 12918 4200 13382
rect 4620 13388 4672 13394
rect 4540 13348 4620 13376
rect 4540 13258 4568 13348
rect 4724 13376 4752 14486
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4816 13818 4844 14418
rect 5368 14346 5396 14894
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5368 14074 5396 14282
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5356 13932 5408 13938
rect 5460 13920 5488 15030
rect 5408 13892 5488 13920
rect 5356 13874 5408 13880
rect 4816 13790 4936 13818
rect 4908 13734 4936 13790
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4896 13728 4948 13734
rect 5264 13728 5316 13734
rect 4948 13688 5028 13716
rect 4896 13670 4948 13676
rect 4672 13348 4752 13376
rect 4620 13330 4672 13336
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4540 12986 4568 13194
rect 4632 12986 4660 13194
rect 4816 13190 4844 13670
rect 5000 13530 5028 13688
rect 5264 13670 5316 13676
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4816 12850 4844 13126
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4620 12844 4672 12850
rect 4804 12844 4856 12850
rect 4672 12804 4752 12832
rect 4620 12786 4672 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12434 4752 12804
rect 4804 12786 4856 12792
rect 5000 12782 5028 12922
rect 5276 12850 5304 13670
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 4988 12776 5040 12782
rect 5368 12730 5396 13874
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12918 5488 13126
rect 5552 12986 5580 15150
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5644 14006 5672 14962
rect 5736 14482 5764 15098
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5828 13734 5856 14758
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 4988 12718 5040 12724
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 5276 12702 5396 12730
rect 4540 12406 4752 12434
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 1320 10305 1348 10610
rect 1306 10296 1362 10305
rect 1306 10231 1308 10240
rect 1360 10231 1362 10240
rect 1308 10202 1360 10208
rect 940 9920 992 9926
rect 940 9862 992 9868
rect 952 9625 980 9862
rect 938 9616 994 9625
rect 938 9551 994 9560
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 7478 2912 8230
rect 3436 7818 3464 11562
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11218 3648 11494
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3896 11098 3924 12038
rect 4356 11694 4384 12174
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4448 11898 4476 12106
rect 4540 12102 4568 12406
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4540 11626 4568 12038
rect 4528 11620 4580 11626
rect 4528 11562 4580 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11354 4660 12038
rect 4724 11558 4752 12310
rect 4816 12306 4844 12650
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 5184 12238 5212 12378
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 3896 11082 4108 11098
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3896 11076 4120 11082
rect 3896 11070 4068 11076
rect 3712 10810 3740 11018
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3896 10674 3924 11070
rect 4068 11018 4120 11024
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3896 9926 3924 10610
rect 4172 10606 4200 11154
rect 4724 10606 4752 11494
rect 4816 11218 4844 11494
rect 5276 11286 5304 12702
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11354 5396 12038
rect 5460 11830 5488 12854
rect 5920 12850 5948 14350
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6196 14074 6224 14282
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6564 13938 6592 14962
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12918 6960 13126
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4816 10130 4844 10950
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5368 10674 5396 11290
rect 5828 11218 5856 12310
rect 6196 12238 6224 12786
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 11694 6224 12174
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 5920 11218 5948 11630
rect 6472 11354 6500 12106
rect 7024 11830 7052 15642
rect 9232 15502 9260 15982
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9232 15162 9260 15438
rect 9876 15162 9904 16390
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7484 14346 7512 15030
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 6564 10674 6592 11630
rect 7392 11218 7420 13262
rect 7484 12918 7512 14282
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 13938 7696 14214
rect 8312 14006 8340 15098
rect 10060 15094 10088 16118
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 8680 14550 8708 14894
rect 9600 14618 9628 14894
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 10060 14090 10088 15030
rect 10704 14958 10732 17070
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10888 15162 10916 15642
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 15162 11100 15370
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10520 14346 10548 14758
rect 10704 14482 10732 14894
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9968 14062 10180 14090
rect 9968 14006 9996 14062
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7484 12646 7512 12854
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7668 12306 7696 13126
rect 8312 12850 8340 13942
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8496 12714 8524 13262
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8036 12434 8064 12582
rect 8036 12406 8248 12434
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 11898 7788 12174
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7852 11286 7880 11630
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 8128 11218 8156 12242
rect 8220 12102 8248 12406
rect 8588 12238 8616 12582
rect 9140 12442 9168 13194
rect 9232 12782 9260 13398
rect 10060 13394 10088 13738
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10152 13258 10180 14062
rect 10244 13938 10272 14214
rect 10520 13938 10548 14282
rect 11072 14074 11100 14350
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11072 13938 11100 14010
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10244 13326 10272 13874
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9600 12986 9628 13126
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9692 12918 9720 13126
rect 10152 12918 10180 13194
rect 9680 12912 9732 12918
rect 10140 12912 10192 12918
rect 9680 12854 9732 12860
rect 10060 12872 10140 12900
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8220 11898 8248 12038
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8404 11830 8432 12038
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6564 10130 6592 10610
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9602 3924 9862
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 3804 9574 3924 9602
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 848 7336 900 7342
rect 848 7278 900 7284
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 860 6769 888 7278
rect 2608 6882 2636 7278
rect 2608 6866 2728 6882
rect 2608 6860 2740 6866
rect 2608 6854 2688 6860
rect 846 6760 902 6769
rect 846 6695 902 6704
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1688 6254 1716 6666
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 2608 5778 2636 6854
rect 2688 6802 2740 6808
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 860 5409 888 5646
rect 846 5400 902 5409
rect 846 5335 902 5344
rect 2884 5234 2912 6190
rect 3160 5642 3188 6734
rect 3804 6730 3832 9574
rect 5276 9518 5304 9930
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4816 8566 4844 9454
rect 6564 8906 6592 10066
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 8220 9874 8248 10678
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8312 10062 8340 10610
rect 8404 10266 8432 11086
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10810 8524 10950
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8680 10470 8708 11086
rect 8864 10674 8892 12038
rect 9784 11898 9812 12174
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10060 11830 10088 12872
rect 10140 12854 10192 12860
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 12442 10180 12582
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10888 11898 10916 12310
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9048 10674 9076 11086
rect 10888 10810 10916 11834
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8588 10130 8616 10406
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8496 10010 8524 10066
rect 8680 10010 8708 10406
rect 8772 10266 8800 10542
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 10336 10062 10364 10474
rect 8496 9982 8708 10010
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 9042 6684 9318
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 5368 8498 5396 8570
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 3896 8090 3924 8434
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7410 4016 7754
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4080 7342 4108 7822
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3252 6254 3280 6666
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6322 3372 6598
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 2976 5370 3004 5510
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3712 5234 3740 5510
rect 3804 5370 3832 6666
rect 3988 6322 4016 6938
rect 4080 6934 4108 7278
rect 4448 7206 4476 7822
rect 4724 7546 4752 8434
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7818 5396 8230
rect 5460 7954 5488 8842
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 8294 6040 8434
rect 6748 8294 6776 9862
rect 6840 9586 6868 9862
rect 8220 9846 8340 9874
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6840 8090 6868 8502
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 6840 7886 6868 8026
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 7024 7750 7052 8774
rect 7208 8090 7236 9522
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8128 9178 8156 9454
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7300 7750 7328 8434
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 8090 7512 8298
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8090 7788 8230
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 8128 7954 8156 9114
rect 8312 8906 8340 9846
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 8090 8340 8502
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8496 7886 8524 9522
rect 8588 8906 8616 9982
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9178 9444 9454
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9692 8974 9720 9862
rect 9864 9648 9916 9654
rect 9784 9596 9864 9602
rect 9784 9590 9916 9596
rect 9784 9574 9904 9590
rect 10692 9580 10744 9586
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 9508 8566 9536 8910
rect 9784 8566 9812 9574
rect 10692 9522 10744 9528
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 8974 10548 9318
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 9496 8560 9548 8566
rect 9772 8560 9824 8566
rect 9548 8520 9772 8548
rect 9496 8502 9548 8508
rect 9772 8502 9824 8508
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 7886 8616 8366
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 7886 9168 8230
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8576 7880 8628 7886
rect 9128 7880 9180 7886
rect 8576 7822 8628 7828
rect 8864 7828 9128 7834
rect 8864 7822 9180 7828
rect 8864 7818 9168 7822
rect 8852 7812 9168 7818
rect 8904 7806 9168 7812
rect 8852 7754 8904 7760
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4816 7410 4844 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4172 6168 4200 6802
rect 4816 6254 4844 7142
rect 4908 7002 4936 7142
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 5276 6186 5304 7346
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6322 5580 6598
rect 7208 6458 7236 6938
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7576 6322 7604 7346
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 6458 7788 7142
rect 8588 6798 8616 7278
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7760 6322 7788 6394
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 4080 6140 4200 6168
rect 5264 6180 5316 6186
rect 4080 5794 4108 6140
rect 5264 6122 5316 6128
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4080 5766 4200 5794
rect 4724 5778 4752 6054
rect 5552 5914 5580 6258
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 848 5160 900 5166
rect 848 5102 900 5108
rect 860 5001 888 5102
rect 846 4992 902 5001
rect 846 4927 902 4936
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 848 4480 900 4486
rect 848 4422 900 4428
rect 860 4321 888 4422
rect 846 4312 902 4321
rect 846 4247 902 4256
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3528 3738 3556 4014
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 848 3664 900 3670
rect 846 3632 848 3641
rect 900 3632 902 3641
rect 846 3567 902 3576
rect 3804 3398 3832 4558
rect 3896 3738 3924 5646
rect 4172 5302 4200 5766
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 7576 5710 7604 6258
rect 7760 5778 7788 6258
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5644 5370 5672 5646
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4172 5012 4200 5238
rect 4080 4984 4200 5012
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 4080 4706 4108 4984
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3896 3534 3924 3674
rect 3988 3534 4016 4694
rect 4080 4690 4200 4706
rect 4068 4684 4200 4690
rect 4120 4678 4200 4684
rect 4068 4626 4120 4632
rect 4172 4282 4200 4678
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4264 4282 4292 4490
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3738 4660 4422
rect 4816 4214 4844 5238
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4816 3738 4844 4150
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 848 2984 900 2990
rect 846 2952 848 2961
rect 900 2952 902 2961
rect 846 2887 902 2896
rect 3988 2854 4016 3334
rect 4172 3126 4200 3538
rect 4632 3534 4660 3674
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4540 3194 4568 3334
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4816 3126 4844 3674
rect 5000 3466 5028 3878
rect 5368 3602 5396 4626
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5552 4078 5580 4558
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5644 4026 5672 5306
rect 5736 5166 5764 5510
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 6012 4826 6040 5646
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6104 4622 6132 5510
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6196 4622 6224 5170
rect 6564 5030 6592 5646
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 5552 3942 5580 4014
rect 5644 3998 5764 4026
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 3602 5672 3878
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 5368 2774 5396 3538
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5644 3194 5672 3402
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5736 3058 5764 3998
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5828 2922 5856 4082
rect 6012 3194 6040 4082
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6104 3466 6132 3674
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6380 3398 6408 4082
rect 6564 3942 6592 4966
rect 6840 4690 6868 4966
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6932 4554 6960 5306
rect 7116 5234 7144 5510
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7392 5234 7420 5306
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 7576 4146 7604 5646
rect 7852 4604 7880 6666
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6254 8064 6598
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8128 5710 8156 6258
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5914 8248 6054
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 7944 5234 7972 5646
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8220 5166 8248 5850
rect 8312 5386 8340 6122
rect 8588 5642 8616 6734
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9232 6458 9260 6666
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8772 6118 8800 6258
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 9140 5914 9168 6190
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9140 5710 9168 5850
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8312 5358 8432 5386
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8312 4826 8340 5170
rect 8404 5166 8432 5358
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 9048 4826 9076 5646
rect 9324 5642 9352 6122
rect 9600 5760 9628 7958
rect 9784 6730 9812 8502
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9876 8090 9904 8366
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9968 7954 9996 8910
rect 10520 8294 10548 8910
rect 10704 8838 10732 9522
rect 10888 9382 10916 9998
rect 10980 9722 11008 10542
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 8906 10916 9318
rect 10980 9178 11008 9658
rect 11072 9450 11100 10066
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9680 5772 9732 5778
rect 9416 5732 9680 5760
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 7932 4616 7984 4622
rect 7852 4576 7932 4604
rect 7932 4558 7984 4564
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 7116 3738 7144 4082
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7116 3534 7144 3674
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 7116 3058 7144 3470
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 3126 7236 3334
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 5368 2746 5488 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5460 2514 5488 2746
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1306 5304 2382
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 7116 800 7144 2790
rect 7300 2514 7328 3878
rect 7576 3670 7604 4082
rect 7852 3738 7880 4082
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7944 2990 7972 4558
rect 8496 3738 8524 4762
rect 9232 4690 9260 5578
rect 9416 5030 9444 5732
rect 9680 5714 9732 5720
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8588 4146 8616 4490
rect 8576 4140 8628 4146
rect 8628 4100 8708 4128
rect 8576 4082 8628 4088
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8312 3398 8340 3470
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8312 3194 8340 3334
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7944 2378 7972 2926
rect 8496 2514 8524 3674
rect 8680 3482 8708 4100
rect 9508 4010 9536 5170
rect 9600 5098 9628 5578
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 9692 4826 9720 5102
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9600 3670 9628 4558
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 8852 3528 8904 3534
rect 8680 3476 8852 3482
rect 8680 3470 8904 3476
rect 8680 3466 8892 3470
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8668 3460 8892 3466
rect 8720 3454 8892 3460
rect 8668 3402 8720 3408
rect 8588 2650 8616 3402
rect 9232 3126 9260 3538
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 8772 2990 8800 3062
rect 9600 2990 9628 3606
rect 9692 3534 9720 3946
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9784 3126 9812 6666
rect 9968 6458 9996 7890
rect 10520 7886 10548 8230
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10336 7546 10364 7754
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10152 6390 10180 7414
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10152 5914 10180 6326
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9876 5234 9904 5646
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10428 4282 10456 7414
rect 10520 7342 10548 7822
rect 11164 7546 11192 14554
rect 11256 12374 11284 17190
rect 11336 17060 11388 17066
rect 11336 17002 11388 17008
rect 11348 16590 11376 17002
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 14482 11376 16186
rect 11440 15094 11468 16390
rect 11808 15434 11836 17546
rect 11992 17338 12020 18022
rect 12544 17746 12572 18158
rect 12636 17882 12664 18226
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 12544 17202 12572 17682
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12728 16794 12756 17138
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12728 15434 12756 15506
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 11808 15162 11836 15370
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11440 14618 11468 15030
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 13938 12204 14418
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 11808 13258 11836 13874
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 12850 11468 13126
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 12268 12102 12296 15098
rect 12728 15026 12756 15370
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12360 14618 12388 14894
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12452 13818 12480 14962
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 13938 12664 14350
rect 12820 14346 12848 25230
rect 13004 24954 13032 25230
rect 12992 24948 13044 24954
rect 12992 24890 13044 24896
rect 13096 24818 13124 25774
rect 13188 25758 13308 25786
rect 13188 25498 13216 25758
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 13280 25294 13308 25638
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13464 24818 13492 26318
rect 13556 25702 13584 27390
rect 13636 27396 13688 27402
rect 13636 27338 13688 27344
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13740 26382 13768 26862
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13648 25770 13676 26182
rect 13832 25838 13860 27950
rect 13924 27878 13952 28358
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13924 27674 13952 27814
rect 13912 27668 13964 27674
rect 13912 27610 13964 27616
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14016 26246 14044 26930
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 14108 26450 14136 26726
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 14004 26240 14056 26246
rect 14004 26182 14056 26188
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 13636 25764 13688 25770
rect 13636 25706 13688 25712
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 13084 24812 13136 24818
rect 13004 24772 13084 24800
rect 13004 24206 13032 24772
rect 13084 24754 13136 24760
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13004 23594 13032 24142
rect 13464 23798 13492 24754
rect 13648 24206 13676 25706
rect 14108 25498 14136 25842
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13924 24410 13952 24754
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13924 23866 13952 24346
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 14200 23594 14228 28358
rect 14372 27668 14424 27674
rect 14372 27610 14424 27616
rect 14384 26994 14412 27610
rect 15120 27606 15148 29446
rect 15212 29034 15240 29582
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15212 28626 15240 28970
rect 16316 28626 16344 30602
rect 15200 28620 15252 28626
rect 15200 28562 15252 28568
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 16304 28620 16356 28626
rect 16304 28562 16356 28568
rect 15212 28150 15240 28562
rect 15476 28416 15528 28422
rect 15476 28358 15528 28364
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15844 28416 15896 28422
rect 15844 28358 15896 28364
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15200 28144 15252 28150
rect 15200 28086 15252 28092
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 15108 27600 15160 27606
rect 15108 27542 15160 27548
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14464 26784 14516 26790
rect 14464 26726 14516 26732
rect 14476 26382 14504 26726
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14372 25900 14424 25906
rect 14372 25842 14424 25848
rect 14292 24410 14320 25842
rect 14384 25226 14412 25842
rect 14476 25838 14504 26182
rect 14464 25832 14516 25838
rect 14464 25774 14516 25780
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14384 23730 14412 24346
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 12992 23588 13044 23594
rect 12992 23530 13044 23536
rect 14188 23588 14240 23594
rect 14188 23530 14240 23536
rect 14464 23588 14516 23594
rect 14464 23530 14516 23536
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 21622 13032 22374
rect 13740 22098 13768 22510
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 13372 21350 13400 21626
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13004 21026 13032 21286
rect 13464 21146 13492 21490
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13556 21146 13584 21422
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13004 21010 13124 21026
rect 13004 21004 13136 21010
rect 13004 20998 13084 21004
rect 13556 20992 13584 21082
rect 13084 20946 13136 20952
rect 13464 20964 13584 20992
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13360 20936 13412 20942
rect 13464 20924 13492 20964
rect 13412 20896 13492 20924
rect 13360 20878 13412 20884
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12912 19378 12940 20538
rect 13004 19446 13032 20878
rect 13648 20874 13676 21490
rect 13740 21146 13768 22034
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13728 20868 13780 20874
rect 13728 20810 13780 20816
rect 13740 20602 13768 20810
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 19922 13492 20198
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13188 18970 13216 19314
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13372 18902 13400 19110
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13372 18766 13400 18838
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13280 18290 13308 18566
rect 13372 18290 13400 18702
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13464 18154 13492 19246
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12912 17678 12940 17818
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12912 14074 12940 15438
rect 13004 15434 13032 18090
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17678 13584 18022
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 13096 17202 13124 17546
rect 13648 17338 13676 18702
rect 13832 18426 13860 21014
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13924 20058 13952 20334
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14108 19990 14136 21626
rect 14200 21554 14228 21966
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14200 21146 14228 21354
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14292 20058 14320 22170
rect 14476 22114 14504 23530
rect 14568 22778 14596 27542
rect 15304 27538 15332 28154
rect 15488 28014 15516 28358
rect 15764 28218 15792 28358
rect 15752 28212 15804 28218
rect 15752 28154 15804 28160
rect 15476 28008 15528 28014
rect 15476 27950 15528 27956
rect 15856 27577 15884 28358
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15842 27568 15898 27577
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 15660 27532 15712 27538
rect 15948 27538 15976 28018
rect 16040 28014 16068 28562
rect 16500 28234 16528 30654
rect 16580 30602 16632 30608
rect 16684 30190 16712 31078
rect 16960 30938 16988 31282
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 17052 30054 17080 31418
rect 17408 31136 17460 31142
rect 17408 31078 17460 31084
rect 17224 30864 17276 30870
rect 17224 30806 17276 30812
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 17236 29850 17264 30806
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17328 29850 17356 30534
rect 17420 30394 17448 31078
rect 17408 30388 17460 30394
rect 17408 30330 17460 30336
rect 17420 29850 17448 30330
rect 17224 29844 17276 29850
rect 17224 29786 17276 29792
rect 17316 29844 17368 29850
rect 17316 29786 17368 29792
rect 17408 29844 17460 29850
rect 17408 29786 17460 29792
rect 17236 29646 17264 29786
rect 17224 29640 17276 29646
rect 17224 29582 17276 29588
rect 17512 29578 17540 31826
rect 17604 31278 17632 31878
rect 17788 31770 17816 31894
rect 17696 31754 17816 31770
rect 17684 31748 17816 31754
rect 17736 31742 17816 31748
rect 17684 31690 17736 31696
rect 17684 31408 17736 31414
rect 17684 31350 17736 31356
rect 17592 31272 17644 31278
rect 17592 31214 17644 31220
rect 17696 30870 17724 31350
rect 17972 31346 18000 32166
rect 18156 31822 18184 32166
rect 18248 31958 18276 32370
rect 18524 32026 18552 32438
rect 18892 32026 18920 32438
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 18248 31822 18276 31894
rect 19168 31890 19196 32370
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 18144 31816 18196 31822
rect 18144 31758 18196 31764
rect 18236 31816 18288 31822
rect 18236 31758 18288 31764
rect 18248 31482 18276 31758
rect 18604 31680 18656 31686
rect 18604 31622 18656 31628
rect 18616 31482 18644 31622
rect 18236 31476 18288 31482
rect 18236 31418 18288 31424
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 17684 30864 17736 30870
rect 17684 30806 17736 30812
rect 18156 30734 18184 31282
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 17880 30394 17908 30602
rect 17868 30388 17920 30394
rect 17868 30330 17920 30336
rect 17500 29572 17552 29578
rect 17500 29514 17552 29520
rect 17880 29510 17908 30330
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 17868 29504 17920 29510
rect 17920 29452 18000 29458
rect 17868 29446 18000 29452
rect 17880 29430 18000 29446
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16408 28206 16528 28234
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 15842 27503 15898 27512
rect 15936 27532 15988 27538
rect 15660 27474 15712 27480
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14844 26926 14872 27270
rect 14832 26920 14884 26926
rect 14832 26862 14884 26868
rect 15212 26314 15240 27406
rect 15304 26994 15332 27474
rect 15672 26994 15700 27474
rect 15292 26988 15344 26994
rect 15476 26988 15528 26994
rect 15344 26948 15424 26976
rect 15292 26930 15344 26936
rect 15396 26518 15424 26948
rect 15476 26930 15528 26936
rect 15660 26988 15712 26994
rect 15712 26948 15792 26976
rect 15660 26930 15712 26936
rect 15488 26518 15516 26930
rect 15384 26512 15436 26518
rect 15384 26454 15436 26460
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 14740 26240 14792 26246
rect 14740 26182 14792 26188
rect 15292 26240 15344 26246
rect 15292 26182 15344 26188
rect 14752 25158 14780 26182
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14844 24886 14872 25434
rect 14936 25430 14964 25842
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 14924 25424 14976 25430
rect 14924 25366 14976 25372
rect 15212 24954 15240 25774
rect 15304 25362 15332 26182
rect 15396 25498 15424 26454
rect 15764 26450 15792 26948
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 15580 25514 15608 26386
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15672 25906 15700 26318
rect 15660 25900 15712 25906
rect 15660 25842 15712 25848
rect 15488 25498 15608 25514
rect 15672 25498 15700 25842
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15488 25492 15620 25498
rect 15488 25486 15568 25492
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14844 24206 14872 24822
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14752 23866 14780 24006
rect 14844 23866 14872 24142
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 15028 23594 15056 24074
rect 15120 23730 15148 24210
rect 15212 24070 15240 24754
rect 15396 24750 15424 25230
rect 15488 25226 15516 25486
rect 15568 25434 15620 25440
rect 15660 25492 15712 25498
rect 15660 25434 15712 25440
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15476 25220 15528 25226
rect 15476 25162 15528 25168
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 15580 24614 15608 25298
rect 15764 25294 15792 26386
rect 15856 26042 15884 27503
rect 15936 27474 15988 27480
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15752 25288 15804 25294
rect 15752 25230 15804 25236
rect 15764 25158 15792 25230
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15764 24970 15792 25094
rect 15672 24942 15792 24970
rect 15844 24948 15896 24954
rect 15672 24818 15700 24942
rect 15844 24890 15896 24896
rect 15856 24818 15884 24890
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15764 24682 15792 24754
rect 15752 24676 15804 24682
rect 15752 24618 15804 24624
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15580 24274 15608 24550
rect 15764 24410 15792 24618
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 15212 23798 15240 24006
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15016 23588 15068 23594
rect 15016 23530 15068 23536
rect 16040 23118 16068 27950
rect 16408 27674 16436 28206
rect 16488 28144 16540 28150
rect 16488 28086 16540 28092
rect 16396 27668 16448 27674
rect 16396 27610 16448 27616
rect 16408 27402 16436 27610
rect 16396 27396 16448 27402
rect 16396 27338 16448 27344
rect 16304 27328 16356 27334
rect 16500 27282 16528 28086
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27674 16896 27814
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16960 27538 16988 28494
rect 17972 28490 18000 29430
rect 18340 29238 18368 29718
rect 18800 29646 18828 30602
rect 19352 30258 19380 32506
rect 19996 31754 20024 33866
rect 20364 33862 20392 34342
rect 20352 33856 20404 33862
rect 20352 33798 20404 33804
rect 20364 32978 20392 33798
rect 20456 33046 20484 34496
rect 21376 33862 21404 34954
rect 21836 34746 21864 35702
rect 21916 35556 21968 35562
rect 21916 35498 21968 35504
rect 21928 34746 21956 35498
rect 22204 35306 22232 36110
rect 22284 36032 22336 36038
rect 22284 35974 22336 35980
rect 22296 35494 22324 35974
rect 22284 35488 22336 35494
rect 22284 35430 22336 35436
rect 22204 35290 22324 35306
rect 22192 35284 22324 35290
rect 22244 35278 22324 35284
rect 22192 35226 22244 35232
rect 22192 35148 22244 35154
rect 22192 35090 22244 35096
rect 21732 34740 21784 34746
rect 21732 34682 21784 34688
rect 21824 34740 21876 34746
rect 21824 34682 21876 34688
rect 21916 34740 21968 34746
rect 21916 34682 21968 34688
rect 21744 34066 21772 34682
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 21824 34468 21876 34474
rect 21824 34410 21876 34416
rect 21732 34060 21784 34066
rect 21732 34002 21784 34008
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 21364 33856 21416 33862
rect 21364 33798 21416 33804
rect 21192 33658 21220 33798
rect 21180 33652 21232 33658
rect 21180 33594 21232 33600
rect 21272 33516 21324 33522
rect 21376 33504 21404 33798
rect 21836 33590 21864 34410
rect 22112 34406 22140 34478
rect 22100 34400 22152 34406
rect 22100 34342 22152 34348
rect 22204 34066 22232 35090
rect 22296 34610 22324 35278
rect 22388 35086 22416 36110
rect 23676 35698 23704 36178
rect 23756 36168 23808 36174
rect 23754 36136 23756 36145
rect 23808 36136 23810 36145
rect 23754 36071 23810 36080
rect 23768 35834 23796 36071
rect 23756 35828 23808 35834
rect 23756 35770 23808 35776
rect 23664 35692 23716 35698
rect 23664 35634 23716 35640
rect 23848 35692 23900 35698
rect 23848 35634 23900 35640
rect 23676 35086 23704 35634
rect 23860 35086 23888 35634
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 23296 35080 23348 35086
rect 23296 35022 23348 35028
rect 23664 35080 23716 35086
rect 23664 35022 23716 35028
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 22928 34944 22980 34950
rect 22928 34886 22980 34892
rect 22940 34746 22968 34886
rect 22928 34740 22980 34746
rect 22928 34682 22980 34688
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22468 34536 22520 34542
rect 22468 34478 22520 34484
rect 22192 34060 22244 34066
rect 22192 34002 22244 34008
rect 21916 33856 21968 33862
rect 21916 33798 21968 33804
rect 21824 33584 21876 33590
rect 21824 33526 21876 33532
rect 21324 33476 21404 33504
rect 21272 33458 21324 33464
rect 20444 33040 20496 33046
rect 20444 32982 20496 32988
rect 20352 32972 20404 32978
rect 20352 32914 20404 32920
rect 21928 32502 21956 33798
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 22020 32774 22048 33254
rect 22204 32910 22232 34002
rect 22284 33924 22336 33930
rect 22284 33866 22336 33872
rect 22296 33114 22324 33866
rect 22480 33658 22508 34478
rect 22848 34406 22876 34546
rect 23020 34468 23072 34474
rect 23020 34410 23072 34416
rect 22836 34400 22888 34406
rect 22836 34342 22888 34348
rect 22468 33652 22520 33658
rect 22468 33594 22520 33600
rect 22480 33522 22508 33594
rect 22468 33516 22520 33522
rect 22468 33458 22520 33464
rect 22848 33386 22876 34342
rect 23032 33522 23060 34410
rect 23204 34060 23256 34066
rect 23204 34002 23256 34008
rect 23216 33590 23244 34002
rect 23204 33584 23256 33590
rect 23204 33526 23256 33532
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 22836 33380 22888 33386
rect 22836 33322 22888 33328
rect 23308 33318 23336 35022
rect 23860 34542 23888 35022
rect 23952 34678 23980 36790
rect 24400 36780 24452 36786
rect 24400 36722 24452 36728
rect 24124 36576 24176 36582
rect 24124 36518 24176 36524
rect 24136 36174 24164 36518
rect 24412 36378 24440 36722
rect 24860 36712 24912 36718
rect 24860 36654 24912 36660
rect 25136 36712 25188 36718
rect 25136 36654 25188 36660
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 24124 36168 24176 36174
rect 24124 36110 24176 36116
rect 24216 36168 24268 36174
rect 24216 36110 24268 36116
rect 24032 35760 24084 35766
rect 24032 35702 24084 35708
rect 24044 35222 24072 35702
rect 24228 35494 24256 36110
rect 24780 35834 24808 36178
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 24780 35698 24808 35770
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 24216 35488 24268 35494
rect 24216 35430 24268 35436
rect 24308 35488 24360 35494
rect 24308 35430 24360 35436
rect 24032 35216 24084 35222
rect 24032 35158 24084 35164
rect 24228 35154 24256 35430
rect 24320 35290 24348 35430
rect 24308 35284 24360 35290
rect 24308 35226 24360 35232
rect 24216 35148 24268 35154
rect 24216 35090 24268 35096
rect 23940 34672 23992 34678
rect 23940 34614 23992 34620
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23676 33658 23704 33798
rect 23952 33658 23980 34614
rect 23664 33652 23716 33658
rect 23664 33594 23716 33600
rect 23940 33652 23992 33658
rect 23940 33594 23992 33600
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 23492 33386 23520 33458
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 23308 33046 23336 33254
rect 23296 33040 23348 33046
rect 23296 32982 23348 32988
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21916 32496 21968 32502
rect 21916 32438 21968 32444
rect 20720 32224 20772 32230
rect 20720 32166 20772 32172
rect 20732 31890 20760 32166
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 19984 31748 20036 31754
rect 19984 31690 20036 31696
rect 19996 31482 20024 31690
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 19996 30258 20024 31418
rect 20088 31414 20116 31826
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 20076 31408 20128 31414
rect 20076 31350 20128 31356
rect 21008 31346 21036 31758
rect 21928 31346 21956 32438
rect 22100 32428 22152 32434
rect 22204 32416 22232 32846
rect 23952 32842 23980 33594
rect 23940 32836 23992 32842
rect 23940 32778 23992 32784
rect 24216 32836 24268 32842
rect 24216 32778 24268 32784
rect 23756 32564 23808 32570
rect 23756 32506 23808 32512
rect 23664 32496 23716 32502
rect 23664 32438 23716 32444
rect 22152 32388 22232 32416
rect 22100 32370 22152 32376
rect 22112 31754 22140 32370
rect 22376 32360 22428 32366
rect 22376 32302 22428 32308
rect 22388 31754 22416 32302
rect 23676 31890 23704 32438
rect 23664 31884 23716 31890
rect 23664 31826 23716 31832
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 22008 31748 22060 31754
rect 22008 31690 22060 31696
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 22296 31726 22416 31754
rect 22560 31748 22612 31754
rect 22020 31482 22048 31690
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 22008 31476 22060 31482
rect 22008 31418 22060 31424
rect 22204 31346 22232 31622
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21916 31340 21968 31346
rect 21916 31282 21968 31288
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 21008 30802 21036 31282
rect 21640 31204 21692 31210
rect 21640 31146 21692 31152
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 21364 30660 21416 30666
rect 21364 30602 21416 30608
rect 21376 30394 21404 30602
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 18788 29640 18840 29646
rect 18788 29582 18840 29588
rect 18328 29232 18380 29238
rect 18328 29174 18380 29180
rect 19168 29170 19196 29990
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19260 29306 19288 29582
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19352 29238 19380 30194
rect 19444 29850 19472 30194
rect 19432 29844 19484 29850
rect 19432 29786 19484 29792
rect 19892 29640 19944 29646
rect 19892 29582 19944 29588
rect 19708 29572 19760 29578
rect 19708 29514 19760 29520
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 19720 29170 19748 29514
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19708 29164 19760 29170
rect 19708 29106 19760 29112
rect 18144 29028 18196 29034
rect 18144 28970 18196 28976
rect 17592 28484 17644 28490
rect 17592 28426 17644 28432
rect 17960 28484 18012 28490
rect 17960 28426 18012 28432
rect 17604 28218 17632 28426
rect 17592 28212 17644 28218
rect 17592 28154 17644 28160
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 17592 27600 17644 27606
rect 17590 27568 17592 27577
rect 17644 27568 17646 27577
rect 16948 27532 17000 27538
rect 17590 27503 17646 27512
rect 16948 27474 17000 27480
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 16356 27276 16528 27282
rect 16304 27270 16528 27276
rect 16316 27254 16528 27270
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16224 26246 16252 26862
rect 16500 26450 16528 27254
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16500 26330 16528 26386
rect 16408 26302 16528 26330
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 16224 25906 16252 26182
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16224 24818 16252 25842
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16316 24954 16344 25230
rect 16408 25226 16436 26302
rect 16488 26240 16540 26246
rect 16488 26182 16540 26188
rect 16396 25220 16448 25226
rect 16396 25162 16448 25168
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16212 24812 16264 24818
rect 16132 24772 16212 24800
rect 16132 23526 16160 24772
rect 16212 24754 16264 24760
rect 16316 24342 16344 24890
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 16316 24206 16344 24278
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16408 24070 16436 25162
rect 16500 24206 16528 26182
rect 17328 25974 17356 26318
rect 17512 26246 17540 26318
rect 17500 26240 17552 26246
rect 17500 26182 17552 26188
rect 17316 25968 17368 25974
rect 17316 25910 17368 25916
rect 17696 25702 17724 27406
rect 17788 27130 17816 27610
rect 17972 27402 18000 28018
rect 18156 28014 18184 28970
rect 19064 28484 19116 28490
rect 19064 28426 19116 28432
rect 19076 28218 19104 28426
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18052 28008 18104 28014
rect 18052 27950 18104 27956
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 17960 27396 18012 27402
rect 17960 27338 18012 27344
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17788 25906 17816 27066
rect 17880 27062 17908 27270
rect 17868 27056 17920 27062
rect 17868 26998 17920 27004
rect 17880 25974 17908 26998
rect 17972 26994 18000 27338
rect 18064 26994 18092 27950
rect 18788 27668 18840 27674
rect 18788 27610 18840 27616
rect 18694 27568 18750 27577
rect 18694 27503 18750 27512
rect 18708 27402 18736 27503
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17972 26382 18000 26930
rect 18156 26382 18184 27270
rect 18432 27130 18460 27270
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18432 26382 18460 27066
rect 18800 26382 18828 27610
rect 18892 27402 18920 28018
rect 19352 27606 19380 28086
rect 19524 28076 19576 28082
rect 19524 28018 19576 28024
rect 19536 27674 19564 28018
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19340 27600 19392 27606
rect 19154 27568 19210 27577
rect 19064 27532 19116 27538
rect 19340 27542 19392 27548
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19154 27503 19210 27512
rect 19064 27474 19116 27480
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18880 27396 18932 27402
rect 18880 27338 18932 27344
rect 18880 26512 18932 26518
rect 18880 26454 18932 26460
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 17868 25968 17920 25974
rect 17868 25910 17920 25916
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17500 24336 17552 24342
rect 17500 24278 17552 24284
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16592 23662 16620 24006
rect 17512 23730 17540 24278
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 16132 22982 16160 23462
rect 16592 23050 16620 23598
rect 16868 23526 16896 23666
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 17696 23186 17724 25638
rect 17788 24818 17816 25842
rect 17972 25294 18000 25978
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18156 25430 18184 25842
rect 18340 25838 18368 26318
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18144 25424 18196 25430
rect 18064 25372 18144 25378
rect 18064 25366 18196 25372
rect 18064 25350 18184 25366
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 17788 24138 17816 24754
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17958 23896 18014 23905
rect 17958 23831 18014 23840
rect 17972 23798 18000 23831
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 18064 23526 18092 25350
rect 18248 25294 18276 25638
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18156 24954 18184 25230
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 18144 24200 18196 24206
rect 18248 24188 18276 25230
rect 18196 24160 18276 24188
rect 18144 24142 18196 24148
rect 18144 23656 18196 23662
rect 18340 23644 18368 25298
rect 18432 24750 18460 26318
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18696 26240 18748 26246
rect 18696 26182 18748 26188
rect 18512 25900 18564 25906
rect 18512 25842 18564 25848
rect 18524 25498 18552 25842
rect 18616 25770 18644 26182
rect 18708 25906 18736 26182
rect 18892 25906 18920 26454
rect 18984 26382 19012 27406
rect 19076 26518 19104 27474
rect 19064 26512 19116 26518
rect 19064 26454 19116 26460
rect 18972 26376 19024 26382
rect 18972 26318 19024 26324
rect 19076 26314 19104 26454
rect 19064 26308 19116 26314
rect 19064 26250 19116 26256
rect 19076 25906 19104 26250
rect 19168 26042 19196 27503
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19352 27062 19380 27406
rect 19444 27402 19472 27542
rect 19536 27470 19564 27610
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19536 27130 19564 27406
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19628 26994 19656 27814
rect 19708 27396 19760 27402
rect 19708 27338 19760 27344
rect 19616 26988 19668 26994
rect 19616 26930 19668 26936
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19156 26036 19208 26042
rect 19156 25978 19208 25984
rect 19536 25906 19564 26726
rect 19628 26382 19656 26930
rect 19720 26926 19748 27338
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 19812 26994 19840 27270
rect 19800 26988 19852 26994
rect 19800 26930 19852 26936
rect 19708 26920 19760 26926
rect 19708 26862 19760 26868
rect 19720 26586 19748 26862
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 19524 25900 19576 25906
rect 19524 25842 19576 25848
rect 18604 25764 18656 25770
rect 18604 25706 18656 25712
rect 18512 25492 18564 25498
rect 18512 25434 18564 25440
rect 18616 25294 18644 25706
rect 18604 25288 18656 25294
rect 18892 25242 18920 25842
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 18972 25696 19024 25702
rect 19260 25684 19288 25774
rect 19024 25656 19288 25684
rect 18972 25638 19024 25644
rect 18604 25230 18656 25236
rect 18708 25214 18920 25242
rect 18708 24936 18736 25214
rect 18892 25158 18920 25214
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18880 25152 18932 25158
rect 18880 25094 18932 25100
rect 18616 24908 18736 24936
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18418 24304 18474 24313
rect 18418 24239 18420 24248
rect 18472 24239 18474 24248
rect 18512 24268 18564 24274
rect 18420 24210 18472 24216
rect 18512 24210 18564 24216
rect 18418 24168 18474 24177
rect 18418 24103 18420 24112
rect 18472 24103 18474 24112
rect 18420 24074 18472 24080
rect 18524 23866 18552 24210
rect 18616 24070 18644 24908
rect 18800 24886 18828 25094
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 18984 24818 19012 25638
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18708 24154 18736 24754
rect 19076 24206 19104 24890
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19352 24410 19380 24686
rect 19147 24404 19199 24410
rect 19248 24404 19300 24410
rect 19199 24364 19248 24392
rect 19147 24346 19199 24352
rect 19248 24346 19300 24352
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19536 24342 19564 25842
rect 19904 25786 19932 29582
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20272 29306 20300 29514
rect 20364 29306 20392 30194
rect 20536 30048 20588 30054
rect 20536 29990 20588 29996
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20548 29646 20576 29990
rect 20536 29640 20588 29646
rect 20536 29582 20588 29588
rect 20824 29510 20852 29990
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20352 29300 20404 29306
rect 20352 29242 20404 29248
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 20732 28150 20760 29242
rect 20824 29238 20852 29446
rect 21100 29306 21128 30194
rect 21652 30190 21680 31146
rect 21732 30252 21784 30258
rect 21732 30194 21784 30200
rect 21640 30184 21692 30190
rect 21640 30126 21692 30132
rect 21088 29300 21140 29306
rect 21088 29242 21140 29248
rect 20812 29232 20864 29238
rect 20812 29174 20864 29180
rect 21652 29170 21680 30126
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21640 29164 21692 29170
rect 21640 29106 21692 29112
rect 20916 28218 20944 29106
rect 21192 29034 21220 29106
rect 21180 29028 21232 29034
rect 21180 28970 21232 28976
rect 21640 29028 21692 29034
rect 21640 28970 21692 28976
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 20904 28212 20956 28218
rect 20904 28154 20956 28160
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20732 28014 20760 28086
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 20720 28008 20772 28014
rect 20720 27950 20772 27956
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 21180 28008 21232 28014
rect 21180 27950 21232 27956
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 20088 26994 20116 27814
rect 20444 27464 20496 27470
rect 20444 27406 20496 27412
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 19812 25758 19932 25786
rect 19812 24410 19840 25758
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19904 25294 19932 25638
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19996 24954 20024 26386
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19800 24404 19852 24410
rect 19800 24346 19852 24352
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 19524 24336 19576 24342
rect 19154 24304 19210 24313
rect 19524 24278 19576 24284
rect 19154 24239 19210 24248
rect 19168 24206 19196 24239
rect 18880 24200 18932 24206
rect 18708 24148 18880 24154
rect 18708 24142 18932 24148
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19246 24168 19302 24177
rect 18708 24126 18920 24142
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18708 23798 18736 24126
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18696 23792 18748 23798
rect 18196 23616 18368 23644
rect 18616 23752 18696 23780
rect 18144 23598 18196 23604
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 18156 22982 18184 23598
rect 18616 23322 18644 23752
rect 18696 23734 18748 23740
rect 18892 23730 18920 24006
rect 19076 23798 19104 24142
rect 19064 23792 19116 23798
rect 19168 23780 19196 24142
rect 19246 24103 19248 24112
rect 19300 24103 19302 24112
rect 19248 24074 19300 24080
rect 19246 23896 19302 23905
rect 19246 23831 19248 23840
rect 19300 23831 19302 23840
rect 19248 23802 19300 23808
rect 19064 23734 19116 23740
rect 19159 23752 19196 23780
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14568 22234 14596 22714
rect 15764 22234 15792 22918
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 14476 22086 14688 22114
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14476 21146 14504 21422
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14016 19378 14044 19654
rect 14108 19530 14136 19926
rect 14108 19502 14228 19530
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14016 19242 14044 19314
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 14016 18834 14044 19178
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14108 18766 14136 19314
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13924 18306 13952 18702
rect 13832 18290 13952 18306
rect 13820 18284 13952 18290
rect 13872 18278 13952 18284
rect 13820 18226 13872 18232
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13740 17542 13768 18158
rect 13832 17882 13860 18226
rect 14200 18222 14228 19502
rect 14384 19446 14412 20198
rect 14660 19854 14688 22086
rect 15120 21690 15148 22170
rect 16132 22098 16160 22918
rect 18708 22506 18736 23462
rect 18800 23186 18828 23598
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18800 22710 18828 23122
rect 18892 23118 18920 23666
rect 19159 23644 19187 23752
rect 19260 23730 19380 23746
rect 19260 23724 19392 23730
rect 19260 23718 19340 23724
rect 19159 23616 19196 23644
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 19168 22642 19196 23616
rect 19260 22982 19288 23718
rect 19340 23666 19392 23672
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 19352 23118 19380 23530
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 19352 22438 19380 23054
rect 19628 22778 19656 23054
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 16684 21622 16712 21898
rect 17420 21690 17448 21966
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 17040 21480 17092 21486
rect 17092 21440 17172 21468
rect 17040 21422 17092 21428
rect 15212 21010 15240 21422
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15580 20942 15608 21286
rect 17144 21146 17172 21440
rect 15936 21140 15988 21146
rect 17132 21140 17184 21146
rect 15936 21082 15988 21088
rect 16776 21100 16988 21128
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15580 20806 15608 20878
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14660 18970 14688 19790
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19378 14780 19654
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 13740 16658 13768 17478
rect 13832 17338 13860 17682
rect 14016 17610 14044 18158
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 13096 15502 13124 16118
rect 13280 15706 13308 16526
rect 13832 16114 13860 16526
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13556 15502 13584 15846
rect 13648 15638 13676 15982
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13832 15502 13860 15846
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 13096 15094 13124 15438
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13648 14958 13676 15098
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13004 14550 13032 14894
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13648 14278 13676 14418
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12900 13932 12952 13938
rect 13360 13932 13412 13938
rect 12900 13874 12952 13880
rect 13280 13892 13360 13920
rect 12360 13790 12480 13818
rect 12360 13394 12388 13790
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13394 12480 13670
rect 12636 13394 12664 13874
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12918 12480 13126
rect 12544 12986 12572 13262
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12820 12850 12848 13194
rect 12912 12986 12940 13874
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13004 13530 13032 13806
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13004 13190 13032 13466
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13096 12442 13124 12786
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12820 12102 12848 12242
rect 13188 12238 13216 13670
rect 13280 13326 13308 13892
rect 13360 13874 13412 13880
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13372 13530 13400 13738
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13464 13394 13492 14214
rect 13648 13734 13676 14214
rect 13740 14074 13768 15438
rect 14292 15162 14320 18702
rect 14752 18290 14780 19314
rect 15488 19310 15516 20198
rect 15672 19922 15700 20334
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15028 18766 15056 19110
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 14924 18352 14976 18358
rect 14924 18294 14976 18300
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14568 17338 14596 18022
rect 14752 17746 14780 18226
rect 14936 17882 14964 18294
rect 15028 18222 15056 18702
rect 15212 18426 15240 18702
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 15212 17202 15240 18362
rect 15304 18358 15332 18566
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15028 16794 15056 17138
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15304 16250 15332 16526
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15570 14412 15846
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14752 15162 14780 16050
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14844 15570 14872 15982
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 13832 14414 13860 15098
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13924 14414 13952 14554
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 14186 14376 14242 14385
rect 14186 14311 14188 14320
rect 14240 14311 14242 14320
rect 14188 14282 14240 14288
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12442 13400 13262
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 11624 11558 11652 12038
rect 11900 11830 11928 12038
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11900 11150 11928 11766
rect 12820 11694 12848 12038
rect 13096 11898 13124 12038
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12636 11286 12664 11494
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12820 11218 12848 11630
rect 12912 11558 12940 11834
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 13188 11218 13216 12174
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11348 10470 11376 10678
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 9654 11284 9862
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11348 7818 11376 10406
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 11624 8974 11652 10066
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11900 9722 11928 9930
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 12636 9518 12664 10066
rect 12912 10062 12940 10406
rect 13188 10130 13216 11154
rect 13372 11150 13400 12378
rect 13464 12374 13492 12582
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13556 12102 13584 12786
rect 13740 12306 13768 13398
rect 14016 13326 14044 13670
rect 14752 13394 14780 14214
rect 14844 14006 14872 15030
rect 15120 14958 15148 15914
rect 15212 15910 15240 16050
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14832 14000 14884 14006
rect 14884 13960 14964 13988
rect 14832 13942 14884 13948
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 10674 13400 11086
rect 13648 10810 13676 12174
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13740 11762 13768 12038
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13832 11626 13860 13262
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 12238 14136 12718
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13924 11762 13952 12106
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 14108 11150 14136 11630
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13096 9654 13124 9862
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11624 8634 11652 8910
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 12820 8566 12848 9318
rect 13188 9042 13216 9862
rect 13372 9722 13400 10610
rect 13832 10266 13860 10610
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13464 8906 13492 9998
rect 14016 9994 14044 10610
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13556 9722 13584 9862
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 14016 9518 14044 9930
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14016 9042 14044 9454
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13464 8566 13492 8842
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 7954 11560 8230
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 6322 10548 6598
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10796 6186 10824 7142
rect 11072 6730 11100 7278
rect 11348 6798 11376 7346
rect 11532 6798 11560 7686
rect 11716 6798 11744 8366
rect 13464 6866 13492 8502
rect 14108 7954 14136 11086
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14384 10810 14412 11018
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14476 10266 14504 13194
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12434 14872 13126
rect 14936 12918 14964 13960
rect 15120 13326 15148 14894
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14844 12406 14964 12434
rect 14936 11218 14964 12406
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14936 10810 14964 11154
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14660 10062 14688 10610
rect 14936 10198 14964 10746
rect 14924 10192 14976 10198
rect 14976 10140 15056 10146
rect 14924 10134 15056 10140
rect 14936 10118 15056 10134
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14200 9518 14228 9998
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 8974 14228 9454
rect 14292 9450 14320 9590
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14292 8430 14320 9386
rect 14568 9178 14596 9998
rect 14660 9654 14688 9998
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14936 8974 14964 9454
rect 15028 9382 15056 10118
rect 15212 9450 15240 15846
rect 15396 15706 15424 15982
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15292 12436 15344 12442
rect 15396 12424 15424 15642
rect 15488 15502 15516 17614
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 16250 15608 16526
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15672 15978 15700 19858
rect 15856 18970 15884 20402
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15948 18834 15976 21082
rect 16672 21072 16724 21078
rect 16776 21060 16804 21100
rect 16724 21032 16804 21060
rect 16960 21060 16988 21100
rect 17132 21082 17184 21088
rect 17040 21072 17092 21078
rect 16960 21032 17040 21060
rect 16672 21014 16724 21020
rect 17040 21014 17092 21020
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16868 20890 16896 20946
rect 16868 20862 16988 20890
rect 16960 20806 16988 20862
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16408 19922 16436 20742
rect 16868 20602 16896 20742
rect 16856 20596 16908 20602
rect 17420 20584 17448 21626
rect 17960 21480 18012 21486
rect 18064 21468 18092 21830
rect 18708 21690 18736 21898
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 18144 21480 18196 21486
rect 18064 21440 18144 21468
rect 17960 21422 18012 21428
rect 18144 21422 18196 21428
rect 17972 21146 18000 21422
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17868 21004 17920 21010
rect 17972 20992 18000 21082
rect 17920 20964 18000 20992
rect 17868 20946 17920 20952
rect 17500 20596 17552 20602
rect 17420 20556 17500 20584
rect 16856 20538 16908 20544
rect 17500 20538 17552 20544
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16592 19378 16620 20402
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16684 19378 16712 19994
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 17882 15792 18566
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15948 17270 15976 18770
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16040 18086 16068 18702
rect 16132 18290 16160 19314
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16132 17542 16160 18226
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 15948 16998 15976 17206
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15752 16720 15804 16726
rect 15752 16662 15804 16668
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 15094 15516 15438
rect 15672 15366 15700 15914
rect 15764 15502 15792 16662
rect 16316 16590 16344 18634
rect 16776 18426 16804 18770
rect 17052 18698 17080 19110
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 17052 18290 17080 18634
rect 17144 18358 17172 18906
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 17610 16988 18022
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 17236 16794 17264 18226
rect 17328 18222 17356 20334
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17420 18970 17448 20198
rect 17512 19786 17540 20538
rect 17972 20534 18000 20964
rect 18156 20806 18184 21422
rect 19260 21010 19288 22034
rect 19904 21894 19932 24346
rect 19996 23730 20024 24754
rect 20088 24342 20116 25434
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 20088 24138 20116 24278
rect 20180 24206 20208 26726
rect 20456 26586 20484 27406
rect 21100 27402 21128 27950
rect 21192 27606 21220 27950
rect 21180 27600 21232 27606
rect 21180 27542 21232 27548
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 26926 20668 27270
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20996 26852 21048 26858
rect 20996 26794 21048 26800
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20364 25906 20392 26522
rect 20628 26240 20680 26246
rect 20628 26182 20680 26188
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20640 25906 20668 26182
rect 20824 26042 20852 26182
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20076 24132 20128 24138
rect 20076 24074 20128 24080
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 20088 23118 20116 23802
rect 20180 23798 20208 24142
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20272 23730 20300 24890
rect 20364 23866 20392 25842
rect 20824 25294 20852 25842
rect 20904 25764 20956 25770
rect 20904 25706 20956 25712
rect 20916 25294 20944 25706
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20444 24880 20496 24886
rect 20444 24822 20496 24828
rect 20456 24274 20484 24822
rect 20548 24818 20576 25230
rect 20720 25220 20772 25226
rect 20720 25162 20772 25168
rect 20732 24834 20760 25162
rect 20916 25129 20944 25230
rect 20902 25120 20958 25129
rect 20902 25055 20958 25064
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20640 24806 20760 24834
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 19996 22778 20024 23054
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 19996 22094 20024 22714
rect 20272 22642 20300 23666
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20456 22234 20484 23462
rect 20548 23322 20576 24754
rect 20640 23866 20668 24806
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20640 23526 20668 23802
rect 20824 23662 20852 24142
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 19996 22066 20116 22094
rect 20088 22030 20116 22066
rect 20640 22030 20668 23462
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20824 22098 20852 23122
rect 20916 22166 20944 24686
rect 21008 24290 21036 26794
rect 21100 24410 21128 27338
rect 21284 25974 21312 28018
rect 21560 27878 21588 28494
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21560 27538 21588 27814
rect 21548 27532 21600 27538
rect 21548 27474 21600 27480
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 21376 27130 21404 27270
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 21468 26994 21496 27406
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21560 26994 21588 27338
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 21548 26988 21600 26994
rect 21548 26930 21600 26936
rect 21272 25968 21324 25974
rect 21272 25910 21324 25916
rect 21284 25158 21312 25910
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21376 25430 21404 25638
rect 21468 25498 21496 26930
rect 21652 26874 21680 28970
rect 21560 26846 21680 26874
rect 21456 25492 21508 25498
rect 21456 25434 21508 25440
rect 21364 25424 21416 25430
rect 21364 25366 21416 25372
rect 21364 25285 21416 25291
rect 21364 25227 21416 25233
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21192 24585 21220 25094
rect 21270 24984 21326 24993
rect 21270 24919 21326 24928
rect 21284 24614 21312 24919
rect 21272 24608 21324 24614
rect 21178 24576 21234 24585
rect 21272 24550 21324 24556
rect 21178 24511 21234 24520
rect 21088 24404 21140 24410
rect 21284 24392 21312 24550
rect 21088 24346 21140 24352
rect 21192 24364 21312 24392
rect 21008 24262 21128 24290
rect 21100 23730 21128 24262
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 21100 23118 21128 23666
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 21008 22778 21036 22986
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21192 22438 21220 24364
rect 21376 24070 21404 25227
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21376 23730 21404 24006
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 20904 22160 20956 22166
rect 20904 22102 20956 22108
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 17972 20058 18000 20470
rect 18156 20330 18184 20742
rect 18248 20602 18276 20810
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18524 20466 18552 20742
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18616 19922 18644 20402
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18708 19854 18736 20742
rect 18800 20330 18828 20946
rect 19260 20534 19288 20946
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17420 18766 17448 18906
rect 17604 18834 17632 19790
rect 18892 19786 18920 20402
rect 19352 20262 19380 21082
rect 19524 20868 19576 20874
rect 19524 20810 19576 20816
rect 19536 20602 19564 20810
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 20088 20398 20116 21830
rect 20732 21622 20760 21898
rect 20916 21894 20944 22102
rect 21376 22030 21404 22646
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20916 21350 20944 21490
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20364 20534 20392 21286
rect 21008 21146 21036 21966
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21008 20874 21036 21082
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 21008 20466 21036 20810
rect 21192 20534 21220 21014
rect 21468 21010 21496 21898
rect 21560 21350 21588 26846
rect 21640 26512 21692 26518
rect 21640 26454 21692 26460
rect 21652 25974 21680 26454
rect 21640 25968 21692 25974
rect 21640 25910 21692 25916
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21652 25158 21680 25298
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21640 24336 21692 24342
rect 21640 24278 21692 24284
rect 21652 24070 21680 24278
rect 21640 24064 21692 24070
rect 21640 24006 21692 24012
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 21652 22030 21680 22102
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21652 21486 21680 21966
rect 21744 21690 21772 30194
rect 21836 28218 21864 31282
rect 22296 31278 22324 31726
rect 22560 31690 22612 31696
rect 22572 31346 22600 31690
rect 22836 31680 22888 31686
rect 22836 31622 22888 31628
rect 22848 31414 22876 31622
rect 22836 31408 22888 31414
rect 22836 31350 22888 31356
rect 22560 31340 22612 31346
rect 22560 31282 22612 31288
rect 22284 31272 22336 31278
rect 22284 31214 22336 31220
rect 22100 30864 22152 30870
rect 22100 30806 22152 30812
rect 22112 30326 22140 30806
rect 22296 30598 22324 31214
rect 23584 30938 23612 31758
rect 23572 30932 23624 30938
rect 23572 30874 23624 30880
rect 23768 30734 23796 32506
rect 23848 32360 23900 32366
rect 23848 32302 23900 32308
rect 23860 30734 23888 32302
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23848 30728 23900 30734
rect 23848 30670 23900 30676
rect 22744 30660 22796 30666
rect 22744 30602 22796 30608
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22652 30592 22704 30598
rect 22652 30534 22704 30540
rect 22100 30320 22152 30326
rect 22100 30262 22152 30268
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 21928 29238 21956 30194
rect 22100 30184 22152 30190
rect 22020 30132 22100 30138
rect 22020 30126 22152 30132
rect 22020 30110 22140 30126
rect 22560 30116 22612 30122
rect 21916 29232 21968 29238
rect 21916 29174 21968 29180
rect 21928 28762 21956 29174
rect 22020 29034 22048 30110
rect 22560 30058 22612 30064
rect 22572 29646 22600 30058
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22468 29572 22520 29578
rect 22468 29514 22520 29520
rect 22100 29096 22152 29102
rect 22100 29038 22152 29044
rect 22008 29028 22060 29034
rect 22008 28970 22060 28976
rect 21916 28756 21968 28762
rect 21916 28698 21968 28704
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 22020 28150 22048 28970
rect 22112 28642 22140 29038
rect 22480 29034 22508 29514
rect 22468 29028 22520 29034
rect 22468 28970 22520 28976
rect 22112 28614 22508 28642
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22008 28144 22060 28150
rect 22008 28086 22060 28092
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 21836 27130 21864 27406
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21836 25498 21864 26930
rect 22204 26926 22232 28018
rect 22388 27062 22416 28494
rect 22376 27056 22428 27062
rect 22376 26998 22428 27004
rect 22192 26920 22244 26926
rect 22112 26880 22192 26908
rect 22112 25702 22140 26880
rect 22192 26862 22244 26868
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22192 25832 22244 25838
rect 22192 25774 22244 25780
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 21824 25492 21876 25498
rect 21824 25434 21876 25440
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 21824 24948 21876 24954
rect 21824 24890 21876 24896
rect 21836 24818 21864 24890
rect 22020 24886 22048 25230
rect 22008 24880 22060 24886
rect 22008 24822 22060 24828
rect 22112 24818 22140 25638
rect 22204 24954 22232 25774
rect 22296 25294 22324 25842
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22296 24993 22324 25230
rect 22282 24984 22338 24993
rect 22192 24948 22244 24954
rect 22282 24919 22338 24928
rect 22192 24890 22244 24896
rect 22480 24834 22508 28614
rect 22572 28082 22600 29582
rect 22664 28558 22692 30534
rect 22756 29850 22784 30602
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23492 30258 23520 30534
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23848 30252 23900 30258
rect 23848 30194 23900 30200
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 23676 29782 23704 30126
rect 23664 29776 23716 29782
rect 23664 29718 23716 29724
rect 23860 29714 23888 30194
rect 24044 29850 24072 30194
rect 24136 30122 24164 30194
rect 24124 30116 24176 30122
rect 24124 30058 24176 30064
rect 24032 29844 24084 29850
rect 24032 29786 24084 29792
rect 23848 29708 23900 29714
rect 23848 29650 23900 29656
rect 24124 29640 24176 29646
rect 24124 29582 24176 29588
rect 23296 29572 23348 29578
rect 24032 29572 24084 29578
rect 23348 29532 23520 29560
rect 23296 29514 23348 29520
rect 23112 29504 23164 29510
rect 23112 29446 23164 29452
rect 23124 29238 23152 29446
rect 23492 29238 23520 29532
rect 24032 29514 24084 29520
rect 24044 29238 24072 29514
rect 23112 29232 23164 29238
rect 23112 29174 23164 29180
rect 23480 29232 23532 29238
rect 23480 29174 23532 29180
rect 24032 29232 24084 29238
rect 24032 29174 24084 29180
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23584 28626 23612 29106
rect 23572 28620 23624 28626
rect 23572 28562 23624 28568
rect 23940 28620 23992 28626
rect 23940 28562 23992 28568
rect 22652 28552 22704 28558
rect 22704 28500 22784 28506
rect 22652 28494 22784 28500
rect 22664 28478 22784 28494
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22572 25906 22600 28018
rect 22756 27334 22784 28478
rect 22928 28484 22980 28490
rect 22928 28426 22980 28432
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 22848 28082 22876 28358
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 22836 27668 22888 27674
rect 22940 27656 22968 28426
rect 23952 28218 23980 28562
rect 23940 28212 23992 28218
rect 23940 28154 23992 28160
rect 22888 27628 22968 27656
rect 22836 27610 22888 27616
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 26994 22784 27270
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22664 25294 22692 25638
rect 22756 25362 22784 26930
rect 22848 25702 22876 27610
rect 24044 27470 24072 29174
rect 24136 29034 24164 29582
rect 24228 29322 24256 32778
rect 24320 32570 24348 35226
rect 24584 34944 24636 34950
rect 24584 34886 24636 34892
rect 24596 34678 24624 34886
rect 24584 34672 24636 34678
rect 24584 34614 24636 34620
rect 24872 34610 24900 36654
rect 25148 36378 25176 36654
rect 25136 36372 25188 36378
rect 25136 36314 25188 36320
rect 25044 36236 25096 36242
rect 25044 36178 25096 36184
rect 24952 35148 25004 35154
rect 25056 35136 25084 36178
rect 25228 36032 25280 36038
rect 25228 35974 25280 35980
rect 25240 35834 25268 35974
rect 25228 35828 25280 35834
rect 25228 35770 25280 35776
rect 25136 35692 25188 35698
rect 25136 35634 25188 35640
rect 25148 35494 25176 35634
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 25004 35108 25084 35136
rect 24952 35090 25004 35096
rect 24964 34678 24992 35090
rect 25228 34944 25280 34950
rect 25228 34886 25280 34892
rect 24952 34672 25004 34678
rect 24952 34614 25004 34620
rect 25240 34610 25268 34886
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 25228 34604 25280 34610
rect 25228 34546 25280 34552
rect 24872 34066 24900 34546
rect 25136 34536 25188 34542
rect 25136 34478 25188 34484
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24872 33522 24900 34002
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24308 32564 24360 32570
rect 24308 32506 24360 32512
rect 24676 32564 24728 32570
rect 24676 32506 24728 32512
rect 24688 32434 24716 32506
rect 25056 32434 25084 33798
rect 25148 32502 25176 34478
rect 25240 33862 25268 34546
rect 25516 34066 25544 37198
rect 25792 37126 25820 39200
rect 26436 37126 26464 39200
rect 27080 37262 27108 39200
rect 27724 37466 27752 39200
rect 27712 37460 27764 37466
rect 27712 37402 27764 37408
rect 28368 37262 28396 39200
rect 29012 37466 29040 39200
rect 29656 37466 29684 39200
rect 29000 37460 29052 37466
rect 29000 37402 29052 37408
rect 29644 37460 29696 37466
rect 29644 37402 29696 37408
rect 30300 37262 30328 39200
rect 30944 37262 30972 39200
rect 31588 37262 31616 39200
rect 32232 37262 32260 39200
rect 32876 37262 32904 39200
rect 33520 37262 33548 39200
rect 34164 37466 34192 39200
rect 34808 37466 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37466 35480 39200
rect 36096 37466 36124 39200
rect 36740 37466 36768 39200
rect 37922 38856 37978 38865
rect 37922 38791 37978 38800
rect 37936 37466 37964 38791
rect 38290 38176 38346 38185
rect 38290 38111 38346 38120
rect 38198 37496 38254 37505
rect 34152 37460 34204 37466
rect 34152 37402 34204 37408
rect 34796 37460 34848 37466
rect 34796 37402 34848 37408
rect 35440 37460 35492 37466
rect 35440 37402 35492 37408
rect 36084 37460 36136 37466
rect 36084 37402 36136 37408
rect 36728 37460 36780 37466
rect 36728 37402 36780 37408
rect 37924 37460 37976 37466
rect 38198 37431 38200 37440
rect 37924 37402 37976 37408
rect 38252 37431 38254 37440
rect 38200 37402 38252 37408
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 27068 37256 27120 37262
rect 27068 37198 27120 37204
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 30288 37256 30340 37262
rect 30288 37198 30340 37204
rect 30932 37256 30984 37262
rect 30932 37198 30984 37204
rect 31576 37256 31628 37262
rect 31576 37198 31628 37204
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 32864 37256 32916 37262
rect 32864 37198 32916 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 25780 37120 25832 37126
rect 25780 37062 25832 37068
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 26988 36922 27016 37198
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 26976 36916 27028 36922
rect 26976 36858 27028 36864
rect 30104 36916 30156 36922
rect 30104 36858 30156 36864
rect 27988 36848 28040 36854
rect 27988 36790 28040 36796
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 26608 36576 26660 36582
rect 26608 36518 26660 36524
rect 26620 36242 26648 36518
rect 27172 36378 27200 36722
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 27160 36372 27212 36378
rect 27160 36314 27212 36320
rect 27540 36258 27568 36654
rect 27620 36304 27672 36310
rect 27540 36252 27620 36258
rect 27540 36246 27672 36252
rect 26608 36236 26660 36242
rect 26608 36178 26660 36184
rect 27540 36230 27660 36246
rect 26148 36168 26200 36174
rect 26146 36136 26148 36145
rect 26200 36136 26202 36145
rect 26146 36071 26202 36080
rect 26160 35698 26188 36071
rect 26620 35698 26648 36178
rect 26976 36100 27028 36106
rect 26976 36042 27028 36048
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26608 35692 26660 35698
rect 26608 35634 26660 35640
rect 26240 35556 26292 35562
rect 26240 35498 26292 35504
rect 26148 35216 26200 35222
rect 26148 35158 26200 35164
rect 26160 34610 26188 35158
rect 26252 35154 26280 35498
rect 26240 35148 26292 35154
rect 26240 35090 26292 35096
rect 26988 35018 27016 36042
rect 27344 36032 27396 36038
rect 27344 35974 27396 35980
rect 27068 35488 27120 35494
rect 27120 35448 27200 35476
rect 27068 35430 27120 35436
rect 27172 35086 27200 35448
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 26976 35012 27028 35018
rect 26976 34954 27028 34960
rect 26148 34604 26200 34610
rect 26148 34546 26200 34552
rect 25504 34060 25556 34066
rect 25504 34002 25556 34008
rect 25228 33856 25280 33862
rect 25228 33798 25280 33804
rect 25516 33114 25544 34002
rect 27172 33522 27200 35022
rect 27264 34898 27292 35226
rect 27356 35018 27384 35974
rect 27540 35766 27568 36230
rect 27620 36100 27672 36106
rect 27620 36042 27672 36048
rect 27804 36100 27856 36106
rect 27804 36042 27856 36048
rect 27528 35760 27580 35766
rect 27528 35702 27580 35708
rect 27436 35488 27488 35494
rect 27436 35430 27488 35436
rect 27448 35290 27476 35430
rect 27436 35284 27488 35290
rect 27436 35226 27488 35232
rect 27344 35012 27396 35018
rect 27344 34954 27396 34960
rect 27436 34944 27488 34950
rect 27264 34892 27436 34898
rect 27264 34886 27488 34892
rect 27264 34870 27476 34886
rect 27356 33522 27384 34870
rect 27436 34060 27488 34066
rect 27540 34048 27568 35702
rect 27632 35630 27660 36042
rect 27620 35624 27672 35630
rect 27620 35566 27672 35572
rect 27632 35086 27660 35566
rect 27816 35154 27844 36042
rect 28000 35766 28028 36790
rect 28356 36712 28408 36718
rect 28356 36654 28408 36660
rect 29368 36712 29420 36718
rect 29368 36654 29420 36660
rect 28368 36378 28396 36654
rect 29380 36378 29408 36654
rect 29460 36576 29512 36582
rect 29460 36518 29512 36524
rect 28356 36372 28408 36378
rect 28356 36314 28408 36320
rect 29276 36372 29328 36378
rect 29276 36314 29328 36320
rect 29368 36372 29420 36378
rect 29368 36314 29420 36320
rect 28172 36100 28224 36106
rect 28172 36042 28224 36048
rect 29000 36100 29052 36106
rect 29000 36042 29052 36048
rect 27988 35760 28040 35766
rect 27988 35702 28040 35708
rect 27804 35148 27856 35154
rect 27804 35090 27856 35096
rect 27620 35080 27672 35086
rect 27620 35022 27672 35028
rect 27896 34468 27948 34474
rect 27896 34410 27948 34416
rect 27488 34020 27568 34048
rect 27436 34002 27488 34008
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 27344 33516 27396 33522
rect 27344 33458 27396 33464
rect 26240 33380 26292 33386
rect 26240 33322 26292 33328
rect 26252 33114 26280 33322
rect 26516 33312 26568 33318
rect 26516 33254 26568 33260
rect 26608 33312 26660 33318
rect 26608 33254 26660 33260
rect 27068 33312 27120 33318
rect 27068 33254 27120 33260
rect 25504 33108 25556 33114
rect 25504 33050 25556 33056
rect 26240 33108 26292 33114
rect 26240 33050 26292 33056
rect 25596 32836 25648 32842
rect 25596 32778 25648 32784
rect 25964 32836 26016 32842
rect 25964 32778 26016 32784
rect 25608 32570 25636 32778
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 25976 32434 26004 32778
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 25044 32428 25096 32434
rect 25044 32370 25096 32376
rect 25228 32428 25280 32434
rect 25228 32370 25280 32376
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25964 32428 26016 32434
rect 25964 32370 26016 32376
rect 26424 32428 26476 32434
rect 26424 32370 26476 32376
rect 24492 32224 24544 32230
rect 24492 32166 24544 32172
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24412 30802 24440 31622
rect 24504 31346 24532 32166
rect 24768 31952 24820 31958
rect 24768 31894 24820 31900
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 24400 30796 24452 30802
rect 24400 30738 24452 30744
rect 24504 30666 24532 31282
rect 24492 30660 24544 30666
rect 24492 30602 24544 30608
rect 24584 30660 24636 30666
rect 24584 30602 24636 30608
rect 24504 29578 24532 30602
rect 24596 30054 24624 30602
rect 24584 30048 24636 30054
rect 24584 29990 24636 29996
rect 24780 29782 24808 31894
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 24964 31482 24992 31758
rect 25056 31482 25084 31758
rect 24952 31476 25004 31482
rect 24952 31418 25004 31424
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 24860 31136 24912 31142
rect 24860 31078 24912 31084
rect 24872 30870 24900 31078
rect 24860 30864 24912 30870
rect 24860 30806 24912 30812
rect 25240 30802 25268 32370
rect 25332 32026 25360 32370
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25596 32020 25648 32026
rect 25596 31962 25648 31968
rect 25228 30796 25280 30802
rect 25228 30738 25280 30744
rect 25608 30734 25636 31962
rect 25976 30734 26004 32370
rect 26240 31408 26292 31414
rect 26240 31350 26292 31356
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 25228 30660 25280 30666
rect 25228 30602 25280 30608
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24872 30190 24900 30534
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 24952 30048 25004 30054
rect 24952 29990 25004 29996
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24584 29708 24636 29714
rect 24584 29650 24636 29656
rect 24492 29572 24544 29578
rect 24492 29514 24544 29520
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 24228 29306 24348 29322
rect 24228 29300 24360 29306
rect 24228 29294 24308 29300
rect 24124 29028 24176 29034
rect 24124 28970 24176 28976
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 22836 25696 22888 25702
rect 22836 25638 22888 25644
rect 22744 25356 22796 25362
rect 22744 25298 22796 25304
rect 22848 25294 22876 25638
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 22650 25120 22706 25129
rect 22650 25055 22706 25064
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 22100 24812 22152 24818
rect 22480 24806 22600 24834
rect 22664 24818 22692 25055
rect 22100 24754 22152 24760
rect 22008 24744 22060 24750
rect 21928 24692 22008 24698
rect 21928 24686 22060 24692
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 21928 24670 22048 24686
rect 21822 24576 21878 24585
rect 21822 24511 21878 24520
rect 21836 24206 21864 24511
rect 21928 24410 21956 24670
rect 22284 24608 22336 24614
rect 22284 24550 22336 24556
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21836 22030 21864 23666
rect 21928 23254 21956 24210
rect 22020 23866 22048 24278
rect 22296 24206 22324 24550
rect 22388 24342 22416 24550
rect 22376 24336 22428 24342
rect 22376 24278 22428 24284
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 22112 23594 22140 24074
rect 22480 24070 22508 24686
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22480 23730 22508 24006
rect 22572 23866 22600 24806
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 21916 23248 21968 23254
rect 21916 23190 21968 23196
rect 22112 22642 22140 23530
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21744 21146 21772 21490
rect 21836 21418 21864 21830
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21180 20528 21232 20534
rect 21180 20470 21232 20476
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19536 19854 19564 20198
rect 19812 20058 19840 20334
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17604 18426 17632 18634
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17696 18358 17724 19722
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18800 19446 18828 19654
rect 18788 19440 18840 19446
rect 18510 19408 18566 19417
rect 18788 19382 18840 19388
rect 18892 19378 18920 19722
rect 18510 19343 18512 19352
rect 18564 19343 18566 19352
rect 18696 19372 18748 19378
rect 18512 19314 18564 19320
rect 18696 19314 18748 19320
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17696 18154 17724 18294
rect 17788 18290 17816 18634
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17880 18358 17908 18566
rect 17868 18352 17920 18358
rect 17868 18294 17920 18300
rect 17972 18290 18000 19246
rect 18708 18902 18736 19314
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17972 17746 18000 18226
rect 18432 17882 18460 18702
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 18708 17678 18736 18838
rect 18892 18834 18920 19314
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19352 18834 19380 19110
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 15856 16182 15884 16526
rect 17972 16522 18000 17478
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15948 15552 15976 16390
rect 17314 16280 17370 16289
rect 17972 16266 18000 16458
rect 17972 16238 18184 16266
rect 17314 16215 17316 16224
rect 17368 16215 17370 16224
rect 17316 16186 17368 16192
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 16040 15706 16068 16050
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 16028 15564 16080 15570
rect 15948 15524 16028 15552
rect 16028 15506 16080 15512
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15488 13530 15516 13806
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15764 13394 15792 13806
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15764 12918 15792 13330
rect 16040 13326 16068 15506
rect 16224 15502 16252 15846
rect 16408 15638 16436 15982
rect 16684 15638 16712 16050
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16672 15632 16724 15638
rect 16672 15574 16724 15580
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16776 15434 16804 16050
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15672 12442 15700 12718
rect 15344 12396 15424 12424
rect 15660 12436 15712 12442
rect 15292 12378 15344 12384
rect 15660 12378 15712 12384
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 10606 15332 12174
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15304 9466 15332 9998
rect 15396 9722 15424 10066
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15200 9444 15252 9450
rect 15304 9438 15424 9466
rect 15200 9386 15252 9392
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14384 7954 14412 8230
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14476 7410 14504 8570
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10888 6322 10916 6394
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10704 5710 10732 6054
rect 10980 5778 11008 6054
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10520 5370 10548 5646
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 9968 3738 9996 3878
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 10520 2990 10548 3878
rect 10980 3670 11008 3878
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 11072 2854 11100 6666
rect 11532 6322 11560 6734
rect 11716 6458 11744 6734
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11808 6390 11836 6734
rect 12912 6730 12940 6802
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12084 6390 12112 6666
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11152 5840 11204 5846
rect 11256 5828 11284 6054
rect 11428 5908 11480 5914
rect 11204 5800 11284 5828
rect 11348 5868 11428 5896
rect 11152 5782 11204 5788
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11164 4826 11192 5646
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11256 5030 11284 5170
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11256 3670 11284 4966
rect 11348 4622 11376 5868
rect 11428 5850 11480 5856
rect 11888 5704 11940 5710
rect 11992 5692 12020 6054
rect 12176 5710 12204 6598
rect 12452 6186 12480 6666
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12268 5710 12296 6122
rect 12544 5710 12572 6326
rect 11940 5664 12020 5692
rect 11888 5646 11940 5652
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11440 4554 11468 5578
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5234 11928 5510
rect 11992 5302 12020 5664
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12728 5642 12756 6666
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6322 14136 6598
rect 12808 6316 12860 6322
rect 12992 6316 13044 6322
rect 12808 6258 12860 6264
rect 12912 6276 12992 6304
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12728 5522 12756 5578
rect 12544 5494 12756 5522
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12176 4690 12204 4966
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11440 4214 11468 4490
rect 12360 4282 12388 4966
rect 12544 4622 12572 5494
rect 12820 5234 12848 6258
rect 12912 5778 12940 6276
rect 12992 6258 13044 6264
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12912 5302 12940 5714
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13372 5574 13400 5646
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5370 13400 5510
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11532 3738 11560 4082
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 11900 3466 11928 4082
rect 12176 3534 12204 4150
rect 12360 4146 12388 4218
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12360 3466 12388 4082
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 3126 11836 3334
rect 12544 3126 12572 4558
rect 12636 4146 12664 4966
rect 13740 4554 13768 5102
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13648 4282 13676 4490
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13280 3194 13308 3470
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 14936 2650 14964 8910
rect 15028 8906 15056 9318
rect 15304 8974 15332 9318
rect 15396 9110 15424 9438
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15108 8832 15160 8838
rect 15488 8820 15516 11086
rect 16224 11082 16252 14350
rect 16592 13841 16620 14350
rect 16578 13832 16634 13841
rect 16578 13767 16634 13776
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16592 13394 16620 13670
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16592 11778 16620 12786
rect 16592 11750 16712 11778
rect 16684 11694 16712 11750
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11218 16712 11630
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 9722 16528 9998
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 15672 8838 15700 9522
rect 16408 9450 16436 9522
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16408 9178 16436 9386
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15108 8774 15160 8780
rect 15396 8792 15516 8820
rect 15568 8832 15620 8838
rect 15120 8566 15148 8774
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15396 7818 15424 8792
rect 15568 8774 15620 8780
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15580 8634 15608 8774
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15396 7698 15424 7754
rect 15212 7670 15424 7698
rect 15212 7478 15240 7670
rect 15672 7546 15700 8230
rect 15856 8090 15884 8910
rect 16408 8566 16436 9114
rect 16500 8838 16528 9522
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 16224 7954 16252 8366
rect 16408 7954 16436 8502
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7546 16436 7890
rect 16500 7750 16528 8774
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7546 16528 7686
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15212 6934 15240 7414
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 16592 6798 16620 11018
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16684 9654 16712 9862
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16776 9178 16804 15370
rect 16868 9926 16896 15574
rect 16960 14346 16988 15642
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 13938 17080 14214
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17144 12442 17172 15370
rect 17972 15026 18000 16050
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17958 14784 18014 14793
rect 17958 14719 18014 14728
rect 17776 14272 17828 14278
rect 17972 14226 18000 14719
rect 18064 14618 18092 15506
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18156 14346 18184 16238
rect 18248 16114 18276 16934
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18432 15706 18460 17138
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18616 16250 18644 16730
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 17776 14214 17828 14220
rect 17788 14074 17816 14214
rect 17880 14198 18000 14226
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 12918 17448 13670
rect 17604 13530 17632 13806
rect 17696 13530 17724 14010
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16960 11830 16988 12106
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17144 11354 17172 12378
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 11694 17540 12174
rect 17696 11898 17724 13194
rect 17880 12434 17908 14198
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17972 13870 18000 14010
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18156 13258 18184 14282
rect 18432 13326 18460 15642
rect 18708 15434 18736 16934
rect 18800 16794 18828 17206
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18800 16114 18828 16730
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18892 15994 18920 18770
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19444 17746 19472 18702
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18800 15966 18920 15994
rect 18696 15428 18748 15434
rect 18696 15370 18748 15376
rect 18800 15162 18828 15966
rect 18880 15496 18932 15502
rect 18984 15450 19012 17206
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 19076 15502 19104 16526
rect 18932 15444 19012 15450
rect 18880 15438 19012 15444
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 18892 15422 19012 15438
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18708 14278 18736 14962
rect 18892 14958 18920 15302
rect 18984 15026 19012 15422
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18892 14822 18920 14894
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18800 14482 18828 14758
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18892 14074 18920 14758
rect 19076 14414 19104 15438
rect 19168 15026 19196 16934
rect 19352 15978 19380 17546
rect 19444 16522 19472 17682
rect 19536 17134 19564 18294
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19628 17678 19656 18022
rect 19812 17882 19840 19246
rect 20088 18290 20116 20334
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20824 18766 20852 19382
rect 21284 19174 21312 20946
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21560 20398 21588 20470
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21468 19718 21496 19994
rect 21652 19922 21680 20266
rect 21744 20058 21772 21082
rect 21824 20936 21876 20942
rect 21928 20924 21956 21490
rect 22112 21486 22140 21898
rect 22100 21480 22152 21486
rect 22100 21422 22152 21428
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 21876 20896 21956 20924
rect 21824 20878 21876 20884
rect 21836 20210 21864 20878
rect 21914 20496 21970 20505
rect 21914 20431 21970 20440
rect 21928 20398 21956 20431
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21916 20256 21968 20262
rect 21836 20204 21916 20210
rect 21836 20198 21968 20204
rect 21836 20182 21956 20198
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21836 19854 21864 20182
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21456 19712 21508 19718
rect 21836 19666 21864 19790
rect 21456 19654 21508 19660
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18766 21312 19110
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 21284 18222 21312 18702
rect 21468 18698 21496 19654
rect 21744 19638 21864 19666
rect 21744 18766 21772 19638
rect 22020 19530 22048 21286
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 20380 22232 20742
rect 22296 20505 22324 22714
rect 22664 22506 22692 24754
rect 22848 24070 22876 25230
rect 22940 24750 22968 27406
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 23308 26994 23336 27270
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23584 26586 23612 26862
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 24136 26382 24164 28970
rect 24228 28626 24256 29294
rect 24308 29242 24360 29248
rect 24216 28620 24268 28626
rect 24216 28562 24268 28568
rect 24216 28484 24268 28490
rect 24216 28426 24268 28432
rect 24228 28150 24256 28426
rect 24216 28144 24268 28150
rect 24216 28086 24268 28092
rect 24228 26994 24256 28086
rect 24412 28082 24440 29446
rect 24596 28082 24624 29650
rect 24780 29578 24808 29718
rect 24768 29572 24820 29578
rect 24768 29514 24820 29520
rect 24676 29300 24728 29306
rect 24676 29242 24728 29248
rect 24688 28694 24716 29242
rect 24676 28688 24728 28694
rect 24676 28630 24728 28636
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24596 27538 24624 28018
rect 24780 28014 24808 29514
rect 24860 29504 24912 29510
rect 24860 29446 24912 29452
rect 24872 28082 24900 29446
rect 24964 28082 24992 29990
rect 25240 29646 25268 30602
rect 25424 30054 25452 30670
rect 26056 30660 26108 30666
rect 26056 30602 26108 30608
rect 26068 30190 26096 30602
rect 26252 30326 26280 31350
rect 26436 31278 26464 32370
rect 26424 31272 26476 31278
rect 26424 31214 26476 31220
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25964 30048 26016 30054
rect 25964 29990 26016 29996
rect 25976 29714 26004 29990
rect 26068 29782 26096 30126
rect 26056 29776 26108 29782
rect 26056 29718 26108 29724
rect 25964 29708 26016 29714
rect 25964 29650 26016 29656
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25228 29096 25280 29102
rect 25228 29038 25280 29044
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25240 28082 25268 29038
rect 25608 28490 25636 29038
rect 25792 29034 25820 29582
rect 26252 29578 26280 30262
rect 26240 29572 26292 29578
rect 26292 29532 26464 29560
rect 26240 29514 26292 29520
rect 26436 29306 26464 29532
rect 26528 29306 26556 33254
rect 26620 32978 26648 33254
rect 26608 32972 26660 32978
rect 26608 32914 26660 32920
rect 26620 31890 26648 32914
rect 26700 32768 26752 32774
rect 26700 32710 26752 32716
rect 26712 32570 26740 32710
rect 26700 32564 26752 32570
rect 26700 32506 26752 32512
rect 27080 32434 27108 33254
rect 27172 32910 27200 33458
rect 27356 33402 27384 33458
rect 27264 33374 27384 33402
rect 27264 32910 27292 33374
rect 27448 33046 27476 34002
rect 27712 33924 27764 33930
rect 27712 33866 27764 33872
rect 27724 33658 27752 33866
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 27908 33522 27936 34410
rect 28000 33930 28028 35702
rect 28184 35018 28212 36042
rect 28816 36032 28868 36038
rect 29012 35986 29040 36042
rect 28868 35980 29040 35986
rect 28816 35974 29040 35980
rect 29184 36032 29236 36038
rect 29184 35974 29236 35980
rect 28828 35958 29040 35974
rect 29012 35494 29040 35958
rect 29196 35834 29224 35974
rect 29184 35828 29236 35834
rect 29184 35770 29236 35776
rect 29000 35488 29052 35494
rect 29000 35430 29052 35436
rect 29288 35086 29316 36314
rect 29472 36174 29500 36518
rect 30116 36174 30144 36858
rect 31852 36848 31904 36854
rect 31852 36790 31904 36796
rect 31864 36174 31892 36790
rect 38304 36786 38332 38111
rect 38476 37120 38528 37126
rect 38476 37062 38528 37068
rect 38488 36825 38516 37062
rect 38474 36816 38530 36825
rect 38292 36780 38344 36786
rect 38580 36786 38608 39471
rect 38474 36751 38530 36760
rect 38568 36780 38620 36786
rect 38292 36722 38344 36728
rect 38568 36722 38620 36728
rect 33140 36712 33192 36718
rect 33140 36654 33192 36660
rect 29460 36168 29512 36174
rect 29460 36110 29512 36116
rect 30104 36168 30156 36174
rect 30104 36110 30156 36116
rect 31852 36168 31904 36174
rect 31852 36110 31904 36116
rect 29472 35766 29500 36110
rect 29460 35760 29512 35766
rect 29460 35702 29512 35708
rect 30116 35698 30144 36110
rect 30748 36100 30800 36106
rect 30748 36042 30800 36048
rect 30760 35834 30788 36042
rect 30748 35828 30800 35834
rect 30748 35770 30800 35776
rect 30472 35760 30524 35766
rect 30472 35702 30524 35708
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 30196 35556 30248 35562
rect 30196 35498 30248 35504
rect 30208 35222 30236 35498
rect 30484 35494 30512 35702
rect 30840 35624 30892 35630
rect 30840 35566 30892 35572
rect 31760 35624 31812 35630
rect 31760 35566 31812 35572
rect 30472 35488 30524 35494
rect 30472 35430 30524 35436
rect 30852 35290 30880 35566
rect 30840 35284 30892 35290
rect 30840 35226 30892 35232
rect 31208 35284 31260 35290
rect 31208 35226 31260 35232
rect 30196 35216 30248 35222
rect 30196 35158 30248 35164
rect 30104 35148 30156 35154
rect 30104 35090 30156 35096
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 29736 35080 29788 35086
rect 29736 35022 29788 35028
rect 28172 35012 28224 35018
rect 28172 34954 28224 34960
rect 28724 35012 28776 35018
rect 28724 34954 28776 34960
rect 28736 34610 28764 34954
rect 29748 34746 29776 35022
rect 29920 35012 29972 35018
rect 29920 34954 29972 34960
rect 29736 34740 29788 34746
rect 29736 34682 29788 34688
rect 28724 34604 28776 34610
rect 29184 34604 29236 34610
rect 28776 34564 28948 34592
rect 28724 34546 28776 34552
rect 28448 34536 28500 34542
rect 28632 34536 28684 34542
rect 28448 34478 28500 34484
rect 28552 34496 28632 34524
rect 27988 33924 28040 33930
rect 27988 33866 28040 33872
rect 27896 33516 27948 33522
rect 27896 33458 27948 33464
rect 27908 33114 27936 33458
rect 28000 33318 28028 33866
rect 28080 33856 28132 33862
rect 28080 33798 28132 33804
rect 28092 33522 28120 33798
rect 28460 33658 28488 34478
rect 28448 33652 28500 33658
rect 28448 33594 28500 33600
rect 28080 33516 28132 33522
rect 28080 33458 28132 33464
rect 28264 33516 28316 33522
rect 28264 33458 28316 33464
rect 27988 33312 28040 33318
rect 27988 33254 28040 33260
rect 27896 33108 27948 33114
rect 27896 33050 27948 33056
rect 27436 33040 27488 33046
rect 27488 32988 27844 32994
rect 27436 32982 27844 32988
rect 27448 32978 27844 32982
rect 27448 32972 27856 32978
rect 27448 32966 27804 32972
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 27252 32904 27304 32910
rect 27252 32846 27304 32852
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 26700 32292 26752 32298
rect 26700 32234 26752 32240
rect 26608 31884 26660 31890
rect 26608 31826 26660 31832
rect 26712 31822 26740 32234
rect 27344 32224 27396 32230
rect 27344 32166 27396 32172
rect 27356 31890 27384 32166
rect 27344 31884 27396 31890
rect 27344 31826 27396 31832
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 27448 31754 27476 32966
rect 27804 32914 27856 32920
rect 27988 32768 28040 32774
rect 27988 32710 28040 32716
rect 27896 32564 27948 32570
rect 27896 32506 27948 32512
rect 27804 32428 27856 32434
rect 27804 32370 27856 32376
rect 27816 32026 27844 32370
rect 27804 32020 27856 32026
rect 27804 31962 27856 31968
rect 27620 31952 27672 31958
rect 27908 31906 27936 32506
rect 27620 31894 27672 31900
rect 27356 31726 27476 31754
rect 27356 31346 27384 31726
rect 27632 31414 27660 31894
rect 27816 31878 27936 31906
rect 28000 31890 28028 32710
rect 28092 32502 28120 33458
rect 28276 32842 28304 33458
rect 28448 33312 28500 33318
rect 28448 33254 28500 33260
rect 28356 33040 28408 33046
rect 28356 32982 28408 32988
rect 28264 32836 28316 32842
rect 28264 32778 28316 32784
rect 28172 32768 28224 32774
rect 28172 32710 28224 32716
rect 28080 32496 28132 32502
rect 28080 32438 28132 32444
rect 28184 32434 28212 32710
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 28080 32360 28132 32366
rect 28080 32302 28132 32308
rect 28092 32026 28120 32302
rect 28276 32230 28304 32778
rect 28264 32224 28316 32230
rect 28264 32166 28316 32172
rect 28080 32020 28132 32026
rect 28080 31962 28132 31968
rect 27988 31884 28040 31890
rect 27816 31822 27844 31878
rect 27988 31826 28040 31832
rect 28276 31822 28304 32166
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28276 31482 28304 31758
rect 28368 31686 28396 32982
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 28460 31498 28488 33254
rect 28552 33046 28580 34496
rect 28920 34524 28948 34564
rect 29184 34546 29236 34552
rect 29276 34604 29328 34610
rect 29276 34546 29328 34552
rect 29000 34536 29052 34542
rect 28920 34496 29000 34524
rect 28632 34478 28684 34484
rect 29000 34478 29052 34484
rect 29000 34400 29052 34406
rect 29000 34342 29052 34348
rect 29012 33590 29040 34342
rect 29196 34202 29224 34546
rect 29184 34196 29236 34202
rect 29184 34138 29236 34144
rect 29000 33584 29052 33590
rect 29000 33526 29052 33532
rect 29196 33522 29224 34138
rect 29288 33658 29316 34546
rect 29932 34542 29960 34954
rect 30116 34610 30144 35090
rect 30208 35086 30236 35158
rect 31220 35086 31248 35226
rect 30196 35080 30248 35086
rect 30196 35022 30248 35028
rect 30656 35080 30708 35086
rect 30656 35022 30708 35028
rect 31208 35080 31260 35086
rect 31208 35022 31260 35028
rect 30208 34678 30236 35022
rect 30380 34944 30432 34950
rect 30380 34886 30432 34892
rect 30196 34672 30248 34678
rect 30196 34614 30248 34620
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 30288 34604 30340 34610
rect 30392 34592 30420 34886
rect 30668 34610 30696 35022
rect 31024 34944 31076 34950
rect 31024 34886 31076 34892
rect 31036 34610 31064 34886
rect 30340 34564 30420 34592
rect 30288 34546 30340 34552
rect 29920 34536 29972 34542
rect 29920 34478 29972 34484
rect 30392 34066 30420 34564
rect 30656 34604 30708 34610
rect 30656 34546 30708 34552
rect 31024 34604 31076 34610
rect 31024 34546 31076 34552
rect 30668 34474 30696 34546
rect 30472 34468 30524 34474
rect 30472 34410 30524 34416
rect 30656 34468 30708 34474
rect 30656 34410 30708 34416
rect 30380 34060 30432 34066
rect 30380 34002 30432 34008
rect 30484 33998 30512 34410
rect 30668 34202 30696 34410
rect 31220 34406 31248 35022
rect 31772 35018 31800 35566
rect 31864 35086 31892 36110
rect 32220 36032 32272 36038
rect 32220 35974 32272 35980
rect 32232 35630 32260 35974
rect 32220 35624 32272 35630
rect 32220 35566 32272 35572
rect 32036 35488 32088 35494
rect 32036 35430 32088 35436
rect 32048 35154 32076 35430
rect 32404 35284 32456 35290
rect 32404 35226 32456 35232
rect 32128 35216 32180 35222
rect 32128 35158 32180 35164
rect 32036 35148 32088 35154
rect 32036 35090 32088 35096
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 31760 35012 31812 35018
rect 31760 34954 31812 34960
rect 31668 34944 31720 34950
rect 31668 34886 31720 34892
rect 31680 34746 31708 34886
rect 31668 34740 31720 34746
rect 31668 34682 31720 34688
rect 31760 34672 31812 34678
rect 31760 34614 31812 34620
rect 31208 34400 31260 34406
rect 31208 34342 31260 34348
rect 30656 34196 30708 34202
rect 30656 34138 30708 34144
rect 31772 34066 31800 34614
rect 31760 34060 31812 34066
rect 31760 34002 31812 34008
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 29828 33924 29880 33930
rect 29828 33866 29880 33872
rect 29276 33652 29328 33658
rect 29276 33594 29328 33600
rect 28724 33516 28776 33522
rect 28724 33458 28776 33464
rect 29184 33516 29236 33522
rect 29184 33458 29236 33464
rect 28632 33108 28684 33114
rect 28632 33050 28684 33056
rect 28540 33040 28592 33046
rect 28540 32982 28592 32988
rect 28644 31822 28672 33050
rect 28736 32910 28764 33458
rect 29288 33454 29316 33594
rect 29736 33584 29788 33590
rect 29840 33572 29868 33866
rect 30380 33856 30432 33862
rect 30380 33798 30432 33804
rect 30656 33856 30708 33862
rect 30656 33798 30708 33804
rect 30392 33658 30420 33798
rect 30380 33652 30432 33658
rect 30380 33594 30432 33600
rect 29788 33544 29868 33572
rect 29736 33526 29788 33532
rect 29276 33448 29328 33454
rect 29276 33390 29328 33396
rect 29552 33380 29604 33386
rect 29552 33322 29604 33328
rect 29564 32910 29592 33322
rect 28724 32904 28776 32910
rect 28724 32846 28776 32852
rect 29552 32904 29604 32910
rect 29552 32846 29604 32852
rect 28736 32570 28764 32846
rect 28724 32564 28776 32570
rect 28724 32506 28776 32512
rect 29276 32496 29328 32502
rect 29276 32438 29328 32444
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28264 31476 28316 31482
rect 28264 31418 28316 31424
rect 28368 31470 28488 31498
rect 28368 31414 28396 31470
rect 27620 31408 27672 31414
rect 27620 31350 27672 31356
rect 28356 31408 28408 31414
rect 28356 31350 28408 31356
rect 27344 31340 27396 31346
rect 27344 31282 27396 31288
rect 28368 31278 28396 31350
rect 26792 31272 26844 31278
rect 26792 31214 26844 31220
rect 28356 31272 28408 31278
rect 28356 31214 28408 31220
rect 26424 29300 26476 29306
rect 26424 29242 26476 29248
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26332 29096 26384 29102
rect 26332 29038 26384 29044
rect 25780 29028 25832 29034
rect 25780 28970 25832 28976
rect 25792 28762 25820 28970
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 25780 28756 25832 28762
rect 25780 28698 25832 28704
rect 25596 28484 25648 28490
rect 25596 28426 25648 28432
rect 26252 28150 26280 28902
rect 26240 28144 26292 28150
rect 26240 28086 26292 28092
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25688 28076 25740 28082
rect 25688 28018 25740 28024
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 24780 27606 24808 27950
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24584 27532 24636 27538
rect 24584 27474 24636 27480
rect 24308 27396 24360 27402
rect 24308 27338 24360 27344
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 24032 26308 24084 26314
rect 24032 26250 24084 26256
rect 24044 26042 24072 26250
rect 24032 26036 24084 26042
rect 24032 25978 24084 25984
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23124 25498 23152 25842
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 24228 24818 24256 26930
rect 24320 26246 24348 27338
rect 24596 26926 24624 27474
rect 24780 27418 24808 27542
rect 25700 27538 25728 28018
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 26252 27606 26280 27950
rect 26344 27946 26372 29038
rect 26436 28558 26464 29242
rect 26528 28626 26556 29242
rect 26804 29170 26832 31214
rect 26976 31204 27028 31210
rect 26976 31146 27028 31152
rect 26988 30938 27016 31146
rect 26976 30932 27028 30938
rect 26976 30874 27028 30880
rect 29288 30326 29316 32438
rect 29276 30320 29328 30326
rect 29276 30262 29328 30268
rect 26976 30184 27028 30190
rect 26976 30126 27028 30132
rect 26988 29850 27016 30126
rect 27528 30048 27580 30054
rect 27528 29990 27580 29996
rect 26976 29844 27028 29850
rect 26976 29786 27028 29792
rect 27540 29714 27568 29990
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 28540 29776 28592 29782
rect 28540 29718 28592 29724
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 28552 29238 28580 29718
rect 28920 29714 28948 29786
rect 28908 29708 28960 29714
rect 28908 29650 28960 29656
rect 28540 29232 28592 29238
rect 28540 29174 28592 29180
rect 26792 29164 26844 29170
rect 26792 29106 26844 29112
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 26516 28620 26568 28626
rect 26516 28562 26568 28568
rect 26424 28552 26476 28558
rect 26424 28494 26476 28500
rect 27632 28422 27660 29038
rect 28920 28642 28948 29650
rect 29288 29238 29316 30262
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29276 29232 29328 29238
rect 29276 29174 29328 29180
rect 28920 28614 29224 28642
rect 28448 28552 28500 28558
rect 28448 28494 28500 28500
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 27632 28082 27660 28358
rect 28276 28150 28304 28358
rect 28460 28218 28488 28494
rect 28448 28212 28500 28218
rect 28448 28154 28500 28160
rect 28264 28144 28316 28150
rect 28264 28086 28316 28092
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 26976 28008 27028 28014
rect 26976 27950 27028 27956
rect 26332 27940 26384 27946
rect 26332 27882 26384 27888
rect 26240 27600 26292 27606
rect 26240 27542 26292 27548
rect 26988 27538 27016 27950
rect 27528 27872 27580 27878
rect 27528 27814 27580 27820
rect 27540 27674 27568 27814
rect 27528 27668 27580 27674
rect 27528 27610 27580 27616
rect 27632 27538 27660 28018
rect 27712 27668 27764 27674
rect 27712 27610 27764 27616
rect 28724 27668 28776 27674
rect 28920 27656 28948 28614
rect 29196 28558 29224 28614
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 29184 28552 29236 28558
rect 29184 28494 29236 28500
rect 28776 27628 28948 27656
rect 28724 27610 28776 27616
rect 25688 27532 25740 27538
rect 25688 27474 25740 27480
rect 26976 27532 27028 27538
rect 26976 27474 27028 27480
rect 27620 27532 27672 27538
rect 27620 27474 27672 27480
rect 25872 27464 25924 27470
rect 24780 27402 24900 27418
rect 25872 27406 25924 27412
rect 24780 27396 24912 27402
rect 24780 27390 24860 27396
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 24596 26518 24624 26862
rect 24584 26512 24636 26518
rect 24584 26454 24636 26460
rect 24780 26382 24808 27390
rect 24860 27338 24912 27344
rect 25884 27062 25912 27406
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 25872 27056 25924 27062
rect 25872 26998 25924 27004
rect 26436 26994 26464 27270
rect 26700 27056 26752 27062
rect 26700 26998 26752 27004
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24872 26382 24900 26726
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 25608 26314 25636 26930
rect 25596 26308 25648 26314
rect 25596 26250 25648 26256
rect 24308 26240 24360 26246
rect 24308 26182 24360 26188
rect 24320 25974 24348 26182
rect 24308 25968 24360 25974
rect 24308 25910 24360 25916
rect 25228 25900 25280 25906
rect 25228 25842 25280 25848
rect 24308 25696 24360 25702
rect 24308 25638 24360 25644
rect 24320 25294 24348 25638
rect 24308 25288 24360 25294
rect 24308 25230 24360 25236
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 24780 24886 24808 25094
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 22928 24744 22980 24750
rect 22928 24686 22980 24692
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22836 23792 22888 23798
rect 22836 23734 22888 23740
rect 22848 23186 22876 23734
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 22940 22574 22968 24686
rect 23308 24410 23336 24754
rect 25056 24410 25084 25094
rect 25240 24614 25268 25842
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 25240 24274 25268 24550
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 24768 24132 24820 24138
rect 24768 24074 24820 24080
rect 23204 23248 23256 23254
rect 23204 23190 23256 23196
rect 23216 22710 23244 23190
rect 23676 22710 23704 24074
rect 24780 23730 24808 24074
rect 25332 23730 25360 25094
rect 25504 24880 25556 24886
rect 25424 24840 25504 24868
rect 24768 23724 24820 23730
rect 24768 23666 24820 23672
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 24308 23588 24360 23594
rect 24308 23530 24360 23536
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23952 23118 23980 23462
rect 24320 23118 24348 23530
rect 24492 23520 24544 23526
rect 24492 23462 24544 23468
rect 24400 23180 24452 23186
rect 24400 23122 24452 23128
rect 23940 23112 23992 23118
rect 23940 23054 23992 23060
rect 24308 23112 24360 23118
rect 24308 23054 24360 23060
rect 23204 22704 23256 22710
rect 23204 22646 23256 22652
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 22928 22568 22980 22574
rect 22928 22510 22980 22516
rect 22652 22500 22704 22506
rect 22652 22442 22704 22448
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 22388 21554 22416 22374
rect 22940 22098 22968 22510
rect 23676 22438 23704 22646
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 22928 22092 22980 22098
rect 22928 22034 22980 22040
rect 24320 21962 24348 22374
rect 24308 21956 24360 21962
rect 24308 21898 24360 21904
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22572 21350 22600 21422
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22282 20496 22338 20505
rect 22282 20431 22338 20440
rect 22284 20392 22336 20398
rect 22204 20352 22284 20380
rect 22204 19786 22232 20352
rect 22284 20334 22336 20340
rect 22388 20262 22416 21082
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 21836 19502 22048 19530
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21456 18692 21508 18698
rect 21456 18634 21508 18640
rect 21744 18630 21772 18702
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19536 16658 19564 16934
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19628 16046 19656 17614
rect 21284 17610 21312 18158
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21560 17338 21588 17546
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19904 16250 19932 17138
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19996 16522 20024 17002
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19996 16425 20024 16458
rect 19982 16416 20038 16425
rect 19982 16351 20038 16360
rect 20180 16250 20208 17070
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20272 16658 20300 16934
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20272 16114 20300 16594
rect 21100 16454 21128 17070
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21100 16182 21128 16390
rect 21192 16250 21220 16390
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19168 14498 19196 14962
rect 19260 14890 19288 15370
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15026 19472 15302
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19260 14793 19288 14826
rect 19246 14784 19302 14793
rect 19246 14719 19302 14728
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19168 14470 19288 14498
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18156 13138 18184 13194
rect 18708 13190 18736 13874
rect 18064 13110 18184 13138
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18064 12918 18092 13110
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17788 12406 17908 12434
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17420 11354 17448 11630
rect 17696 11354 17724 11834
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17052 11082 17080 11290
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 17604 10674 17632 11154
rect 17788 11150 17816 12406
rect 18708 12306 18736 13126
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11898 18460 12038
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 18432 11014 18460 11834
rect 18616 11694 18644 12106
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 17144 9586 17172 10134
rect 17236 10130 17264 10610
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17328 9722 17356 9862
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17328 9586 17356 9658
rect 17604 9586 17632 10610
rect 17788 10130 17816 10950
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17880 10062 17908 10406
rect 17972 10266 18000 10950
rect 18328 10736 18380 10742
rect 18248 10696 18328 10724
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18156 10266 18184 10542
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 17972 10062 18000 10202
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 18248 9722 18276 10696
rect 18328 10678 18380 10684
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 10062 18552 10406
rect 18708 10130 18736 12242
rect 19076 12170 19104 14350
rect 19168 12986 19196 14350
rect 19260 13852 19288 14470
rect 19352 14006 19380 14554
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19444 13852 19472 13942
rect 19536 13870 19564 15098
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19720 14074 19748 14962
rect 19996 14890 20024 14962
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19996 13938 20024 14554
rect 20180 14074 20208 15982
rect 20272 15162 20300 16050
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20548 15366 20576 15982
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15570 20760 15846
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20364 14618 20392 14962
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19260 13824 19472 13852
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19168 12238 19196 12922
rect 19444 12850 19472 13466
rect 19536 13326 19564 13806
rect 19628 13734 19656 13806
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19628 13326 19656 13670
rect 20180 13530 20208 14010
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20180 13326 20208 13466
rect 20272 13394 20300 13942
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19904 12850 19932 13126
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 20272 12714 20300 13330
rect 20456 12782 20484 13874
rect 20548 13734 20576 14758
rect 20732 13802 20760 15030
rect 20824 14958 20852 16050
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15094 21312 15846
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 21100 13530 21128 14282
rect 21560 14074 21588 14282
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 19352 11694 19380 12582
rect 19628 12306 19656 12650
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11762 20392 12038
rect 20456 11898 20484 12718
rect 20732 12238 20760 13466
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12850 21128 13126
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 12442 20852 12650
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 18786 11520 18842 11529
rect 18786 11455 18842 11464
rect 18800 11150 18828 11455
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 20996 11076 21048 11082
rect 21192 11064 21220 13194
rect 21560 12986 21588 13262
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21652 12986 21680 13194
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21048 11036 21220 11064
rect 20996 11018 21048 11024
rect 21008 10742 21036 11018
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16960 9178 16988 9454
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17328 8634 17356 9522
rect 17604 9382 17632 9522
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17972 9178 18000 9454
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17236 7954 17264 8230
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 7342 16712 7822
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 7478 16988 7686
rect 17788 7546 17816 8366
rect 18248 7818 18276 9658
rect 18340 8974 18368 9930
rect 18708 9042 18736 10066
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19260 9450 19288 9930
rect 19720 9518 19748 10542
rect 20732 10266 20760 10542
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 21008 9654 21036 10678
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18328 8968 18380 8974
rect 18708 8922 18736 8978
rect 18328 8910 18380 8916
rect 18616 8894 18736 8922
rect 18616 8430 18644 8894
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8634 18736 8774
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18708 8090 18736 8570
rect 21008 8566 21036 9590
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 18248 7478 18276 7754
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16684 6322 16712 7278
rect 19628 6730 19656 8366
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 18524 6322 18552 6666
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 16684 5710 16712 6258
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 15856 4690 15884 5646
rect 18524 5234 18552 6258
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18524 4690 18552 5170
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 19996 4554 20024 7414
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20732 7002 20760 7142
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 21008 6866 21036 8502
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21192 7410 21220 7958
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21192 5166 21220 5510
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 21284 2774 21312 11494
rect 21468 11150 21496 11562
rect 21836 11354 21864 19502
rect 22480 18834 22508 20878
rect 22572 20262 22600 21286
rect 22652 21072 22704 21078
rect 22652 21014 22704 21020
rect 22664 20466 22692 21014
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 23032 20398 23060 20878
rect 23308 20505 23336 20878
rect 23480 20868 23532 20874
rect 23480 20810 23532 20816
rect 23294 20496 23350 20505
rect 23492 20466 23520 20810
rect 23860 20534 23888 21286
rect 24320 20534 24348 21898
rect 24412 21010 24440 23122
rect 24504 22982 24532 23462
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24780 22710 24808 23666
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24964 23050 24992 23462
rect 25424 23050 25452 24840
rect 25608 24868 25636 26250
rect 26068 26042 26096 26930
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26528 26586 26556 26862
rect 26712 26858 26740 26998
rect 26700 26852 26752 26858
rect 26700 26794 26752 26800
rect 26516 26580 26568 26586
rect 26516 26522 26568 26528
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 25872 25832 25924 25838
rect 25872 25774 25924 25780
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25556 24840 25636 24868
rect 25504 24822 25556 24828
rect 25700 24410 25728 25434
rect 25884 25158 25912 25774
rect 26344 25226 26372 25842
rect 26896 25770 26924 27338
rect 27632 26450 27660 27474
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 27724 25838 27752 27610
rect 29012 27606 29040 28494
rect 29288 28150 29316 29174
rect 29276 28144 29328 28150
rect 29276 28086 29328 28092
rect 29000 27600 29052 27606
rect 29000 27542 29052 27548
rect 28264 27396 28316 27402
rect 28264 27338 28316 27344
rect 27988 27328 28040 27334
rect 27988 27270 28040 27276
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28000 27062 28028 27270
rect 27988 27056 28040 27062
rect 27988 26998 28040 27004
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 27896 26852 27948 26858
rect 27896 26794 27948 26800
rect 27804 26512 27856 26518
rect 27804 26454 27856 26460
rect 27816 25906 27844 26454
rect 27908 26450 27936 26794
rect 27896 26444 27948 26450
rect 27896 26386 27948 26392
rect 27804 25900 27856 25906
rect 27804 25842 27856 25848
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 26884 25764 26936 25770
rect 26884 25706 26936 25712
rect 27528 25764 27580 25770
rect 27528 25706 27580 25712
rect 26896 25226 26924 25706
rect 26976 25492 27028 25498
rect 26976 25434 27028 25440
rect 26332 25220 26384 25226
rect 26332 25162 26384 25168
rect 26884 25220 26936 25226
rect 26884 25162 26936 25168
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 26252 24342 26280 24550
rect 26344 24410 26372 25162
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 26332 24404 26384 24410
rect 26332 24346 26384 24352
rect 26240 24336 26292 24342
rect 26240 24278 26292 24284
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25608 24070 25636 24142
rect 26436 24070 26464 24754
rect 26988 24750 27016 25434
rect 27540 25430 27568 25706
rect 27528 25424 27580 25430
rect 27528 25366 27580 25372
rect 27436 25152 27488 25158
rect 27436 25094 27488 25100
rect 27448 24818 27476 25094
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 26976 24744 27028 24750
rect 26976 24686 27028 24692
rect 26700 24676 26752 24682
rect 26700 24618 26752 24624
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 26712 24206 26740 24618
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26712 24070 26740 24142
rect 27172 24138 27200 24618
rect 27252 24268 27304 24274
rect 27252 24210 27304 24216
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 26424 24064 26476 24070
rect 26424 24006 26476 24012
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 25424 22094 25452 22986
rect 25516 22778 25544 23666
rect 25608 23594 25636 24006
rect 26240 23656 26292 23662
rect 26240 23598 26292 23604
rect 25596 23588 25648 23594
rect 25596 23530 25648 23536
rect 26252 23186 26280 23598
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26436 23118 26464 24006
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26620 23118 26648 23462
rect 26424 23112 26476 23118
rect 26422 23080 26424 23089
rect 26608 23112 26660 23118
rect 26476 23080 26478 23089
rect 26608 23054 26660 23060
rect 26422 23015 26478 23024
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 26436 22574 26464 23015
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26424 22568 26476 22574
rect 26424 22510 26476 22516
rect 25424 22066 25544 22094
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 21146 25176 21422
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 24400 21004 24452 21010
rect 24400 20946 24452 20952
rect 25516 20874 25544 22066
rect 26620 22030 26648 22578
rect 26712 22574 26740 24006
rect 27172 23730 27200 24074
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 26884 23588 26936 23594
rect 26884 23530 26936 23536
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26804 22778 26832 23054
rect 26792 22772 26844 22778
rect 26792 22714 26844 22720
rect 26700 22568 26752 22574
rect 26700 22510 26752 22516
rect 26896 22506 26924 23530
rect 27172 22642 27200 23666
rect 27264 23118 27292 24210
rect 27448 24206 27476 24754
rect 27436 24200 27488 24206
rect 27356 24160 27436 24188
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 26884 22500 26936 22506
rect 26884 22442 26936 22448
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 25872 21956 25924 21962
rect 25872 21898 25924 21904
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25792 21554 25820 21830
rect 25884 21554 25912 21898
rect 25964 21616 26016 21622
rect 25964 21558 26016 21564
rect 25780 21548 25832 21554
rect 25780 21490 25832 21496
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25504 20868 25556 20874
rect 25504 20810 25556 20816
rect 25516 20534 25544 20810
rect 23848 20528 23900 20534
rect 23848 20470 23900 20476
rect 24308 20528 24360 20534
rect 24308 20470 24360 20476
rect 25504 20528 25556 20534
rect 25504 20470 25556 20476
rect 23294 20431 23296 20440
rect 23348 20431 23350 20440
rect 23480 20460 23532 20466
rect 23296 20402 23348 20408
rect 23480 20402 23532 20408
rect 23020 20392 23072 20398
rect 23388 20392 23440 20398
rect 23072 20352 23244 20380
rect 23020 20334 23072 20340
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22756 19854 22784 20198
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 21928 18086 21956 18702
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 22020 17592 22048 18770
rect 22480 18290 22508 18770
rect 22756 18766 22784 19790
rect 22940 19446 22968 19790
rect 22928 19440 22980 19446
rect 22928 19382 22980 19388
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22940 18426 22968 19382
rect 23032 19378 23060 20198
rect 23216 19854 23244 20352
rect 23388 20334 23440 20340
rect 23400 20058 23428 20334
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23664 19984 23716 19990
rect 23664 19926 23716 19932
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23204 19848 23256 19854
rect 23204 19790 23256 19796
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23020 19372 23072 19378
rect 23020 19314 23072 19320
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22100 17604 22152 17610
rect 22020 17564 22100 17592
rect 22020 16590 22048 17564
rect 22100 17546 22152 17552
rect 22836 17604 22888 17610
rect 22836 17546 22888 17552
rect 22848 17338 22876 17546
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22020 15434 22048 16526
rect 22112 15434 22140 16526
rect 23032 16522 23060 16594
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 23020 16516 23072 16522
rect 23020 16458 23072 16464
rect 22572 16250 22600 16458
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 23124 15706 23152 19110
rect 23216 18766 23244 19654
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23216 15978 23244 17070
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22020 15162 22048 15370
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22020 14278 22048 15098
rect 22112 14958 22140 15370
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22112 14414 22140 14894
rect 22480 14618 22508 14894
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22100 14408 22152 14414
rect 23124 14385 23152 15642
rect 23216 14822 23244 15914
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23400 14498 23428 18770
rect 23492 18358 23520 19858
rect 23676 19718 23704 19926
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23676 19174 23704 19654
rect 23952 19378 23980 19722
rect 24044 19378 24072 19790
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23952 18970 23980 19314
rect 23940 18964 23992 18970
rect 23940 18906 23992 18912
rect 23952 18766 23980 18906
rect 23940 18760 23992 18766
rect 24044 18748 24072 19314
rect 24124 18760 24176 18766
rect 24044 18720 24124 18748
rect 23940 18702 23992 18708
rect 24124 18702 24176 18708
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23492 17202 23520 18294
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23584 17746 23612 18226
rect 23768 18154 23796 18566
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23584 17134 23612 17682
rect 23768 17542 23796 18090
rect 23952 17678 23980 18158
rect 24136 17678 24164 18566
rect 23940 17672 23992 17678
rect 24124 17672 24176 17678
rect 23992 17632 24072 17660
rect 23940 17614 23992 17620
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23860 17184 23888 17546
rect 23940 17196 23992 17202
rect 23860 17156 23940 17184
rect 23940 17138 23992 17144
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 24044 16658 24072 17632
rect 24124 17614 24176 17620
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24136 17202 24164 17478
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23952 15366 23980 16458
rect 24044 16454 24072 16594
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24044 16250 24072 16390
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24136 16182 24164 17138
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24136 15366 24164 15506
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 23676 14906 23704 15302
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23584 14878 23704 14906
rect 23400 14482 23520 14498
rect 23400 14476 23532 14482
rect 23400 14470 23480 14476
rect 22100 14350 22152 14356
rect 23110 14376 23166 14385
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22112 14006 22140 14350
rect 23110 14311 23166 14320
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 23400 13954 23428 14470
rect 23480 14418 23532 14424
rect 23584 14346 23612 14878
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 23400 13938 23520 13954
rect 23400 13932 23532 13938
rect 23400 13926 23480 13932
rect 22100 13864 22152 13870
rect 21914 13832 21970 13841
rect 22100 13806 22152 13812
rect 21914 13767 21970 13776
rect 21928 13530 21956 13767
rect 22112 13530 22140 13806
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 23400 13326 23428 13926
rect 23480 13874 23532 13880
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23124 12306 23152 13126
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23492 12306 23520 12582
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 22020 11762 22048 12038
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 23124 11626 23152 12242
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 22296 10810 22324 11494
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21376 8022 21404 10066
rect 21468 10062 21496 10406
rect 21836 10198 21864 10406
rect 21824 10192 21876 10198
rect 21824 10134 21876 10140
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21928 9926 21956 10134
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 21560 9518 21588 9862
rect 21928 9654 21956 9862
rect 22204 9654 22232 9862
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 22388 9586 22416 10406
rect 22480 10305 22508 10542
rect 22756 10538 22784 10950
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 22940 10674 22968 10746
rect 23216 10674 23244 12038
rect 23400 11830 23428 12174
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23492 11762 23520 12242
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 22744 10532 22796 10538
rect 22744 10474 22796 10480
rect 22466 10296 22522 10305
rect 22466 10231 22522 10240
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23124 10033 23152 10066
rect 23216 10062 23244 10610
rect 23308 10062 23336 10746
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23400 10169 23428 10202
rect 23386 10160 23442 10169
rect 23386 10095 23442 10104
rect 23204 10056 23256 10062
rect 23110 10024 23166 10033
rect 23204 9998 23256 10004
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23110 9959 23166 9968
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9586 22968 9862
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 23032 9518 23060 9658
rect 23124 9568 23152 9959
rect 23492 9722 23520 10610
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 23204 9580 23256 9586
rect 23124 9540 23204 9568
rect 23204 9522 23256 9528
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21640 8900 21692 8906
rect 21640 8842 21692 8848
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21468 7886 21496 8366
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21376 7546 21404 7822
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21652 7342 21680 8842
rect 21744 7886 21772 9046
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21836 8566 21864 8774
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 21824 8560 21876 8566
rect 21824 8502 21876 8508
rect 21732 7880 21784 7886
rect 22296 7834 22324 8570
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 21732 7822 21784 7828
rect 22020 7818 22324 7834
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 22008 7812 22324 7818
rect 22060 7806 22324 7812
rect 22008 7754 22060 7760
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21468 7002 21496 7278
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21376 5302 21404 6666
rect 21744 5778 21772 7210
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 21744 5098 21772 5714
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21744 4690 21772 5034
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21744 4146 21772 4626
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 21836 4078 21864 7754
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22112 7410 22140 7686
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22020 5642 22048 6258
rect 22296 6254 22324 7806
rect 22388 7750 22416 8298
rect 22480 7886 22508 8434
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22008 5636 22060 5642
rect 22008 5578 22060 5584
rect 22020 5370 22048 5578
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 22020 4554 22048 5306
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22008 4548 22060 4554
rect 22008 4490 22060 4496
rect 22020 4214 22048 4490
rect 22008 4208 22060 4214
rect 22008 4150 22060 4156
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 22204 3398 22232 4966
rect 22296 4622 22324 6190
rect 22376 5840 22428 5846
rect 22376 5782 22428 5788
rect 22388 5234 22416 5782
rect 22572 5778 22600 6598
rect 22652 6180 22704 6186
rect 22652 6122 22704 6128
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22664 5710 22692 6122
rect 22756 6118 22784 7482
rect 22940 7410 22968 9318
rect 23032 8090 23060 9454
rect 23216 8974 23244 9522
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23216 8498 23244 8910
rect 23478 8528 23534 8537
rect 23204 8492 23256 8498
rect 23478 8463 23480 8472
rect 23204 8434 23256 8440
rect 23532 8463 23534 8472
rect 23480 8434 23532 8440
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23308 7886 23336 8026
rect 23020 7880 23072 7886
rect 23296 7880 23348 7886
rect 23020 7822 23072 7828
rect 23216 7840 23296 7868
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22756 5794 22784 6054
rect 22940 5930 22968 7346
rect 23032 6458 23060 7822
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 22848 5914 22968 5930
rect 22836 5908 22968 5914
rect 22888 5902 22968 5908
rect 22836 5850 22888 5856
rect 22756 5778 22876 5794
rect 22756 5772 22888 5778
rect 22756 5766 22836 5772
rect 22836 5714 22888 5720
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22296 4282 22324 4558
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22388 3942 22416 4490
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22664 3466 22692 5306
rect 22848 5234 22876 5714
rect 22940 5370 22968 5902
rect 23032 5710 23060 6394
rect 23216 6254 23244 7840
rect 23296 7822 23348 7828
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23308 7478 23336 7686
rect 23296 7472 23348 7478
rect 23296 7414 23348 7420
rect 23296 7268 23348 7274
rect 23296 7210 23348 7216
rect 23204 6248 23256 6254
rect 23204 6190 23256 6196
rect 23216 5710 23244 6190
rect 23308 5778 23336 7210
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23492 6458 23520 6734
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 23308 5302 23336 5510
rect 23296 5296 23348 5302
rect 23296 5238 23348 5244
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22756 4554 22784 5170
rect 23492 4826 23520 5646
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 23112 4548 23164 4554
rect 23112 4490 23164 4496
rect 23124 4282 23152 4490
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22652 3460 22704 3466
rect 22652 3402 22704 3408
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22756 3126 22784 3878
rect 23400 3738 23428 4558
rect 23584 3738 23612 14282
rect 23860 14006 23888 15030
rect 24136 14958 24164 15302
rect 24228 15026 24256 19382
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24872 18766 24900 19246
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24872 18426 24900 18702
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24872 17882 24900 18226
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 24504 17202 24532 17546
rect 24780 17202 24808 17614
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24872 17338 24900 17478
rect 24964 17338 24992 20198
rect 25792 19496 25820 21490
rect 25884 20602 25912 21490
rect 25976 20602 26004 21558
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25964 20596 26016 20602
rect 25964 20538 26016 20544
rect 26252 20466 26280 21354
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26344 20466 26372 20742
rect 26620 20602 26648 21966
rect 26792 21684 26844 21690
rect 26792 21626 26844 21632
rect 26700 21344 26752 21350
rect 26700 21286 26752 21292
rect 26608 20596 26660 20602
rect 26608 20538 26660 20544
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 26068 19854 26096 20334
rect 26252 19854 26280 20402
rect 26344 19854 26372 20402
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26068 19514 26096 19790
rect 26056 19508 26108 19514
rect 25792 19468 25912 19496
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25332 18766 25360 19314
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25424 18766 25452 19246
rect 25792 18970 25820 19314
rect 25780 18964 25832 18970
rect 25780 18906 25832 18912
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25332 18426 25360 18702
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25424 18086 25452 18702
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25516 17678 25544 18158
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24872 16726 24900 16934
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24964 16114 24992 17274
rect 25240 17202 25268 17614
rect 25608 17202 25636 17682
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25240 16794 25268 17138
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 25424 16658 25452 17138
rect 25884 16998 25912 19468
rect 26056 19450 26108 19456
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 25976 18834 26004 19314
rect 26344 19242 26372 19790
rect 26712 19378 26740 21286
rect 26804 20942 26832 21626
rect 26896 21146 26924 22442
rect 26976 22432 27028 22438
rect 27264 22420 27292 23054
rect 27356 22574 27384 24160
rect 27436 24142 27488 24148
rect 27540 23662 27568 25366
rect 27908 25362 27936 25842
rect 28092 25838 28120 26930
rect 28184 26586 28212 27270
rect 28276 26790 28304 27338
rect 29656 27334 29684 30194
rect 29840 30138 29868 33544
rect 30668 33114 30696 33798
rect 31024 33448 31076 33454
rect 31024 33390 31076 33396
rect 30748 33312 30800 33318
rect 30748 33254 30800 33260
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30760 32910 30788 33254
rect 31036 32978 31064 33390
rect 31668 33108 31720 33114
rect 31668 33050 31720 33056
rect 31024 32972 31076 32978
rect 31024 32914 31076 32920
rect 30748 32904 30800 32910
rect 30748 32846 30800 32852
rect 31036 32842 31064 32914
rect 31680 32910 31708 33050
rect 31668 32904 31720 32910
rect 31668 32846 31720 32852
rect 30012 32836 30064 32842
rect 30012 32778 30064 32784
rect 31024 32836 31076 32842
rect 31024 32778 31076 32784
rect 30024 32434 30052 32778
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 30288 32428 30340 32434
rect 30288 32370 30340 32376
rect 31392 32428 31444 32434
rect 31392 32370 31444 32376
rect 30300 31890 30328 32370
rect 30564 32360 30616 32366
rect 30564 32302 30616 32308
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 29920 31136 29972 31142
rect 29920 31078 29972 31084
rect 29932 30666 29960 31078
rect 30300 30802 30328 31826
rect 30472 31136 30524 31142
rect 30472 31078 30524 31084
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 29920 30660 29972 30666
rect 29920 30602 29972 30608
rect 30300 30326 30328 30738
rect 30484 30326 30512 31078
rect 30288 30320 30340 30326
rect 30288 30262 30340 30268
rect 30472 30320 30524 30326
rect 30472 30262 30524 30268
rect 29840 30110 29960 30138
rect 29932 30054 29960 30110
rect 29920 30048 29972 30054
rect 29920 29990 29972 29996
rect 29736 29708 29788 29714
rect 29736 29650 29788 29656
rect 29748 28558 29776 29650
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29840 29306 29868 29582
rect 29828 29300 29880 29306
rect 29828 29242 29880 29248
rect 29736 28552 29788 28558
rect 29788 28500 29868 28506
rect 29736 28494 29868 28500
rect 29748 28478 29868 28494
rect 29840 28422 29868 28478
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 29828 28416 29880 28422
rect 29828 28358 29880 28364
rect 29748 28218 29776 28358
rect 29736 28212 29788 28218
rect 29736 28154 29788 28160
rect 29932 28150 29960 29990
rect 30300 29782 30328 30262
rect 30576 29850 30604 32302
rect 30656 32224 30708 32230
rect 30656 32166 30708 32172
rect 30668 31890 30696 32166
rect 31404 32026 31432 32370
rect 31392 32020 31444 32026
rect 31392 31962 31444 31968
rect 30656 31884 30708 31890
rect 30656 31826 30708 31832
rect 30840 30320 30892 30326
rect 30840 30262 30892 30268
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 30288 29776 30340 29782
rect 30288 29718 30340 29724
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 30024 28762 30052 29242
rect 30196 29164 30248 29170
rect 30300 29152 30328 29718
rect 30380 29504 30432 29510
rect 30380 29446 30432 29452
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30392 29238 30420 29446
rect 30380 29232 30432 29238
rect 30380 29174 30432 29180
rect 30248 29124 30328 29152
rect 30196 29106 30248 29112
rect 30484 28762 30512 29446
rect 30852 29306 30880 30262
rect 31116 29504 31168 29510
rect 31116 29446 31168 29452
rect 30840 29300 30892 29306
rect 30840 29242 30892 29248
rect 30012 28756 30064 28762
rect 30012 28698 30064 28704
rect 30472 28756 30524 28762
rect 30472 28698 30524 28704
rect 30024 28558 30052 28698
rect 30196 28688 30248 28694
rect 30196 28630 30248 28636
rect 30208 28558 30236 28630
rect 31128 28626 31156 29446
rect 31484 29096 31536 29102
rect 31484 29038 31536 29044
rect 31496 28762 31524 29038
rect 31680 28762 31708 32846
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 31772 31278 31800 32370
rect 31864 31890 31892 35022
rect 31944 34944 31996 34950
rect 31944 34886 31996 34892
rect 31956 34542 31984 34886
rect 32048 34610 32076 35090
rect 32036 34604 32088 34610
rect 32036 34546 32088 34552
rect 32140 34542 32168 35158
rect 32416 34610 32444 35226
rect 33152 35170 33180 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 38474 36136 38530 36145
rect 38474 36071 38476 36080
rect 38528 36071 38530 36080
rect 38476 36042 38528 36048
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 38476 35488 38528 35494
rect 38474 35456 38476 35465
rect 38528 35456 38530 35465
rect 34934 35388 35242 35397
rect 38474 35391 38530 35400
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 33152 35154 33364 35170
rect 33152 35148 33376 35154
rect 33152 35142 33324 35148
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 33152 34542 33180 35142
rect 33324 35090 33376 35096
rect 38476 34944 38528 34950
rect 38476 34886 38528 34892
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 38488 34785 38516 34886
rect 38474 34776 38530 34785
rect 38474 34711 38530 34720
rect 31944 34536 31996 34542
rect 31944 34478 31996 34484
rect 32128 34536 32180 34542
rect 32128 34478 32180 34484
rect 32772 34536 32824 34542
rect 32772 34478 32824 34484
rect 33140 34536 33192 34542
rect 33140 34478 33192 34484
rect 32784 33114 32812 34478
rect 33152 34066 33180 34478
rect 38476 34400 38528 34406
rect 38476 34342 38528 34348
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 38488 34105 38516 34342
rect 38474 34096 38530 34105
rect 33140 34060 33192 34066
rect 38474 34031 38530 34040
rect 33140 34002 33192 34008
rect 33152 33522 33180 34002
rect 34796 33856 34848 33862
rect 34796 33798 34848 33804
rect 34808 33590 34836 33798
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 34796 33584 34848 33590
rect 34796 33526 34848 33532
rect 35532 33584 35584 33590
rect 35532 33526 35584 33532
rect 33140 33516 33192 33522
rect 33140 33458 33192 33464
rect 33508 33448 33560 33454
rect 33508 33390 33560 33396
rect 33600 33448 33652 33454
rect 33600 33390 33652 33396
rect 34244 33448 34296 33454
rect 34244 33390 34296 33396
rect 33520 33114 33548 33390
rect 32772 33108 32824 33114
rect 32772 33050 32824 33056
rect 33508 33108 33560 33114
rect 33508 33050 33560 33056
rect 33324 32972 33376 32978
rect 33324 32914 33376 32920
rect 32128 32836 32180 32842
rect 32128 32778 32180 32784
rect 32140 32570 32168 32778
rect 32128 32564 32180 32570
rect 32128 32506 32180 32512
rect 33140 32360 33192 32366
rect 33140 32302 33192 32308
rect 33152 32008 33180 32302
rect 33336 32298 33364 32914
rect 33508 32768 33560 32774
rect 33508 32710 33560 32716
rect 33520 32434 33548 32710
rect 33612 32434 33640 33390
rect 34256 32910 34284 33390
rect 34520 33380 34572 33386
rect 34520 33322 34572 33328
rect 34336 33040 34388 33046
rect 34336 32982 34388 32988
rect 33876 32904 33928 32910
rect 33876 32846 33928 32852
rect 34244 32904 34296 32910
rect 34244 32846 34296 32852
rect 33888 32570 33916 32846
rect 33876 32564 33928 32570
rect 33876 32506 33928 32512
rect 33508 32428 33560 32434
rect 33508 32370 33560 32376
rect 33600 32428 33652 32434
rect 33600 32370 33652 32376
rect 33876 32428 33928 32434
rect 33876 32370 33928 32376
rect 33324 32292 33376 32298
rect 33324 32234 33376 32240
rect 33416 32224 33468 32230
rect 33416 32166 33468 32172
rect 33232 32020 33284 32026
rect 33152 31980 33232 32008
rect 31852 31884 31904 31890
rect 31852 31826 31904 31832
rect 31760 31272 31812 31278
rect 31760 31214 31812 31220
rect 31772 30938 31800 31214
rect 31760 30932 31812 30938
rect 31760 30874 31812 30880
rect 31864 30666 31892 31826
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 32784 31346 32812 31758
rect 33152 31346 33180 31980
rect 33232 31962 33284 31968
rect 33428 31754 33456 32166
rect 33336 31726 33456 31754
rect 32772 31340 32824 31346
rect 32772 31282 32824 31288
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 32588 31136 32640 31142
rect 32588 31078 32640 31084
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 31852 30660 31904 30666
rect 31852 30602 31904 30608
rect 32128 30660 32180 30666
rect 32128 30602 32180 30608
rect 31864 30394 31892 30602
rect 31852 30388 31904 30394
rect 31852 30330 31904 30336
rect 32140 30258 32168 30602
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 32324 30122 32352 30670
rect 32600 30258 32628 31078
rect 32784 30870 32812 31282
rect 33140 31136 33192 31142
rect 33140 31078 33192 31084
rect 32772 30864 32824 30870
rect 32772 30806 32824 30812
rect 33152 30734 33180 31078
rect 33336 30938 33364 31726
rect 33520 31498 33548 32370
rect 33612 32026 33640 32370
rect 33600 32020 33652 32026
rect 33600 31962 33652 31968
rect 33428 31470 33548 31498
rect 33428 31142 33456 31470
rect 33508 31340 33560 31346
rect 33508 31282 33560 31288
rect 33416 31136 33468 31142
rect 33416 31078 33468 31084
rect 33324 30932 33376 30938
rect 33324 30874 33376 30880
rect 32864 30728 32916 30734
rect 32864 30670 32916 30676
rect 33140 30728 33192 30734
rect 33140 30670 33192 30676
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 32588 30252 32640 30258
rect 32588 30194 32640 30200
rect 32312 30116 32364 30122
rect 32312 30058 32364 30064
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 31852 29572 31904 29578
rect 31852 29514 31904 29520
rect 31864 28966 31892 29514
rect 31852 28960 31904 28966
rect 31852 28902 31904 28908
rect 31484 28756 31536 28762
rect 31484 28698 31536 28704
rect 31668 28756 31720 28762
rect 31668 28698 31720 28704
rect 31116 28620 31168 28626
rect 31116 28562 31168 28568
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 30748 28484 30800 28490
rect 30748 28426 30800 28432
rect 31116 28484 31168 28490
rect 31116 28426 31168 28432
rect 30760 28218 30788 28426
rect 30748 28212 30800 28218
rect 30748 28154 30800 28160
rect 29920 28144 29972 28150
rect 29920 28086 29972 28092
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 29828 27668 29880 27674
rect 29828 27610 29880 27616
rect 28816 27328 28868 27334
rect 28816 27270 28868 27276
rect 29644 27328 29696 27334
rect 29644 27270 29696 27276
rect 28264 26784 28316 26790
rect 28264 26726 28316 26732
rect 28172 26580 28224 26586
rect 28172 26522 28224 26528
rect 28276 26382 28304 26726
rect 28828 26518 28856 27270
rect 29656 27062 29684 27270
rect 29644 27056 29696 27062
rect 29644 26998 29696 27004
rect 29656 26586 29684 26998
rect 29644 26580 29696 26586
rect 29644 26522 29696 26528
rect 28816 26512 28868 26518
rect 28816 26454 28868 26460
rect 28264 26376 28316 26382
rect 28264 26318 28316 26324
rect 29092 26376 29144 26382
rect 29092 26318 29144 26324
rect 28540 26308 28592 26314
rect 28540 26250 28592 26256
rect 28080 25832 28132 25838
rect 28080 25774 28132 25780
rect 27896 25356 27948 25362
rect 27896 25298 27948 25304
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28000 24410 28028 25230
rect 27988 24404 28040 24410
rect 27988 24346 28040 24352
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27528 23656 27580 23662
rect 27528 23598 27580 23604
rect 27540 23497 27568 23598
rect 27526 23488 27582 23497
rect 27526 23423 27582 23432
rect 27724 22778 27752 24006
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27816 23118 27844 23462
rect 28184 23322 28212 25230
rect 28264 24336 28316 24342
rect 28264 24278 28316 24284
rect 28276 23322 28304 24278
rect 28552 23798 28580 26250
rect 29104 25702 29132 26318
rect 29184 26240 29236 26246
rect 29184 26182 29236 26188
rect 29196 26042 29224 26182
rect 29184 26036 29236 26042
rect 29184 25978 29236 25984
rect 29656 25974 29684 26522
rect 29840 26450 29868 27610
rect 30760 27470 30788 28018
rect 31128 28014 31156 28426
rect 31496 28150 31524 28698
rect 31484 28144 31536 28150
rect 31404 28104 31484 28132
rect 30840 28008 30892 28014
rect 30840 27950 30892 27956
rect 31116 28008 31168 28014
rect 31116 27950 31168 27956
rect 30852 27538 30880 27950
rect 31404 27674 31432 28104
rect 31484 28086 31536 28092
rect 31484 27872 31536 27878
rect 31484 27814 31536 27820
rect 31392 27668 31444 27674
rect 31392 27610 31444 27616
rect 30840 27532 30892 27538
rect 30840 27474 30892 27480
rect 31116 27532 31168 27538
rect 31116 27474 31168 27480
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30852 26874 30880 27474
rect 31024 26988 31076 26994
rect 31024 26930 31076 26936
rect 30760 26846 30880 26874
rect 30760 26790 30788 26846
rect 30748 26784 30800 26790
rect 30748 26726 30800 26732
rect 29828 26444 29880 26450
rect 29828 26386 29880 26392
rect 30104 26444 30156 26450
rect 30104 26386 30156 26392
rect 29840 26042 29868 26386
rect 30116 26314 30144 26386
rect 30104 26308 30156 26314
rect 30104 26250 30156 26256
rect 29828 26036 29880 26042
rect 29828 25978 29880 25984
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29828 25900 29880 25906
rect 29828 25842 29880 25848
rect 29092 25696 29144 25702
rect 29092 25638 29144 25644
rect 29092 25220 29144 25226
rect 29092 25162 29144 25168
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28644 24410 28672 24754
rect 29104 24750 29132 25162
rect 29840 25158 29868 25842
rect 30116 25480 30144 26250
rect 30288 26036 30340 26042
rect 30288 25978 30340 25984
rect 29932 25452 30144 25480
rect 29828 25152 29880 25158
rect 29828 25094 29880 25100
rect 29092 24744 29144 24750
rect 29092 24686 29144 24692
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29000 24676 29052 24682
rect 29000 24618 29052 24624
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28816 24268 28868 24274
rect 28816 24210 28868 24216
rect 28828 24070 28856 24210
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 28908 24064 28960 24070
rect 28908 24006 28960 24012
rect 28540 23792 28592 23798
rect 28540 23734 28592 23740
rect 28172 23316 28224 23322
rect 28172 23258 28224 23264
rect 28264 23316 28316 23322
rect 28264 23258 28316 23264
rect 27896 23248 27948 23254
rect 27896 23190 27948 23196
rect 27908 23118 27936 23190
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 28356 23112 28408 23118
rect 28448 23112 28500 23118
rect 28356 23054 28408 23060
rect 28446 23080 28448 23089
rect 28540 23112 28592 23118
rect 28500 23080 28502 23089
rect 27712 22772 27764 22778
rect 27712 22714 27764 22720
rect 27724 22574 27752 22714
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27436 22500 27488 22506
rect 27436 22442 27488 22448
rect 27344 22432 27396 22438
rect 27264 22392 27344 22420
rect 26976 22374 27028 22380
rect 27344 22374 27396 22380
rect 26988 22234 27016 22374
rect 27448 22234 27476 22442
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 26988 21554 27016 22170
rect 27908 22098 27936 23054
rect 28080 22568 28132 22574
rect 28080 22510 28132 22516
rect 28092 22234 28120 22510
rect 28080 22228 28132 22234
rect 28080 22170 28132 22176
rect 27896 22092 27948 22098
rect 27896 22034 27948 22040
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 26884 21140 26936 21146
rect 26884 21082 26936 21088
rect 26988 20942 27016 21490
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26804 19446 26832 20198
rect 26884 19712 26936 19718
rect 26884 19654 26936 19660
rect 27080 19666 27108 20946
rect 27264 20466 27292 21286
rect 27816 20942 27844 21490
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27620 20868 27672 20874
rect 27620 20810 27672 20816
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27160 19712 27212 19718
rect 27080 19660 27160 19666
rect 27080 19654 27212 19660
rect 26792 19440 26844 19446
rect 26792 19382 26844 19388
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26332 19236 26384 19242
rect 26332 19178 26384 19184
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 26896 18766 26924 19654
rect 27080 19638 27200 19654
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 27080 19310 27108 19450
rect 27172 19378 27200 19638
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 27080 18902 27108 19246
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 27264 18834 27292 20402
rect 27540 19378 27568 20538
rect 27632 20466 27660 20810
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27816 20398 27844 20878
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 27816 19854 27844 20334
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 27528 19372 27580 19378
rect 27528 19314 27580 19320
rect 27632 19310 27660 19790
rect 27712 19780 27764 19786
rect 27712 19722 27764 19728
rect 27620 19304 27672 19310
rect 27620 19246 27672 19252
rect 27724 18970 27752 19722
rect 27908 19378 27936 22034
rect 28368 21894 28396 23054
rect 28540 23054 28592 23060
rect 28446 23015 28502 23024
rect 28552 22710 28580 23054
rect 28828 22778 28856 24006
rect 28920 23730 28948 24006
rect 29012 23866 29040 24618
rect 29564 24410 29592 24686
rect 29552 24404 29604 24410
rect 29552 24346 29604 24352
rect 29460 24268 29512 24274
rect 29460 24210 29512 24216
rect 29368 24132 29420 24138
rect 29368 24074 29420 24080
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 29380 23730 29408 24074
rect 29472 23730 29500 24210
rect 28908 23724 28960 23730
rect 29276 23724 29328 23730
rect 28908 23666 28960 23672
rect 29196 23684 29276 23712
rect 28816 22772 28868 22778
rect 28816 22714 28868 22720
rect 28540 22704 28592 22710
rect 28540 22646 28592 22652
rect 28920 22642 28948 23666
rect 29196 22710 29224 23684
rect 29276 23666 29328 23672
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29460 23724 29512 23730
rect 29460 23666 29512 23672
rect 29380 22778 29408 23666
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29184 22704 29236 22710
rect 29184 22646 29236 22652
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 28644 22234 28672 22578
rect 28816 22500 28868 22506
rect 28816 22442 28868 22448
rect 28632 22228 28684 22234
rect 28632 22170 28684 22176
rect 28828 22098 28856 22442
rect 28816 22092 28868 22098
rect 28816 22034 28868 22040
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 28368 21690 28396 21830
rect 28356 21684 28408 21690
rect 28356 21626 28408 21632
rect 28460 21486 28488 21966
rect 28644 21554 28672 21966
rect 28816 21956 28868 21962
rect 28816 21898 28868 21904
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28080 21072 28132 21078
rect 28080 21014 28132 21020
rect 28092 20058 28120 21014
rect 28080 20052 28132 20058
rect 28080 19994 28132 20000
rect 27988 19712 28040 19718
rect 27988 19654 28040 19660
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27804 19168 27856 19174
rect 27804 19110 27856 19116
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27816 18834 27844 19110
rect 27252 18828 27304 18834
rect 27252 18770 27304 18776
rect 27804 18828 27856 18834
rect 27804 18770 27856 18776
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26988 18340 27016 18634
rect 26896 18312 27016 18340
rect 27252 18352 27304 18358
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26160 17678 26188 18226
rect 26792 17808 26844 17814
rect 26792 17750 26844 17756
rect 26804 17678 26832 17750
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 26068 16726 26096 17070
rect 26160 17066 26188 17614
rect 26620 17338 26648 17614
rect 26896 17542 26924 18312
rect 27356 18340 27384 18702
rect 27712 18692 27764 18698
rect 27712 18634 27764 18640
rect 27304 18312 27384 18340
rect 27252 18294 27304 18300
rect 27264 17882 27292 18294
rect 27724 18222 27752 18634
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 27816 17678 27844 18770
rect 27908 18766 27936 19314
rect 27896 18760 27948 18766
rect 27896 18702 27948 18708
rect 28000 17882 28028 19654
rect 28184 19446 28212 21082
rect 28828 20942 28856 21898
rect 28920 21690 28948 22578
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 28920 20942 28948 21626
rect 29012 21418 29040 22510
rect 29196 22438 29224 22646
rect 29184 22432 29236 22438
rect 29184 22374 29236 22380
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 29000 21412 29052 21418
rect 29000 21354 29052 21360
rect 29012 21078 29040 21354
rect 29184 21344 29236 21350
rect 29184 21286 29236 21292
rect 29000 21072 29052 21078
rect 29000 21014 29052 21020
rect 29196 20942 29224 21286
rect 29288 21078 29316 21490
rect 29380 21146 29408 22714
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29460 21956 29512 21962
rect 29460 21898 29512 21904
rect 29472 21554 29500 21898
rect 29656 21554 29684 21966
rect 29460 21548 29512 21554
rect 29460 21490 29512 21496
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29276 21072 29328 21078
rect 29276 21014 29328 21020
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 29184 20936 29236 20942
rect 29184 20878 29236 20884
rect 28368 20398 28396 20878
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 28080 19236 28132 19242
rect 28080 19178 28132 19184
rect 28092 18766 28120 19178
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 28092 18170 28120 18702
rect 28184 18290 28212 19382
rect 28460 18766 28488 20742
rect 29012 20466 29040 20878
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29012 19854 29040 20402
rect 29196 20058 29224 20878
rect 29288 20534 29316 21014
rect 29276 20528 29328 20534
rect 29276 20470 29328 20476
rect 29380 20466 29408 21082
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29368 19916 29420 19922
rect 29472 19904 29500 20878
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29564 19922 29592 20402
rect 29656 20262 29684 21490
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29644 20256 29696 20262
rect 29644 20198 29696 20204
rect 29656 20058 29684 20198
rect 29644 20052 29696 20058
rect 29644 19994 29696 20000
rect 29420 19876 29500 19904
rect 29552 19916 29604 19922
rect 29368 19858 29420 19864
rect 29552 19858 29604 19864
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28828 19174 28856 19790
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 28816 19168 28868 19174
rect 28816 19110 28868 19116
rect 29012 18766 29040 19450
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 29104 18970 29132 19314
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29380 19258 29408 19858
rect 29656 19854 29684 19994
rect 29748 19854 29776 20334
rect 29840 19990 29868 25094
rect 29932 21622 29960 25452
rect 30300 25362 30328 25978
rect 30288 25356 30340 25362
rect 30288 25298 30340 25304
rect 30760 25226 30788 26726
rect 31036 26382 31064 26930
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 30932 26240 30984 26246
rect 30932 26182 30984 26188
rect 30944 25294 30972 26182
rect 31128 25906 31156 27474
rect 31496 27470 31524 27814
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31208 27056 31260 27062
rect 31208 26998 31260 27004
rect 31220 26518 31248 26998
rect 31208 26512 31260 26518
rect 31208 26454 31260 26460
rect 31220 26382 31248 26454
rect 31208 26376 31260 26382
rect 31208 26318 31260 26324
rect 31680 26314 31708 28698
rect 31864 28218 31892 28902
rect 31852 28212 31904 28218
rect 31852 28154 31904 28160
rect 31760 27668 31812 27674
rect 31760 27610 31812 27616
rect 31772 26926 31800 27610
rect 31864 27538 31892 28154
rect 32140 27606 32168 29582
rect 32876 29306 32904 30670
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 32968 29850 32996 30194
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 33244 29646 33272 30670
rect 33336 30326 33364 30874
rect 33520 30802 33548 31282
rect 33888 30938 33916 32370
rect 34348 32314 34376 32982
rect 34532 32774 34560 33322
rect 34796 33312 34848 33318
rect 34796 33254 34848 33260
rect 34808 32978 34836 33254
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35544 33114 35572 33526
rect 38474 33416 38530 33425
rect 38474 33351 38476 33360
rect 38528 33351 38530 33360
rect 38476 33322 38528 33328
rect 35532 33108 35584 33114
rect 35532 33050 35584 33056
rect 35544 32978 35572 33050
rect 34796 32972 34848 32978
rect 34796 32914 34848 32920
rect 35532 32972 35584 32978
rect 35532 32914 35584 32920
rect 34612 32904 34664 32910
rect 34612 32846 34664 32852
rect 34520 32768 34572 32774
rect 34520 32710 34572 32716
rect 34624 32570 34652 32846
rect 36176 32836 36228 32842
rect 36176 32778 36228 32784
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 34612 32564 34664 32570
rect 34612 32506 34664 32512
rect 34612 32360 34664 32366
rect 34348 32308 34612 32314
rect 34348 32302 34664 32308
rect 34348 32286 34652 32302
rect 34348 31754 34376 32286
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34348 31726 34468 31754
rect 34440 31278 34468 31726
rect 34612 31408 34664 31414
rect 34612 31350 34664 31356
rect 34428 31272 34480 31278
rect 34428 31214 34480 31220
rect 33876 30932 33928 30938
rect 33876 30874 33928 30880
rect 34244 30932 34296 30938
rect 34244 30874 34296 30880
rect 33508 30796 33560 30802
rect 33508 30738 33560 30744
rect 33968 30796 34020 30802
rect 33968 30738 34020 30744
rect 33692 30728 33744 30734
rect 33692 30670 33744 30676
rect 33324 30320 33376 30326
rect 33324 30262 33376 30268
rect 33508 29844 33560 29850
rect 33508 29786 33560 29792
rect 33048 29640 33100 29646
rect 33048 29582 33100 29588
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 32864 29300 32916 29306
rect 32864 29242 32916 29248
rect 32772 29164 32824 29170
rect 32772 29106 32824 29112
rect 32784 28490 32812 29106
rect 33060 29102 33088 29582
rect 33140 29232 33192 29238
rect 33140 29174 33192 29180
rect 33048 29096 33100 29102
rect 33048 29038 33100 29044
rect 33152 28966 33180 29174
rect 33140 28960 33192 28966
rect 33140 28902 33192 28908
rect 33520 28626 33548 29786
rect 33704 29646 33732 30670
rect 33980 30598 34008 30738
rect 34256 30734 34284 30874
rect 34440 30802 34468 31214
rect 34428 30796 34480 30802
rect 34428 30738 34480 30744
rect 34244 30728 34296 30734
rect 34440 30682 34468 30738
rect 34244 30670 34296 30676
rect 33968 30592 34020 30598
rect 33968 30534 34020 30540
rect 33876 30252 33928 30258
rect 33980 30240 34008 30534
rect 34256 30394 34284 30670
rect 34348 30654 34468 30682
rect 34244 30388 34296 30394
rect 34244 30330 34296 30336
rect 33928 30212 34008 30240
rect 33876 30194 33928 30200
rect 33888 29646 33916 30194
rect 34348 29850 34376 30654
rect 34520 30592 34572 30598
rect 34520 30534 34572 30540
rect 34532 30326 34560 30534
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 34428 30184 34480 30190
rect 34428 30126 34480 30132
rect 34336 29844 34388 29850
rect 34336 29786 34388 29792
rect 33692 29640 33744 29646
rect 33692 29582 33744 29588
rect 33876 29640 33928 29646
rect 33876 29582 33928 29588
rect 33888 29306 33916 29582
rect 34152 29504 34204 29510
rect 34152 29446 34204 29452
rect 34336 29504 34388 29510
rect 34336 29446 34388 29452
rect 33876 29300 33928 29306
rect 33876 29242 33928 29248
rect 34164 29238 34192 29446
rect 34348 29306 34376 29446
rect 34336 29300 34388 29306
rect 34336 29242 34388 29248
rect 33600 29232 33652 29238
rect 33600 29174 33652 29180
rect 34152 29232 34204 29238
rect 34152 29174 34204 29180
rect 33508 28620 33560 28626
rect 33508 28562 33560 28568
rect 33140 28552 33192 28558
rect 33140 28494 33192 28500
rect 32772 28484 32824 28490
rect 32772 28426 32824 28432
rect 32784 28014 32812 28426
rect 33048 28416 33100 28422
rect 33048 28358 33100 28364
rect 32956 28144 33008 28150
rect 32956 28086 33008 28092
rect 32772 28008 32824 28014
rect 32772 27950 32824 27956
rect 32680 27872 32732 27878
rect 32680 27814 32732 27820
rect 32128 27600 32180 27606
rect 32128 27542 32180 27548
rect 31852 27532 31904 27538
rect 31852 27474 31904 27480
rect 32140 27062 32168 27542
rect 32404 27396 32456 27402
rect 32404 27338 32456 27344
rect 32128 27056 32180 27062
rect 32128 26998 32180 27004
rect 31760 26920 31812 26926
rect 31760 26862 31812 26868
rect 31668 26308 31720 26314
rect 31668 26250 31720 26256
rect 31680 26042 31708 26250
rect 31668 26036 31720 26042
rect 31668 25978 31720 25984
rect 32416 25974 32444 27338
rect 32692 26994 32720 27814
rect 32784 27538 32812 27950
rect 32772 27532 32824 27538
rect 32772 27474 32824 27480
rect 32968 27334 32996 28086
rect 33060 27470 33088 28358
rect 33152 27606 33180 28494
rect 33612 28490 33640 29174
rect 34060 29096 34112 29102
rect 34060 29038 34112 29044
rect 34072 28966 34100 29038
rect 34060 28960 34112 28966
rect 34060 28902 34112 28908
rect 34072 28694 34100 28902
rect 33968 28688 34020 28694
rect 33968 28630 34020 28636
rect 34060 28688 34112 28694
rect 34060 28630 34112 28636
rect 33980 28558 34008 28630
rect 34164 28558 34192 29174
rect 34440 29170 34468 30126
rect 34624 30122 34652 31350
rect 34716 30258 34744 31758
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 36188 31414 36216 32778
rect 36728 32768 36780 32774
rect 36728 32710 36780 32716
rect 36740 32434 36768 32710
rect 36728 32428 36780 32434
rect 36728 32370 36780 32376
rect 36636 31816 36688 31822
rect 36636 31758 36688 31764
rect 36648 31482 36676 31758
rect 36636 31476 36688 31482
rect 36636 31418 36688 31424
rect 36176 31408 36228 31414
rect 36096 31356 36176 31362
rect 36096 31350 36228 31356
rect 36096 31334 36216 31350
rect 35348 31136 35400 31142
rect 35348 31078 35400 31084
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30734 35388 31078
rect 35992 30796 36044 30802
rect 35992 30738 36044 30744
rect 35348 30728 35400 30734
rect 35348 30670 35400 30676
rect 35072 30592 35124 30598
rect 35072 30534 35124 30540
rect 35084 30394 35112 30534
rect 35072 30388 35124 30394
rect 35072 30330 35124 30336
rect 35360 30258 35388 30670
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 34704 30252 34756 30258
rect 34704 30194 34756 30200
rect 35348 30252 35400 30258
rect 35348 30194 35400 30200
rect 35440 30252 35492 30258
rect 35440 30194 35492 30200
rect 34612 30116 34664 30122
rect 34612 30058 34664 30064
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35360 29714 35388 30194
rect 35452 29850 35480 30194
rect 36004 30190 36032 30738
rect 36096 30666 36124 31334
rect 36084 30660 36136 30666
rect 36084 30602 36136 30608
rect 35992 30184 36044 30190
rect 35992 30126 36044 30132
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 35348 29708 35400 29714
rect 35348 29650 35400 29656
rect 34428 29164 34480 29170
rect 34428 29106 34480 29112
rect 34612 29164 34664 29170
rect 34612 29106 34664 29112
rect 34336 29028 34388 29034
rect 34336 28970 34388 28976
rect 34348 28626 34376 28970
rect 34624 28762 34652 29106
rect 35360 29084 35388 29650
rect 35452 29186 35480 29786
rect 36096 29646 36124 30602
rect 36648 30258 36676 31418
rect 36636 30252 36688 30258
rect 36636 30194 36688 30200
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 36452 29504 36504 29510
rect 36452 29446 36504 29452
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 35992 29232 36044 29238
rect 35452 29158 35572 29186
rect 35992 29174 36044 29180
rect 35440 29096 35492 29102
rect 35360 29056 35440 29084
rect 35440 29038 35492 29044
rect 34796 28960 34848 28966
rect 34796 28902 34848 28908
rect 34612 28756 34664 28762
rect 34612 28698 34664 28704
rect 34336 28620 34388 28626
rect 34336 28562 34388 28568
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33968 28552 34020 28558
rect 33968 28494 34020 28500
rect 34152 28552 34204 28558
rect 34152 28494 34204 28500
rect 33600 28484 33652 28490
rect 33600 28426 33652 28432
rect 33692 28416 33744 28422
rect 33692 28358 33744 28364
rect 33704 28150 33732 28358
rect 33692 28144 33744 28150
rect 33692 28086 33744 28092
rect 33140 27600 33192 27606
rect 33140 27542 33192 27548
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 32956 27328 33008 27334
rect 32956 27270 33008 27276
rect 32968 27062 32996 27270
rect 33796 27130 33824 28494
rect 34336 28484 34388 28490
rect 34336 28426 34388 28432
rect 34348 28082 34376 28426
rect 34808 28422 34836 28902
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34888 28756 34940 28762
rect 34888 28698 34940 28704
rect 34900 28626 34928 28698
rect 34888 28620 34940 28626
rect 34888 28562 34940 28568
rect 35348 28552 35400 28558
rect 35268 28500 35348 28506
rect 35268 28494 35400 28500
rect 35268 28478 35388 28494
rect 34796 28416 34848 28422
rect 34796 28358 34848 28364
rect 34808 28218 34836 28358
rect 34796 28212 34848 28218
rect 34796 28154 34848 28160
rect 34336 28076 34388 28082
rect 34336 28018 34388 28024
rect 33968 28008 34020 28014
rect 33968 27950 34020 27956
rect 33980 27674 34008 27950
rect 34520 27872 34572 27878
rect 34520 27814 34572 27820
rect 33968 27668 34020 27674
rect 33968 27610 34020 27616
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 32956 27056 33008 27062
rect 32956 26998 33008 27004
rect 32680 26988 32732 26994
rect 32680 26930 32732 26936
rect 32692 26314 32720 26930
rect 33600 26784 33652 26790
rect 33600 26726 33652 26732
rect 32680 26308 32732 26314
rect 32680 26250 32732 26256
rect 32404 25968 32456 25974
rect 32404 25910 32456 25916
rect 33612 25906 33640 26726
rect 33796 26382 33824 27066
rect 34532 26926 34560 27814
rect 34808 27656 34836 28154
rect 35268 27946 35296 28478
rect 35348 28416 35400 28422
rect 35348 28358 35400 28364
rect 35256 27940 35308 27946
rect 35256 27882 35308 27888
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34808 27628 34928 27656
rect 34796 27328 34848 27334
rect 34796 27270 34848 27276
rect 34520 26920 34572 26926
rect 34520 26862 34572 26868
rect 33784 26376 33836 26382
rect 33784 26318 33836 26324
rect 34808 25974 34836 27270
rect 34900 27130 34928 27628
rect 35360 27606 35388 28358
rect 35452 28014 35480 29038
rect 35544 28694 35572 29158
rect 36004 28762 36032 29174
rect 35992 28756 36044 28762
rect 35992 28698 36044 28704
rect 35532 28688 35584 28694
rect 35532 28630 35584 28636
rect 36464 28626 36492 29446
rect 36648 29306 36676 30194
rect 36740 29646 36768 32370
rect 38476 31816 38528 31822
rect 38476 31758 38528 31764
rect 38488 31385 38516 31758
rect 38474 31376 38530 31385
rect 38474 31311 38530 31320
rect 38476 30728 38528 30734
rect 38474 30696 38476 30705
rect 38528 30696 38530 30705
rect 38474 30631 38530 30640
rect 37188 30592 37240 30598
rect 37188 30534 37240 30540
rect 37200 30190 37228 30534
rect 37188 30184 37240 30190
rect 37188 30126 37240 30132
rect 36728 29640 36780 29646
rect 36728 29582 36780 29588
rect 36820 29640 36872 29646
rect 36820 29582 36872 29588
rect 36636 29300 36688 29306
rect 36636 29242 36688 29248
rect 36648 29170 36676 29242
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 36832 28966 36860 29582
rect 37200 29510 37228 30126
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37280 29776 37332 29782
rect 37280 29718 37332 29724
rect 37188 29504 37240 29510
rect 37188 29446 37240 29452
rect 37200 29170 37228 29446
rect 37188 29164 37240 29170
rect 37188 29106 37240 29112
rect 36820 28960 36872 28966
rect 36820 28902 36872 28908
rect 37004 28960 37056 28966
rect 37004 28902 37056 28908
rect 36832 28626 36860 28902
rect 36452 28620 36504 28626
rect 36452 28562 36504 28568
rect 36820 28620 36872 28626
rect 36820 28562 36872 28568
rect 37016 28558 37044 28902
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 36176 28552 36228 28558
rect 36176 28494 36228 28500
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 37004 28552 37056 28558
rect 37004 28494 37056 28500
rect 35544 28422 35572 28494
rect 36188 28422 36216 28494
rect 35532 28416 35584 28422
rect 35532 28358 35584 28364
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 36372 28218 36400 28494
rect 36360 28212 36412 28218
rect 36360 28154 36412 28160
rect 37292 28082 37320 29718
rect 37476 28558 37504 29990
rect 37648 28960 37700 28966
rect 37648 28902 37700 28908
rect 37464 28552 37516 28558
rect 37464 28494 37516 28500
rect 37556 28484 37608 28490
rect 37556 28426 37608 28432
rect 37568 28150 37596 28426
rect 37660 28150 37688 28902
rect 37740 28552 37792 28558
rect 37740 28494 37792 28500
rect 37924 28552 37976 28558
rect 37924 28494 37976 28500
rect 37752 28218 37780 28494
rect 37740 28212 37792 28218
rect 37740 28154 37792 28160
rect 37556 28144 37608 28150
rect 37556 28086 37608 28092
rect 37648 28144 37700 28150
rect 37648 28086 37700 28092
rect 37280 28076 37332 28082
rect 37280 28018 37332 28024
rect 35440 28008 35492 28014
rect 35440 27950 35492 27956
rect 35348 27600 35400 27606
rect 35348 27542 35400 27548
rect 35256 27464 35308 27470
rect 35256 27406 35308 27412
rect 34888 27124 34940 27130
rect 34888 27066 34940 27072
rect 35268 27062 35296 27406
rect 35348 27328 35400 27334
rect 35348 27270 35400 27276
rect 35256 27056 35308 27062
rect 35256 26998 35308 27004
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26586 35388 27270
rect 35452 26994 35480 27950
rect 37568 27606 37596 28086
rect 37556 27600 37608 27606
rect 37556 27542 37608 27548
rect 37372 27464 37424 27470
rect 37660 27452 37688 28086
rect 37740 28076 37792 28082
rect 37740 28018 37792 28024
rect 37752 27674 37780 28018
rect 37936 27674 37964 28494
rect 38016 28416 38068 28422
rect 38016 28358 38068 28364
rect 38028 28082 38056 28358
rect 38016 28076 38068 28082
rect 38016 28018 38068 28024
rect 38016 27940 38068 27946
rect 38016 27882 38068 27888
rect 37740 27668 37792 27674
rect 37740 27610 37792 27616
rect 37924 27668 37976 27674
rect 37924 27610 37976 27616
rect 37424 27424 37688 27452
rect 37372 27406 37424 27412
rect 37464 27328 37516 27334
rect 37464 27270 37516 27276
rect 37556 27328 37608 27334
rect 37556 27270 37608 27276
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 36544 26988 36596 26994
rect 36544 26930 36596 26936
rect 36728 26988 36780 26994
rect 36728 26930 36780 26936
rect 35624 26920 35676 26926
rect 35624 26862 35676 26868
rect 36176 26920 36228 26926
rect 36176 26862 36228 26868
rect 35636 26586 35664 26862
rect 35348 26580 35400 26586
rect 35348 26522 35400 26528
rect 35624 26580 35676 26586
rect 35624 26522 35676 26528
rect 36188 26382 36216 26862
rect 36556 26586 36584 26930
rect 36544 26580 36596 26586
rect 36544 26522 36596 26528
rect 36740 26382 36768 26930
rect 37476 26926 37504 27270
rect 37372 26920 37424 26926
rect 37372 26862 37424 26868
rect 37464 26920 37516 26926
rect 37464 26862 37516 26868
rect 37384 26518 37412 26862
rect 37568 26858 37596 27270
rect 37660 26994 37688 27424
rect 37648 26988 37700 26994
rect 37648 26930 37700 26936
rect 37556 26852 37608 26858
rect 37556 26794 37608 26800
rect 37464 26784 37516 26790
rect 37464 26726 37516 26732
rect 37372 26512 37424 26518
rect 37372 26454 37424 26460
rect 37476 26450 37504 26726
rect 37464 26444 37516 26450
rect 37464 26386 37516 26392
rect 35992 26376 36044 26382
rect 35992 26318 36044 26324
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 36176 26376 36228 26382
rect 36176 26318 36228 26324
rect 36728 26376 36780 26382
rect 36728 26318 36780 26324
rect 37372 26376 37424 26382
rect 37372 26318 37424 26324
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 36004 26042 36032 26318
rect 36096 26042 36124 26318
rect 35992 26036 36044 26042
rect 35992 25978 36044 25984
rect 36084 26036 36136 26042
rect 36084 25978 36136 25984
rect 34796 25968 34848 25974
rect 34796 25910 34848 25916
rect 31116 25900 31168 25906
rect 31116 25842 31168 25848
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 32312 25900 32364 25906
rect 32312 25842 32364 25848
rect 32956 25900 33008 25906
rect 32956 25842 33008 25848
rect 33600 25900 33652 25906
rect 33600 25842 33652 25848
rect 34336 25900 34388 25906
rect 34336 25842 34388 25848
rect 35440 25900 35492 25906
rect 35440 25842 35492 25848
rect 31588 25362 31616 25842
rect 32324 25498 32352 25842
rect 32312 25492 32364 25498
rect 32312 25434 32364 25440
rect 31576 25356 31628 25362
rect 31576 25298 31628 25304
rect 30932 25288 30984 25294
rect 30852 25248 30932 25276
rect 30748 25220 30800 25226
rect 30748 25162 30800 25168
rect 30760 24954 30788 25162
rect 30748 24948 30800 24954
rect 30748 24890 30800 24896
rect 30852 24818 30880 25248
rect 30932 25230 30984 25236
rect 31208 25288 31260 25294
rect 31208 25230 31260 25236
rect 32220 25288 32272 25294
rect 32220 25230 32272 25236
rect 32680 25288 32732 25294
rect 32680 25230 32732 25236
rect 31116 25220 31168 25226
rect 31116 25162 31168 25168
rect 31128 24818 31156 25162
rect 31220 24954 31248 25230
rect 32128 25220 32180 25226
rect 32128 25162 32180 25168
rect 31208 24948 31260 24954
rect 31208 24890 31260 24896
rect 31576 24880 31628 24886
rect 31576 24822 31628 24828
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31588 24750 31616 24822
rect 32140 24818 32168 25162
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 31576 24744 31628 24750
rect 31576 24686 31628 24692
rect 31588 24410 31616 24686
rect 32140 24614 32168 24754
rect 32232 24682 32260 25230
rect 32588 25220 32640 25226
rect 32588 25162 32640 25168
rect 32600 24954 32628 25162
rect 32692 24954 32720 25230
rect 32968 25158 32996 25842
rect 33140 25832 33192 25838
rect 33140 25774 33192 25780
rect 33152 25702 33180 25774
rect 33140 25696 33192 25702
rect 33140 25638 33192 25644
rect 33152 25498 33180 25638
rect 34348 25498 34376 25842
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 33140 25492 33192 25498
rect 33140 25434 33192 25440
rect 34336 25492 34388 25498
rect 34336 25434 34388 25440
rect 33416 25288 33468 25294
rect 33416 25230 33468 25236
rect 33600 25288 33652 25294
rect 33600 25230 33652 25236
rect 32956 25152 33008 25158
rect 32956 25094 33008 25100
rect 33428 24954 33456 25230
rect 32588 24948 32640 24954
rect 32588 24890 32640 24896
rect 32680 24948 32732 24954
rect 32680 24890 32732 24896
rect 33416 24948 33468 24954
rect 33416 24890 33468 24896
rect 33612 24886 33640 25230
rect 34704 25220 34756 25226
rect 34704 25162 34756 25168
rect 34888 25220 34940 25226
rect 34888 25162 34940 25168
rect 34716 24954 34744 25162
rect 34704 24948 34756 24954
rect 34704 24890 34756 24896
rect 33600 24880 33652 24886
rect 33600 24822 33652 24828
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 34796 24812 34848 24818
rect 34796 24754 34848 24760
rect 32220 24676 32272 24682
rect 32220 24618 32272 24624
rect 32312 24676 32364 24682
rect 32312 24618 32364 24624
rect 32128 24608 32180 24614
rect 32128 24550 32180 24556
rect 31576 24404 31628 24410
rect 31576 24346 31628 24352
rect 32324 24206 32352 24618
rect 32692 24410 32720 24754
rect 33796 24698 33824 24754
rect 33704 24682 33824 24698
rect 33692 24676 33824 24682
rect 33744 24670 33824 24676
rect 33876 24676 33928 24682
rect 33692 24618 33744 24624
rect 33876 24618 33928 24624
rect 32680 24404 32732 24410
rect 32680 24346 32732 24352
rect 33704 24274 33732 24618
rect 33784 24608 33836 24614
rect 33784 24550 33836 24556
rect 33692 24268 33744 24274
rect 33692 24210 33744 24216
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 30012 24064 30064 24070
rect 30012 24006 30064 24012
rect 30024 23798 30052 24006
rect 30208 23866 30236 24142
rect 30196 23860 30248 23866
rect 30196 23802 30248 23808
rect 30392 23798 30420 24142
rect 31576 24132 31628 24138
rect 31576 24074 31628 24080
rect 31588 23866 31616 24074
rect 32876 23866 32904 24142
rect 33704 23866 33732 24210
rect 33796 24206 33824 24550
rect 33888 24410 33916 24618
rect 33876 24404 33928 24410
rect 33876 24346 33928 24352
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 33796 23866 33824 24142
rect 34532 23866 34560 24142
rect 34808 23866 34836 24754
rect 34900 24682 34928 25162
rect 35452 24954 35480 25842
rect 35992 25764 36044 25770
rect 35992 25706 36044 25712
rect 36004 25430 36032 25706
rect 36740 25498 36768 26318
rect 36728 25492 36780 25498
rect 36728 25434 36780 25440
rect 35992 25424 36044 25430
rect 35992 25366 36044 25372
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 36004 24954 36032 25366
rect 37096 25356 37148 25362
rect 37096 25298 37148 25304
rect 36912 25288 36964 25294
rect 36832 25236 36912 25242
rect 36832 25230 36964 25236
rect 36832 25214 36952 25230
rect 35440 24948 35492 24954
rect 35440 24890 35492 24896
rect 35992 24948 36044 24954
rect 35992 24890 36044 24896
rect 36832 24818 36860 25214
rect 37108 25158 37136 25298
rect 37004 25152 37056 25158
rect 37004 25094 37056 25100
rect 37096 25152 37148 25158
rect 37096 25094 37148 25100
rect 37016 24818 37044 25094
rect 35440 24812 35492 24818
rect 35440 24754 35492 24760
rect 36820 24812 36872 24818
rect 36820 24754 36872 24760
rect 37004 24812 37056 24818
rect 37004 24754 37056 24760
rect 34888 24676 34940 24682
rect 34888 24618 34940 24624
rect 35452 24614 35480 24754
rect 35532 24744 35584 24750
rect 35532 24686 35584 24692
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 32864 23860 32916 23866
rect 32864 23802 32916 23808
rect 33692 23860 33744 23866
rect 33692 23802 33744 23808
rect 33784 23860 33836 23866
rect 33784 23802 33836 23808
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 30012 23792 30064 23798
rect 30012 23734 30064 23740
rect 30380 23792 30432 23798
rect 30380 23734 30432 23740
rect 33048 23792 33100 23798
rect 33048 23734 33100 23740
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 32128 23724 32180 23730
rect 32128 23666 32180 23672
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 30010 23488 30066 23497
rect 30010 23423 30066 23432
rect 29920 21616 29972 21622
rect 29920 21558 29972 21564
rect 29828 19984 29880 19990
rect 29828 19926 29880 19932
rect 30024 19922 30052 23423
rect 30116 23254 30144 23598
rect 30104 23248 30156 23254
rect 30104 23190 30156 23196
rect 30208 22778 30236 23666
rect 31588 23322 31616 23666
rect 32140 23322 32168 23666
rect 33060 23322 33088 23734
rect 35452 23730 35480 24550
rect 35544 24410 35572 24686
rect 35532 24404 35584 24410
rect 35532 24346 35584 24352
rect 36832 24342 36860 24754
rect 37016 24410 37044 24754
rect 37108 24682 37136 25094
rect 37096 24676 37148 24682
rect 37096 24618 37148 24624
rect 37004 24404 37056 24410
rect 37004 24346 37056 24352
rect 36176 24336 36228 24342
rect 36176 24278 36228 24284
rect 36820 24336 36872 24342
rect 36820 24278 36872 24284
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 34336 23724 34388 23730
rect 34336 23666 34388 23672
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 31576 23316 31628 23322
rect 31576 23258 31628 23264
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30300 22778 30328 23122
rect 30840 23112 30892 23118
rect 30840 23054 30892 23060
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 30852 22778 30880 23054
rect 30196 22772 30248 22778
rect 30196 22714 30248 22720
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30104 22568 30156 22574
rect 30104 22510 30156 22516
rect 30116 22234 30144 22510
rect 30104 22228 30156 22234
rect 30104 22170 30156 22176
rect 30196 22092 30248 22098
rect 30196 22034 30248 22040
rect 30208 21554 30236 22034
rect 30196 21548 30248 21554
rect 30196 21490 30248 21496
rect 30392 21350 30420 22578
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30392 20942 30420 21286
rect 30852 21010 30880 22714
rect 31772 22506 31800 23054
rect 32140 22778 32168 23054
rect 32128 22772 32180 22778
rect 32128 22714 32180 22720
rect 33048 22704 33100 22710
rect 33048 22646 33100 22652
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 32036 22568 32088 22574
rect 32036 22510 32088 22516
rect 31760 22500 31812 22506
rect 31760 22442 31812 22448
rect 32048 22234 32076 22510
rect 32324 22234 32352 22578
rect 32876 22438 32904 22578
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32036 22228 32088 22234
rect 32036 22170 32088 22176
rect 32312 22228 32364 22234
rect 32312 22170 32364 22176
rect 32876 22030 32904 22374
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 31760 21480 31812 21486
rect 31760 21422 31812 21428
rect 31772 21146 31800 21422
rect 31760 21140 31812 21146
rect 31760 21082 31812 21088
rect 30840 21004 30892 21010
rect 30840 20946 30892 20952
rect 32324 20942 32352 21490
rect 32692 21486 32720 21966
rect 33060 21962 33088 22646
rect 33152 22234 33180 23054
rect 33244 22778 33272 23054
rect 34348 22778 34376 23666
rect 34624 22778 34652 23666
rect 34808 22778 34836 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 33232 22772 33284 22778
rect 33232 22714 33284 22720
rect 34336 22772 34388 22778
rect 34336 22714 34388 22720
rect 34612 22772 34664 22778
rect 34612 22714 34664 22720
rect 34796 22772 34848 22778
rect 34796 22714 34848 22720
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 33968 22568 34020 22574
rect 33968 22510 34020 22516
rect 33140 22228 33192 22234
rect 33140 22170 33192 22176
rect 33048 21956 33100 21962
rect 33048 21898 33100 21904
rect 32680 21480 32732 21486
rect 32680 21422 32732 21428
rect 33060 21146 33088 21898
rect 33980 21690 34008 22510
rect 34440 22234 34468 22578
rect 34624 22234 34652 22578
rect 35360 22438 35388 22578
rect 35452 22506 35480 23666
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35900 22636 35952 22642
rect 35900 22578 35952 22584
rect 35440 22500 35492 22506
rect 35440 22442 35492 22448
rect 35348 22432 35400 22438
rect 35348 22374 35400 22380
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34428 22228 34480 22234
rect 34428 22170 34480 22176
rect 34612 22228 34664 22234
rect 34612 22170 34664 22176
rect 35256 22094 35308 22098
rect 35360 22094 35388 22374
rect 35256 22092 35388 22094
rect 35308 22066 35388 22092
rect 35912 22094 35940 22578
rect 35912 22066 36032 22094
rect 35256 22034 35308 22040
rect 34428 22024 34480 22030
rect 34428 21966 34480 21972
rect 33968 21684 34020 21690
rect 33968 21626 34020 21632
rect 34336 21616 34388 21622
rect 34336 21558 34388 21564
rect 33876 21548 33928 21554
rect 33876 21490 33928 21496
rect 33888 21146 33916 21490
rect 34348 21146 34376 21558
rect 33048 21140 33100 21146
rect 33048 21082 33100 21088
rect 33876 21140 33928 21146
rect 33876 21082 33928 21088
rect 34336 21140 34388 21146
rect 34336 21082 34388 21088
rect 30380 20936 30432 20942
rect 31392 20936 31444 20942
rect 30380 20878 30432 20884
rect 31390 20904 31392 20913
rect 31576 20936 31628 20942
rect 31444 20904 31446 20913
rect 31576 20878 31628 20884
rect 32312 20936 32364 20942
rect 33876 20936 33928 20942
rect 32312 20878 32364 20884
rect 33046 20904 33102 20913
rect 31390 20839 31446 20848
rect 31588 20806 31616 20878
rect 31944 20868 31996 20874
rect 31944 20810 31996 20816
rect 32588 20868 32640 20874
rect 33876 20878 33928 20884
rect 33046 20839 33048 20848
rect 32588 20810 32640 20816
rect 33100 20839 33102 20848
rect 33048 20810 33100 20816
rect 30196 20800 30248 20806
rect 30196 20742 30248 20748
rect 31576 20800 31628 20806
rect 31576 20742 31628 20748
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 30012 19916 30064 19922
rect 30012 19858 30064 19864
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29460 19780 29512 19786
rect 29460 19722 29512 19728
rect 29472 19378 29500 19722
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 29092 18964 29144 18970
rect 29092 18906 29144 18912
rect 29196 18766 29224 19110
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 28276 18426 28304 18702
rect 28264 18420 28316 18426
rect 28264 18362 28316 18368
rect 28276 18290 28304 18362
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28460 18222 28488 18702
rect 28828 18426 28856 18702
rect 29092 18692 29144 18698
rect 29092 18634 29144 18640
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28448 18216 28500 18222
rect 28092 18142 28304 18170
rect 28448 18158 28500 18164
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 28000 17678 28028 17818
rect 28276 17814 28304 18142
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28264 17808 28316 17814
rect 28264 17750 28316 17756
rect 28276 17678 28304 17750
rect 28736 17678 28764 18022
rect 28920 17678 28948 18566
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 29012 17678 29040 18226
rect 29104 18222 29132 18634
rect 29196 18358 29224 18702
rect 29288 18698 29316 19246
rect 29380 19230 29500 19258
rect 29276 18692 29328 18698
rect 29276 18634 29328 18640
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29184 18352 29236 18358
rect 29184 18294 29236 18300
rect 29092 18216 29144 18222
rect 29092 18158 29144 18164
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28724 17672 28776 17678
rect 28724 17614 28776 17620
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 26884 17536 26936 17542
rect 26884 17478 26936 17484
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26896 17202 26924 17478
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 25688 16720 25740 16726
rect 25688 16662 25740 16668
rect 26056 16720 26108 16726
rect 26056 16662 26108 16668
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25148 16250 25176 16526
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25240 15638 25268 15982
rect 25228 15632 25280 15638
rect 25228 15574 25280 15580
rect 25700 15570 25728 16662
rect 26804 16658 26832 17138
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24044 14414 24072 14758
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 24136 14362 24164 14894
rect 24228 14498 24256 14962
rect 24412 14618 24440 15302
rect 24964 15162 24992 15438
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24228 14470 24348 14498
rect 24320 14414 24348 14470
rect 24216 14408 24268 14414
rect 24136 14356 24216 14362
rect 24136 14350 24268 14356
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24136 14334 24256 14350
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23940 13796 23992 13802
rect 23940 13738 23992 13744
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13326 23704 13670
rect 23952 13394 23980 13738
rect 24228 13462 24256 14334
rect 24320 14074 24348 14350
rect 24688 14346 24716 14758
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24676 14340 24728 14346
rect 24676 14282 24728 14288
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24688 14006 24716 14282
rect 24780 14074 24808 14418
rect 24964 14278 24992 15098
rect 26804 15026 26832 16594
rect 27816 15978 27844 17614
rect 28184 17338 28212 17614
rect 28356 17604 28408 17610
rect 28356 17546 28408 17552
rect 28264 17536 28316 17542
rect 28264 17478 28316 17484
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 28080 16652 28132 16658
rect 28080 16594 28132 16600
rect 27988 16516 28040 16522
rect 27988 16458 28040 16464
rect 28000 16046 28028 16458
rect 28092 16250 28120 16594
rect 28276 16250 28304 17478
rect 28368 17338 28396 17546
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 29104 17202 29132 17614
rect 29196 17610 29224 18294
rect 29380 18290 29408 18566
rect 29368 18284 29420 18290
rect 29368 18226 29420 18232
rect 29472 18170 29500 19230
rect 29564 18766 29592 19654
rect 29656 19446 29684 19790
rect 29644 19440 29696 19446
rect 29644 19382 29696 19388
rect 29840 19378 29868 19790
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 29932 19446 29960 19654
rect 30116 19446 30144 20198
rect 30208 19922 30236 20742
rect 31852 20528 31904 20534
rect 31852 20470 31904 20476
rect 31576 20256 31628 20262
rect 31576 20198 31628 20204
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 29920 19440 29972 19446
rect 29920 19382 29972 19388
rect 30104 19440 30156 19446
rect 30104 19382 30156 19388
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 30208 18766 30236 19858
rect 31588 19854 31616 20198
rect 31864 19990 31892 20470
rect 31956 20466 31984 20810
rect 32312 20800 32364 20806
rect 32312 20742 32364 20748
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 31852 19984 31904 19990
rect 31852 19926 31904 19932
rect 31576 19848 31628 19854
rect 31576 19790 31628 19796
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 29552 18760 29604 18766
rect 30196 18760 30248 18766
rect 29552 18702 29604 18708
rect 30116 18720 30196 18748
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29920 18624 29972 18630
rect 29920 18566 29972 18572
rect 29380 18142 29500 18170
rect 29184 17604 29236 17610
rect 29184 17546 29236 17552
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 28632 16720 28684 16726
rect 28632 16662 28684 16668
rect 28080 16244 28132 16250
rect 28080 16186 28132 16192
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 27804 15972 27856 15978
rect 27804 15914 27856 15920
rect 26884 15904 26936 15910
rect 26884 15846 26936 15852
rect 26896 15502 26924 15846
rect 27804 15632 27856 15638
rect 27804 15574 27856 15580
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 26804 14906 26832 14962
rect 25516 14618 25544 14894
rect 26804 14878 26924 14906
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25056 14482 25084 14554
rect 25228 14544 25280 14550
rect 25228 14486 25280 14492
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24952 14272 25004 14278
rect 25056 14260 25084 14418
rect 25056 14232 25176 14260
rect 24952 14214 25004 14220
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24676 14000 24728 14006
rect 24676 13942 24728 13948
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23768 12238 23796 13194
rect 23848 12844 23900 12850
rect 23952 12832 23980 13330
rect 24872 13326 24900 13806
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24964 13530 24992 13670
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24228 12850 24256 13262
rect 24964 12918 24992 13330
rect 25148 13326 25176 14232
rect 25240 13530 25268 14486
rect 26896 14482 26924 14878
rect 26988 14618 27016 15438
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27712 15360 27764 15366
rect 27712 15302 27764 15308
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 27632 14482 27660 15302
rect 27724 14958 27752 15302
rect 27712 14952 27764 14958
rect 27712 14894 27764 14900
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 27620 14476 27672 14482
rect 27620 14418 27672 14424
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26516 14408 26568 14414
rect 26516 14350 26568 14356
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 23900 12804 23980 12832
rect 24216 12844 24268 12850
rect 23848 12786 23900 12792
rect 24216 12786 24268 12792
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23860 12170 23888 12786
rect 24492 12368 24544 12374
rect 24492 12310 24544 12316
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 23952 11898 23980 12174
rect 24124 12164 24176 12170
rect 24124 12106 24176 12112
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 24136 11082 24164 12106
rect 24504 12102 24532 12310
rect 24688 12238 24716 12786
rect 24964 12306 24992 12854
rect 25148 12850 25176 13262
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 26252 12782 26280 14350
rect 26528 13802 26556 14350
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27080 14074 27108 14282
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27540 14074 27568 14214
rect 27068 14068 27120 14074
rect 27068 14010 27120 14016
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26516 13796 26568 13802
rect 26516 13738 26568 13744
rect 26528 13326 26556 13738
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26424 12912 26476 12918
rect 26424 12854 26476 12860
rect 26240 12776 26292 12782
rect 26240 12718 26292 12724
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 24136 10742 24164 11018
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23662 10296 23718 10305
rect 23662 10231 23664 10240
rect 23716 10231 23718 10240
rect 23664 10202 23716 10208
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23676 9722 23704 9998
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23664 9580 23716 9586
rect 23768 9568 23796 10610
rect 24032 10532 24084 10538
rect 24032 10474 24084 10480
rect 23938 10296 23994 10305
rect 24044 10266 24072 10474
rect 23938 10231 23940 10240
rect 23992 10231 23994 10240
rect 24032 10260 24084 10266
rect 23940 10202 23992 10208
rect 24032 10202 24084 10208
rect 23848 10022 23900 10028
rect 23900 9982 23980 10010
rect 23848 9964 23900 9970
rect 23846 9888 23902 9897
rect 23846 9823 23902 9832
rect 23716 9540 23796 9568
rect 23664 9522 23716 9528
rect 23676 7818 23704 9522
rect 23860 8498 23888 9823
rect 23952 9654 23980 9982
rect 23940 9648 23992 9654
rect 23940 9590 23992 9596
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23952 7868 23980 9590
rect 24044 9450 24072 10202
rect 24124 10056 24176 10062
rect 24122 10024 24124 10033
rect 24176 10024 24178 10033
rect 24122 9959 24178 9968
rect 24228 9897 24256 11086
rect 24320 10674 24348 11630
rect 24596 11558 24624 12106
rect 24688 11762 24716 12174
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11150 24624 11494
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24872 10810 24900 11086
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24214 9888 24270 9897
rect 24214 9823 24270 9832
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 24320 8480 24348 10610
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24490 10160 24546 10169
rect 24490 10095 24546 10104
rect 24504 10062 24532 10095
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24412 9722 24440 9998
rect 24400 9716 24452 9722
rect 24400 9658 24452 9664
rect 24596 9382 24624 10542
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24688 10130 24716 10406
rect 24858 10296 24914 10305
rect 24858 10231 24914 10240
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24584 8492 24636 8498
rect 24320 8452 24584 8480
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24214 7984 24270 7993
rect 24214 7919 24216 7928
rect 24268 7919 24270 7928
rect 24216 7890 24268 7896
rect 24320 7886 24348 8230
rect 24124 7880 24176 7886
rect 23952 7840 24124 7868
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 23860 5710 23888 7142
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23952 5234 23980 7840
rect 24124 7822 24176 7828
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24228 7546 24256 7754
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24412 6746 24440 8452
rect 24584 8434 24636 8440
rect 24676 8016 24728 8022
rect 24780 8004 24808 10066
rect 24872 9654 24900 10231
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24964 9586 24992 12038
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24872 8362 24900 8570
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24728 7976 24808 8004
rect 24676 7958 24728 7964
rect 24584 7744 24636 7750
rect 24584 7686 24636 7692
rect 24596 7410 24624 7686
rect 24780 7410 24808 7976
rect 24872 7886 24900 8298
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 24964 8022 24992 8230
rect 24952 8016 25004 8022
rect 24952 7958 25004 7964
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24964 7410 24992 7754
rect 25056 7546 25084 11494
rect 25148 10062 25176 12378
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25700 11762 25728 12038
rect 26436 11762 26464 12854
rect 26528 12850 26556 13262
rect 26620 12850 26648 13262
rect 26712 13258 26740 13874
rect 27816 13870 27844 15574
rect 28000 15094 28028 15982
rect 28644 15978 28672 16662
rect 29000 16516 29052 16522
rect 29000 16458 29052 16464
rect 29012 16046 29040 16458
rect 29104 16046 29132 17138
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29196 16794 29224 17070
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 29380 16522 29408 18142
rect 29656 17678 29684 18566
rect 29644 17672 29696 17678
rect 29644 17614 29696 17620
rect 29460 17536 29512 17542
rect 29460 17478 29512 17484
rect 29472 17202 29500 17478
rect 29932 17338 29960 18566
rect 30012 17672 30064 17678
rect 30012 17614 30064 17620
rect 29920 17332 29972 17338
rect 29920 17274 29972 17280
rect 29932 17202 29960 17274
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29920 17196 29972 17202
rect 29920 17138 29972 17144
rect 30024 16998 30052 17614
rect 30116 16998 30144 18720
rect 30196 18702 30248 18708
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30656 18352 30708 18358
rect 30656 18294 30708 18300
rect 30196 17876 30248 17882
rect 30196 17818 30248 17824
rect 30208 17678 30236 17818
rect 30288 17808 30340 17814
rect 30340 17756 30420 17762
rect 30288 17750 30420 17756
rect 30300 17734 30420 17750
rect 30392 17678 30420 17734
rect 30668 17678 30696 18294
rect 30852 17882 30880 18634
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 30944 17882 30972 18158
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 30932 17876 30984 17882
rect 30932 17818 30984 17824
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30656 17672 30708 17678
rect 30656 17614 30708 17620
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30208 17202 30236 17478
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30012 16992 30064 16998
rect 30012 16934 30064 16940
rect 30104 16992 30156 16998
rect 30104 16934 30156 16940
rect 30116 16658 30144 16934
rect 30300 16794 30328 17138
rect 30288 16788 30340 16794
rect 30288 16730 30340 16736
rect 30104 16652 30156 16658
rect 30104 16594 30156 16600
rect 29368 16516 29420 16522
rect 29368 16458 29420 16464
rect 30576 16454 30604 17478
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30668 17105 30696 17138
rect 30654 17096 30710 17105
rect 30654 17031 30710 17040
rect 30668 16454 30696 17031
rect 30944 16726 30972 17614
rect 31036 17610 31064 18770
rect 31024 17604 31076 17610
rect 31024 17546 31076 17552
rect 31036 17270 31064 17546
rect 31024 17264 31076 17270
rect 31024 17206 31076 17212
rect 30932 16720 30984 16726
rect 30932 16662 30984 16668
rect 29460 16448 29512 16454
rect 29460 16390 29512 16396
rect 30472 16448 30524 16454
rect 30472 16390 30524 16396
rect 30564 16448 30616 16454
rect 30564 16390 30616 16396
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 29472 16114 29500 16390
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 29092 16040 29144 16046
rect 29092 15982 29144 15988
rect 28632 15972 28684 15978
rect 28632 15914 28684 15920
rect 28172 15428 28224 15434
rect 28172 15370 28224 15376
rect 28184 15162 28212 15370
rect 29472 15162 29500 16050
rect 30484 16046 30512 16390
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 30472 16040 30524 16046
rect 30472 15982 30524 15988
rect 28172 15156 28224 15162
rect 28172 15098 28224 15104
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 27988 15088 28040 15094
rect 27988 15030 28040 15036
rect 28000 14362 28028 15030
rect 27908 14346 28028 14362
rect 27896 14340 28028 14346
rect 27948 14334 28028 14340
rect 27896 14282 27948 14288
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27908 13462 27936 14282
rect 28184 13802 28212 15098
rect 29564 14482 29592 15982
rect 30668 15910 30696 16390
rect 31220 16182 31248 19722
rect 31588 19446 31616 19790
rect 32324 19786 32352 20742
rect 32600 19854 32628 20810
rect 33048 20528 33100 20534
rect 33046 20496 33048 20505
rect 33100 20496 33102 20505
rect 33046 20431 33102 20440
rect 33888 20398 33916 20878
rect 34440 20602 34468 21966
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34428 20596 34480 20602
rect 34428 20538 34480 20544
rect 33968 20460 34020 20466
rect 33968 20402 34020 20408
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 33600 20392 33652 20398
rect 33600 20334 33652 20340
rect 33876 20392 33928 20398
rect 33876 20334 33928 20340
rect 33612 19990 33640 20334
rect 33692 20324 33744 20330
rect 33692 20266 33744 20272
rect 33600 19984 33652 19990
rect 33600 19926 33652 19932
rect 32588 19848 32640 19854
rect 32588 19790 32640 19796
rect 32680 19848 32732 19854
rect 32680 19790 32732 19796
rect 32128 19780 32180 19786
rect 32128 19722 32180 19728
rect 32312 19780 32364 19786
rect 32312 19722 32364 19728
rect 32140 19514 32168 19722
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 32128 19508 32180 19514
rect 32128 19450 32180 19456
rect 31576 19440 31628 19446
rect 31576 19382 31628 19388
rect 31392 19168 31444 19174
rect 31392 19110 31444 19116
rect 31404 18358 31432 19110
rect 31772 18902 31800 19450
rect 32324 19378 32352 19722
rect 32600 19514 32628 19790
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 32692 19446 32720 19790
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 32680 19440 32732 19446
rect 32680 19382 32732 19388
rect 33244 19378 33272 19654
rect 33324 19508 33376 19514
rect 33324 19450 33376 19456
rect 33600 19508 33652 19514
rect 33600 19450 33652 19456
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 33232 19372 33284 19378
rect 33232 19314 33284 19320
rect 31760 18896 31812 18902
rect 32324 18850 32352 19314
rect 33140 19236 33192 19242
rect 33140 19178 33192 19184
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 33048 19168 33100 19174
rect 33048 19110 33100 19116
rect 31760 18838 31812 18844
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31956 18822 32352 18850
rect 32496 18896 32548 18902
rect 32496 18838 32548 18844
rect 31496 18698 31524 18770
rect 31484 18692 31536 18698
rect 31484 18634 31536 18640
rect 31392 18352 31444 18358
rect 31392 18294 31444 18300
rect 31668 18148 31720 18154
rect 31668 18090 31720 18096
rect 31680 17678 31708 18090
rect 31668 17672 31720 17678
rect 31668 17614 31720 17620
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 31392 16992 31444 16998
rect 31392 16934 31444 16940
rect 31760 16992 31812 16998
rect 31956 16980 31984 18822
rect 32128 18760 32180 18766
rect 32128 18702 32180 18708
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32140 18358 32168 18702
rect 32128 18352 32180 18358
rect 32128 18294 32180 18300
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 32048 17678 32076 18226
rect 32140 17746 32168 18294
rect 32232 17746 32260 18702
rect 32128 17740 32180 17746
rect 32128 17682 32180 17688
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 32036 17672 32088 17678
rect 32036 17614 32088 17620
rect 32324 17218 32352 17682
rect 32508 17678 32536 18838
rect 32784 18766 32812 19110
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32588 18692 32640 18698
rect 32588 18634 32640 18640
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 32496 17672 32548 17678
rect 32496 17614 32548 17620
rect 32416 17338 32444 17614
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32232 17202 32352 17218
rect 32220 17196 32352 17202
rect 32272 17190 32352 17196
rect 32220 17138 32272 17144
rect 31812 16952 31984 16980
rect 31760 16934 31812 16940
rect 31312 16726 31340 16934
rect 31300 16720 31352 16726
rect 31300 16662 31352 16668
rect 31404 16590 31432 16934
rect 31772 16658 31800 16934
rect 31760 16652 31812 16658
rect 31760 16594 31812 16600
rect 31392 16584 31444 16590
rect 31392 16526 31444 16532
rect 31404 16250 31432 16526
rect 31668 16448 31720 16454
rect 31668 16390 31720 16396
rect 31392 16244 31444 16250
rect 31392 16186 31444 16192
rect 31680 16182 31708 16390
rect 32232 16250 32260 17138
rect 32416 16658 32444 17274
rect 32496 17264 32548 17270
rect 32496 17206 32548 17212
rect 32508 16726 32536 17206
rect 32600 17202 32628 18634
rect 32680 17536 32732 17542
rect 32680 17478 32732 17484
rect 32588 17196 32640 17202
rect 32588 17138 32640 17144
rect 32496 16720 32548 16726
rect 32496 16662 32548 16668
rect 32692 16658 32720 17478
rect 32784 17116 32812 18702
rect 33060 18290 33088 19110
rect 33152 18834 33180 19178
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33048 18284 33100 18290
rect 33048 18226 33100 18232
rect 33232 18216 33284 18222
rect 33232 18158 33284 18164
rect 33244 17882 33272 18158
rect 33336 17882 33364 19450
rect 33508 19372 33560 19378
rect 33508 19314 33560 19320
rect 33520 18970 33548 19314
rect 33508 18964 33560 18970
rect 33508 18906 33560 18912
rect 33416 18896 33468 18902
rect 33416 18838 33468 18844
rect 33428 18290 33456 18838
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 33416 18284 33468 18290
rect 33416 18226 33468 18232
rect 33520 18086 33548 18702
rect 33612 18630 33640 19450
rect 33704 18698 33732 20266
rect 33980 19990 34008 20402
rect 33968 19984 34020 19990
rect 33968 19926 34020 19932
rect 34164 19854 34192 20402
rect 34152 19848 34204 19854
rect 34152 19790 34204 19796
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33796 19378 33824 19654
rect 34164 19514 34192 19790
rect 34336 19780 34388 19786
rect 34336 19722 34388 19728
rect 34152 19508 34204 19514
rect 34152 19450 34204 19456
rect 33784 19372 33836 19378
rect 33784 19314 33836 19320
rect 34348 19310 34376 19722
rect 34336 19304 34388 19310
rect 34336 19246 34388 19252
rect 34152 19168 34204 19174
rect 34152 19110 34204 19116
rect 34164 18834 34192 19110
rect 34152 18828 34204 18834
rect 34152 18770 34204 18776
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33600 18624 33652 18630
rect 33600 18566 33652 18572
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33508 18080 33560 18086
rect 33508 18022 33560 18028
rect 33612 17882 33640 18158
rect 33232 17876 33284 17882
rect 33232 17818 33284 17824
rect 33324 17876 33376 17882
rect 33324 17818 33376 17824
rect 33600 17876 33652 17882
rect 33600 17818 33652 17824
rect 33336 17678 33364 17818
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 33140 17196 33192 17202
rect 33140 17138 33192 17144
rect 32956 17128 33008 17134
rect 32784 17088 32956 17116
rect 32956 17070 33008 17076
rect 33152 16794 33180 17138
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 32404 16652 32456 16658
rect 32404 16594 32456 16600
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 32772 16584 32824 16590
rect 32824 16544 32904 16572
rect 32772 16526 32824 16532
rect 32220 16244 32272 16250
rect 32220 16186 32272 16192
rect 31208 16176 31260 16182
rect 31208 16118 31260 16124
rect 31668 16176 31720 16182
rect 31668 16118 31720 16124
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30104 15360 30156 15366
rect 30104 15302 30156 15308
rect 30116 15162 30144 15302
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 29828 15020 29880 15026
rect 29828 14962 29880 14968
rect 30748 15020 30800 15026
rect 30748 14962 30800 14968
rect 29840 14618 29868 14962
rect 29828 14612 29880 14618
rect 29828 14554 29880 14560
rect 30760 14600 30788 14962
rect 31024 14816 31076 14822
rect 31024 14758 31076 14764
rect 30840 14612 30892 14618
rect 30760 14572 30840 14600
rect 29552 14476 29604 14482
rect 29552 14418 29604 14424
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28644 13938 28672 14214
rect 29380 14074 29408 14350
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29840 14006 29868 14554
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 29828 14000 29880 14006
rect 29828 13942 29880 13948
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28540 13864 28592 13870
rect 28540 13806 28592 13812
rect 28172 13796 28224 13802
rect 28172 13738 28224 13744
rect 27896 13456 27948 13462
rect 27896 13398 27948 13404
rect 26700 13252 26752 13258
rect 26700 13194 26752 13200
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 26712 12918 26740 13194
rect 26884 13184 26936 13190
rect 26884 13126 26936 13132
rect 26700 12912 26752 12918
rect 26700 12854 26752 12860
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26528 12238 26556 12786
rect 26516 12232 26568 12238
rect 26516 12174 26568 12180
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 25976 11354 26004 11698
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25688 10736 25740 10742
rect 25688 10678 25740 10684
rect 25700 10130 25728 10678
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25688 10124 25740 10130
rect 25688 10066 25740 10072
rect 25136 10056 25188 10062
rect 25188 10004 25360 10010
rect 25136 9998 25360 10004
rect 25148 9982 25360 9998
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 7546 25176 9862
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25240 8634 25268 8910
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25226 8528 25282 8537
rect 25226 8463 25228 8472
rect 25280 8463 25282 8472
rect 25228 8434 25280 8440
rect 25228 8016 25280 8022
rect 25226 7984 25228 7993
rect 25280 7984 25282 7993
rect 25226 7919 25282 7928
rect 25332 7886 25360 9982
rect 25700 9654 25728 10066
rect 25792 9994 25820 10610
rect 25976 10062 26004 11086
rect 26056 10600 26108 10606
rect 26056 10542 26108 10548
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 25780 9988 25832 9994
rect 25780 9930 25832 9936
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25792 9586 25820 9930
rect 25976 9722 26004 9998
rect 25964 9716 26016 9722
rect 25964 9658 26016 9664
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25792 9110 25820 9522
rect 25780 9104 25832 9110
rect 25780 9046 25832 9052
rect 25976 8906 26004 9658
rect 26068 9518 26096 10542
rect 26160 10538 26188 11698
rect 26252 11150 26280 11698
rect 26528 11150 26556 12174
rect 26620 11762 26648 12786
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26804 12170 26832 12582
rect 26896 12442 26924 13126
rect 27632 12986 27660 13194
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27908 12918 27936 13398
rect 28184 13394 28212 13738
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27896 12912 27948 12918
rect 27896 12854 27948 12860
rect 27252 12776 27304 12782
rect 27252 12718 27304 12724
rect 27264 12442 27292 12718
rect 26884 12436 26936 12442
rect 26884 12378 26936 12384
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 27540 12170 27568 12854
rect 28276 12442 28304 13126
rect 28552 12866 28580 13806
rect 28644 13462 28672 13874
rect 30208 13818 30236 14418
rect 30208 13790 30420 13818
rect 30196 13728 30248 13734
rect 30196 13670 30248 13676
rect 29828 13524 29880 13530
rect 29828 13466 29880 13472
rect 28632 13456 28684 13462
rect 28632 13398 28684 13404
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28644 12986 28672 13262
rect 28724 13252 28776 13258
rect 28724 13194 28776 13200
rect 29092 13252 29144 13258
rect 29092 13194 29144 13200
rect 28632 12980 28684 12986
rect 28632 12922 28684 12928
rect 28552 12838 28672 12866
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 28264 12436 28316 12442
rect 28264 12378 28316 12384
rect 28552 12374 28580 12718
rect 28540 12368 28592 12374
rect 28540 12310 28592 12316
rect 26792 12164 26844 12170
rect 26792 12106 26844 12112
rect 27528 12164 27580 12170
rect 27528 12106 27580 12112
rect 28356 12096 28408 12102
rect 28644 12084 28672 12838
rect 28736 12646 28764 13194
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 28736 12374 28764 12582
rect 28828 12374 28856 12922
rect 28724 12368 28776 12374
rect 28724 12310 28776 12316
rect 28816 12368 28868 12374
rect 28816 12310 28868 12316
rect 28408 12056 28672 12084
rect 28356 12038 28408 12044
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 26988 11626 27016 11698
rect 26608 11620 26660 11626
rect 26608 11562 26660 11568
rect 26976 11620 27028 11626
rect 26976 11562 27028 11568
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26332 11144 26384 11150
rect 26332 11086 26384 11092
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26344 11014 26372 11086
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26344 10674 26372 10950
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26148 10532 26200 10538
rect 26148 10474 26200 10480
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 26160 9178 26188 10066
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26148 9172 26200 9178
rect 26068 9132 26148 9160
rect 26068 9042 26096 9132
rect 26148 9114 26200 9120
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 25596 8900 25648 8906
rect 25596 8842 25648 8848
rect 25964 8900 26016 8906
rect 25964 8842 26016 8848
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25056 7410 25084 7482
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 24676 7268 24728 7274
rect 24676 7210 24728 7216
rect 24412 6718 24532 6746
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24412 6458 24440 6598
rect 24504 6458 24532 6718
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24504 6338 24532 6394
rect 24688 6390 24716 7210
rect 24964 7206 24992 7346
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 24228 6322 24532 6338
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 24216 6316 24532 6322
rect 24268 6310 24532 6316
rect 24216 6258 24268 6264
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 24320 5370 24348 5714
rect 24688 5642 24716 6326
rect 25056 6322 25084 7346
rect 25148 6798 25176 7346
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25148 6322 25176 6734
rect 25424 6730 25452 8774
rect 25516 8498 25544 8774
rect 25608 8566 25636 8842
rect 25596 8560 25648 8566
rect 25596 8502 25648 8508
rect 26252 8498 26280 9522
rect 26436 9382 26464 10610
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 26344 8634 26372 8910
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 25504 8492 25556 8498
rect 25504 8434 25556 8440
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 26620 8294 26648 11562
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28276 11218 28304 11494
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28540 11212 28592 11218
rect 28540 11154 28592 11160
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27896 11144 27948 11150
rect 27896 11086 27948 11092
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27172 10266 27200 10610
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 27816 10198 27844 11086
rect 27908 10538 27936 11086
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 27896 10532 27948 10538
rect 27896 10474 27948 10480
rect 27804 10192 27856 10198
rect 27804 10134 27856 10140
rect 27436 9988 27488 9994
rect 27436 9930 27488 9936
rect 27448 8566 27476 9930
rect 27816 9654 27844 10134
rect 27804 9648 27856 9654
rect 27804 9590 27856 9596
rect 27988 8900 28040 8906
rect 27988 8842 28040 8848
rect 28000 8634 28028 8842
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 27436 8560 27488 8566
rect 27436 8502 27488 8508
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 27080 8090 27108 8366
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26804 7546 26832 7822
rect 27172 7818 27200 8434
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 27160 7812 27212 7818
rect 27160 7754 27212 7760
rect 27356 7546 27384 7822
rect 26792 7540 26844 7546
rect 26792 7482 26844 7488
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27448 7274 27476 8502
rect 28092 8498 28120 10950
rect 28552 10742 28580 11154
rect 28828 11150 28856 12310
rect 28816 11144 28868 11150
rect 28816 11086 28868 11092
rect 29104 11082 29132 13194
rect 29736 13184 29788 13190
rect 29736 13126 29788 13132
rect 29748 12238 29776 13126
rect 29840 12918 29868 13466
rect 29828 12912 29880 12918
rect 29828 12854 29880 12860
rect 29840 12374 29868 12854
rect 30208 12646 30236 13670
rect 30392 13394 30420 13790
rect 30656 13796 30708 13802
rect 30656 13738 30708 13744
rect 30380 13388 30432 13394
rect 30380 13330 30432 13336
rect 30392 12918 30420 13330
rect 30668 12986 30696 13738
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30196 12640 30248 12646
rect 30196 12582 30248 12588
rect 30208 12442 30236 12582
rect 30196 12436 30248 12442
rect 30196 12378 30248 12384
rect 29828 12368 29880 12374
rect 29828 12310 29880 12316
rect 30760 12238 30788 14572
rect 30840 14554 30892 14560
rect 30932 14544 30984 14550
rect 30932 14486 30984 14492
rect 30944 13938 30972 14486
rect 31036 14074 31064 14758
rect 31220 14498 31248 16118
rect 32876 16046 32904 16544
rect 33336 16522 33364 17614
rect 33704 17202 33732 18634
rect 34348 18578 34376 19246
rect 34716 19174 34744 21830
rect 35268 21690 35296 22034
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 35360 21690 35388 21966
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 36004 21146 36032 22066
rect 35992 21140 36044 21146
rect 35992 21082 36044 21088
rect 35440 20936 35492 20942
rect 35440 20878 35492 20884
rect 35992 20936 36044 20942
rect 36044 20896 36124 20924
rect 35992 20878 36044 20884
rect 35452 20602 35480 20878
rect 35992 20800 36044 20806
rect 35992 20742 36044 20748
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35440 20596 35492 20602
rect 35440 20538 35492 20544
rect 36004 20505 36032 20742
rect 36096 20534 36124 20896
rect 36188 20602 36216 24278
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36372 23866 36400 24142
rect 36636 24132 36688 24138
rect 36636 24074 36688 24080
rect 36360 23860 36412 23866
rect 36360 23802 36412 23808
rect 36648 23798 36676 24074
rect 36636 23792 36688 23798
rect 36636 23734 36688 23740
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 36280 23322 36308 23666
rect 36636 23656 36688 23662
rect 36636 23598 36688 23604
rect 36268 23316 36320 23322
rect 36268 23258 36320 23264
rect 36648 23186 36676 23598
rect 36912 23520 36964 23526
rect 36912 23462 36964 23468
rect 36924 23322 36952 23462
rect 37292 23322 37320 23666
rect 36912 23316 36964 23322
rect 36912 23258 36964 23264
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 36636 23180 36688 23186
rect 36636 23122 36688 23128
rect 36648 22778 36676 23122
rect 37384 23118 37412 26318
rect 37476 25974 37504 26386
rect 37464 25968 37516 25974
rect 37464 25910 37516 25916
rect 37476 25498 37504 25910
rect 37568 25838 37596 26794
rect 37752 26586 37780 27610
rect 38028 27470 38056 27882
rect 38200 27872 38252 27878
rect 38200 27814 38252 27820
rect 37924 27464 37976 27470
rect 37924 27406 37976 27412
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 37936 27130 37964 27406
rect 37924 27124 37976 27130
rect 37924 27066 37976 27072
rect 38028 26926 38056 27406
rect 38212 26994 38240 27814
rect 38382 27296 38438 27305
rect 38382 27231 38438 27240
rect 38396 27130 38424 27231
rect 38384 27124 38436 27130
rect 38384 27066 38436 27072
rect 38200 26988 38252 26994
rect 38200 26930 38252 26936
rect 38016 26920 38068 26926
rect 38016 26862 38068 26868
rect 37740 26580 37792 26586
rect 37740 26522 37792 26528
rect 38016 26512 38068 26518
rect 38016 26454 38068 26460
rect 37648 26308 37700 26314
rect 37648 26250 37700 26256
rect 37556 25832 37608 25838
rect 37556 25774 37608 25780
rect 37464 25492 37516 25498
rect 37464 25434 37516 25440
rect 37464 23724 37516 23730
rect 37464 23666 37516 23672
rect 37476 23254 37504 23666
rect 37464 23248 37516 23254
rect 37660 23202 37688 26250
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 37844 25498 37872 25842
rect 37832 25492 37884 25498
rect 37832 25434 37884 25440
rect 37740 25288 37792 25294
rect 37924 25288 37976 25294
rect 37792 25236 37872 25242
rect 37740 25230 37872 25236
rect 37924 25230 37976 25236
rect 37752 25214 37872 25230
rect 37844 25158 37872 25214
rect 37832 25152 37884 25158
rect 37832 25094 37884 25100
rect 37464 23190 37516 23196
rect 37568 23174 37688 23202
rect 36728 23112 36780 23118
rect 36728 23054 36780 23060
rect 36912 23112 36964 23118
rect 36912 23054 36964 23060
rect 37188 23112 37240 23118
rect 37188 23054 37240 23060
rect 37372 23112 37424 23118
rect 37372 23054 37424 23060
rect 36740 22778 36768 23054
rect 36636 22772 36688 22778
rect 36636 22714 36688 22720
rect 36728 22772 36780 22778
rect 36728 22714 36780 22720
rect 36452 22636 36504 22642
rect 36452 22578 36504 22584
rect 36636 22636 36688 22642
rect 36636 22578 36688 22584
rect 36464 22234 36492 22578
rect 36648 22506 36676 22578
rect 36636 22500 36688 22506
rect 36636 22442 36688 22448
rect 36452 22228 36504 22234
rect 36452 22170 36504 22176
rect 36360 21344 36412 21350
rect 36360 21286 36412 21292
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36084 20528 36136 20534
rect 35990 20496 36046 20505
rect 36084 20470 36136 20476
rect 35990 20431 36046 20440
rect 35808 20392 35860 20398
rect 35808 20334 35860 20340
rect 35992 20392 36044 20398
rect 35992 20334 36044 20340
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35820 19990 35848 20334
rect 36004 20262 36032 20334
rect 35900 20256 35952 20262
rect 35900 20198 35952 20204
rect 35992 20256 36044 20262
rect 35992 20198 36044 20204
rect 35808 19984 35860 19990
rect 35808 19926 35860 19932
rect 35912 19854 35940 20198
rect 36004 19922 36032 20198
rect 35992 19916 36044 19922
rect 35992 19858 36044 19864
rect 35900 19848 35952 19854
rect 35900 19790 35952 19796
rect 36096 19786 36124 20470
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 36084 19780 36136 19786
rect 36084 19722 36136 19728
rect 36188 19718 36216 20402
rect 36372 20330 36400 21286
rect 36544 20936 36596 20942
rect 36544 20878 36596 20884
rect 36452 20800 36504 20806
rect 36452 20742 36504 20748
rect 36360 20324 36412 20330
rect 36360 20266 36412 20272
rect 36268 19848 36320 19854
rect 36268 19790 36320 19796
rect 35440 19712 35492 19718
rect 35440 19654 35492 19660
rect 36176 19712 36228 19718
rect 36176 19654 36228 19660
rect 35452 19514 35480 19654
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 36280 19514 36308 19790
rect 35440 19508 35492 19514
rect 35440 19450 35492 19456
rect 35716 19508 35768 19514
rect 35716 19450 35768 19456
rect 36268 19508 36320 19514
rect 36268 19450 36320 19456
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 34704 19168 34756 19174
rect 34704 19110 34756 19116
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34440 18698 34468 18906
rect 34428 18692 34480 18698
rect 34428 18634 34480 18640
rect 34716 18630 34744 19110
rect 34612 18624 34664 18630
rect 34348 18550 34468 18578
rect 34612 18566 34664 18572
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34440 18426 34468 18550
rect 34428 18420 34480 18426
rect 34428 18362 34480 18368
rect 34520 18352 34572 18358
rect 34520 18294 34572 18300
rect 34428 18216 34480 18222
rect 34428 18158 34480 18164
rect 34244 18080 34296 18086
rect 34244 18022 34296 18028
rect 34256 17202 34284 18022
rect 34440 17678 34468 18158
rect 34532 17814 34560 18294
rect 34624 18290 34652 18566
rect 34612 18284 34664 18290
rect 34612 18226 34664 18232
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 34520 17808 34572 17814
rect 34520 17750 34572 17756
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 34440 17270 34468 17614
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 33692 17196 33744 17202
rect 33692 17138 33744 17144
rect 34244 17196 34296 17202
rect 34244 17138 34296 17144
rect 33414 17096 33470 17105
rect 33414 17031 33416 17040
rect 33468 17031 33470 17040
rect 33416 17002 33468 17008
rect 33704 16998 33732 17138
rect 34532 17066 34560 17750
rect 34612 17672 34664 17678
rect 34612 17614 34664 17620
rect 34624 17134 34652 17614
rect 34716 17610 34744 18226
rect 34808 17746 34836 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35728 18970 35756 19450
rect 36084 19440 36136 19446
rect 35990 19408 36046 19417
rect 36084 19382 36136 19388
rect 35990 19343 35992 19352
rect 36044 19343 36046 19352
rect 35992 19314 36044 19320
rect 36096 18970 36124 19382
rect 36372 19378 36400 20266
rect 36464 20058 36492 20742
rect 36452 20052 36504 20058
rect 36452 19994 36504 20000
rect 36464 19786 36492 19994
rect 36556 19922 36584 20878
rect 36544 19916 36596 19922
rect 36544 19858 36596 19864
rect 36452 19780 36504 19786
rect 36452 19722 36504 19728
rect 36648 19514 36676 22442
rect 36728 21548 36780 21554
rect 36728 21490 36780 21496
rect 36740 21146 36768 21490
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36728 20936 36780 20942
rect 36728 20878 36780 20884
rect 36740 20262 36768 20878
rect 36728 20256 36780 20262
rect 36728 20198 36780 20204
rect 36740 20058 36768 20198
rect 36728 20052 36780 20058
rect 36728 19994 36780 20000
rect 36636 19508 36688 19514
rect 36636 19450 36688 19456
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 36360 19372 36412 19378
rect 36360 19314 36412 19320
rect 36176 19168 36228 19174
rect 36280 19156 36308 19314
rect 36228 19128 36308 19156
rect 36176 19110 36228 19116
rect 35716 18964 35768 18970
rect 35716 18906 35768 18912
rect 36084 18964 36136 18970
rect 36084 18906 36136 18912
rect 36188 18902 36216 19110
rect 36176 18896 36228 18902
rect 36176 18838 36228 18844
rect 36372 18834 36400 19314
rect 36648 19242 36676 19450
rect 36924 19446 36952 23054
rect 37200 22094 37228 23054
rect 37372 22976 37424 22982
rect 37372 22918 37424 22924
rect 37280 22704 37332 22710
rect 37280 22646 37332 22652
rect 37292 22098 37320 22646
rect 37108 22066 37228 22094
rect 37280 22092 37332 22098
rect 37108 22030 37136 22066
rect 37280 22034 37332 22040
rect 37384 22030 37412 22918
rect 37568 22642 37596 23174
rect 37648 23112 37700 23118
rect 37648 23054 37700 23060
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37464 22568 37516 22574
rect 37464 22510 37516 22516
rect 37096 22024 37148 22030
rect 37096 21966 37148 21972
rect 37372 22024 37424 22030
rect 37372 21966 37424 21972
rect 36912 19440 36964 19446
rect 36818 19408 36874 19417
rect 36912 19382 36964 19388
rect 36818 19343 36820 19352
rect 36872 19343 36874 19352
rect 37004 19372 37056 19378
rect 36820 19314 36872 19320
rect 37004 19314 37056 19320
rect 36636 19236 36688 19242
rect 36636 19178 36688 19184
rect 37016 19174 37044 19314
rect 37004 19168 37056 19174
rect 37004 19110 37056 19116
rect 34980 18828 35032 18834
rect 34980 18770 35032 18776
rect 36360 18828 36412 18834
rect 36360 18770 36412 18776
rect 34992 18290 35020 18770
rect 36636 18760 36688 18766
rect 36636 18702 36688 18708
rect 35256 18624 35308 18630
rect 35256 18566 35308 18572
rect 35268 18290 35296 18566
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 34980 18284 35032 18290
rect 34980 18226 35032 18232
rect 35256 18284 35308 18290
rect 35256 18226 35308 18232
rect 35808 18080 35860 18086
rect 35808 18022 35860 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35820 17746 35848 18022
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 35808 17740 35860 17746
rect 35808 17682 35860 17688
rect 34704 17604 34756 17610
rect 34704 17546 34756 17552
rect 36176 17604 36228 17610
rect 36176 17546 36228 17552
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 34612 17128 34664 17134
rect 34612 17070 34664 17076
rect 34520 17060 34572 17066
rect 34520 17002 34572 17008
rect 33692 16992 33744 16998
rect 33692 16934 33744 16940
rect 33324 16516 33376 16522
rect 33324 16458 33376 16464
rect 34624 16046 34652 17070
rect 34808 16794 34836 17478
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35992 17196 36044 17202
rect 35992 17138 36044 17144
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35348 16108 35400 16114
rect 35348 16050 35400 16056
rect 32864 16040 32916 16046
rect 32864 15982 32916 15988
rect 34612 16040 34664 16046
rect 34612 15982 34664 15988
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 32876 15570 32904 15982
rect 33140 15972 33192 15978
rect 33140 15914 33192 15920
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 32864 15564 32916 15570
rect 32864 15506 32916 15512
rect 32876 15026 32904 15506
rect 32968 15434 32996 15846
rect 32956 15428 33008 15434
rect 32956 15370 33008 15376
rect 33152 15094 33180 15914
rect 34428 15428 34480 15434
rect 34428 15370 34480 15376
rect 34520 15428 34572 15434
rect 34520 15370 34572 15376
rect 34440 15094 34468 15370
rect 33140 15088 33192 15094
rect 33140 15030 33192 15036
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 32864 15020 32916 15026
rect 32864 14962 32916 14968
rect 32876 14550 32904 14962
rect 34532 14618 34560 15370
rect 34704 15360 34756 15366
rect 34704 15302 34756 15308
rect 34612 14816 34664 14822
rect 34612 14758 34664 14764
rect 34520 14612 34572 14618
rect 34520 14554 34572 14560
rect 34624 14550 34652 14758
rect 31128 14470 31248 14498
rect 32864 14544 32916 14550
rect 32864 14486 32916 14492
rect 34612 14544 34664 14550
rect 34612 14486 34664 14492
rect 34716 14482 34744 15302
rect 34808 14958 34836 15982
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 14952 34848 14958
rect 34796 14894 34848 14900
rect 34808 14482 34836 14894
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34704 14476 34756 14482
rect 31128 14346 31156 14470
rect 34704 14418 34756 14424
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 35072 14408 35124 14414
rect 35072 14350 35124 14356
rect 31116 14340 31168 14346
rect 31116 14282 31168 14288
rect 31208 14340 31260 14346
rect 31208 14282 31260 14288
rect 34796 14340 34848 14346
rect 34796 14282 34848 14288
rect 31220 14074 31248 14282
rect 31300 14272 31352 14278
rect 31300 14214 31352 14220
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 31208 14068 31260 14074
rect 31208 14010 31260 14016
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30944 12238 30972 13874
rect 31312 13530 31340 14214
rect 34612 14000 34664 14006
rect 34612 13942 34664 13948
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 33508 13932 33560 13938
rect 33508 13874 33560 13880
rect 31576 13728 31628 13734
rect 31576 13670 31628 13676
rect 31300 13524 31352 13530
rect 31300 13466 31352 13472
rect 31312 13258 31340 13466
rect 31116 13252 31168 13258
rect 31116 13194 31168 13200
rect 31300 13252 31352 13258
rect 31300 13194 31352 13200
rect 31128 12986 31156 13194
rect 31208 13184 31260 13190
rect 31208 13126 31260 13132
rect 31116 12980 31168 12986
rect 31116 12922 31168 12928
rect 31220 12866 31248 13126
rect 31312 12986 31340 13194
rect 31300 12980 31352 12986
rect 31300 12922 31352 12928
rect 31128 12850 31248 12866
rect 31588 12850 31616 13670
rect 31116 12844 31248 12850
rect 31168 12838 31248 12844
rect 31484 12844 31536 12850
rect 31116 12786 31168 12792
rect 31484 12786 31536 12792
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 31128 12434 31156 12786
rect 31208 12776 31260 12782
rect 31208 12718 31260 12724
rect 31220 12442 31248 12718
rect 31300 12640 31352 12646
rect 31300 12582 31352 12588
rect 31036 12406 31156 12434
rect 31208 12436 31260 12442
rect 29736 12232 29788 12238
rect 29736 12174 29788 12180
rect 30748 12232 30800 12238
rect 30748 12174 30800 12180
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 29748 11830 29776 12174
rect 30840 12096 30892 12102
rect 30840 12038 30892 12044
rect 29736 11824 29788 11830
rect 29736 11766 29788 11772
rect 30196 11348 30248 11354
rect 30196 11290 30248 11296
rect 30208 11150 30236 11290
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 30104 11144 30156 11150
rect 30104 11086 30156 11092
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 29092 11076 29144 11082
rect 29092 11018 29144 11024
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 29196 10810 29224 11018
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 28540 10736 28592 10742
rect 28540 10678 28592 10684
rect 28264 10464 28316 10470
rect 28264 10406 28316 10412
rect 28276 10062 28304 10406
rect 28552 10266 28580 10678
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 29012 10266 29040 10610
rect 30024 10606 30052 11086
rect 30116 11014 30144 11086
rect 30104 11008 30156 11014
rect 30104 10950 30156 10956
rect 30208 10810 30236 11086
rect 30472 11008 30524 11014
rect 30472 10950 30524 10956
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30484 10674 30512 10950
rect 30668 10674 30696 10950
rect 30852 10674 30880 12038
rect 30944 11286 30972 12174
rect 31036 12170 31064 12406
rect 31208 12378 31260 12384
rect 31312 12170 31340 12582
rect 31392 12368 31444 12374
rect 31392 12310 31444 12316
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 31300 12164 31352 12170
rect 31300 12106 31352 12112
rect 31036 11762 31064 12106
rect 31208 12096 31260 12102
rect 31404 12050 31432 12310
rect 31260 12044 31432 12050
rect 31208 12038 31432 12044
rect 31220 12022 31432 12038
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 30932 11280 30984 11286
rect 30932 11222 30984 11228
rect 30944 11082 30972 11222
rect 31036 11150 31064 11698
rect 31404 11694 31432 12022
rect 31496 11762 31524 12786
rect 31680 12102 31708 13874
rect 31760 13796 31812 13802
rect 31760 13738 31812 13744
rect 31772 12850 31800 13738
rect 32864 13728 32916 13734
rect 32864 13670 32916 13676
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 32680 12708 32732 12714
rect 32680 12650 32732 12656
rect 32692 12374 32720 12650
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31668 12096 31720 12102
rect 31668 12038 31720 12044
rect 31484 11756 31536 11762
rect 31484 11698 31536 11704
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31576 11620 31628 11626
rect 31576 11562 31628 11568
rect 31024 11144 31076 11150
rect 31024 11086 31076 11092
rect 30932 11076 30984 11082
rect 30932 11018 30984 11024
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 30472 10668 30524 10674
rect 30472 10610 30524 10616
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 31024 10668 31076 10674
rect 31024 10610 31076 10616
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 28540 10260 28592 10266
rect 28540 10202 28592 10208
rect 29000 10260 29052 10266
rect 29000 10202 29052 10208
rect 29104 10198 29132 10542
rect 30116 10266 30144 10610
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 30300 10198 30328 10542
rect 30748 10464 30800 10470
rect 30748 10406 30800 10412
rect 29092 10192 29144 10198
rect 29092 10134 29144 10140
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 28448 9988 28500 9994
rect 28448 9930 28500 9936
rect 28460 9722 28488 9930
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 29104 9586 29132 10134
rect 29644 10124 29696 10130
rect 29644 10066 29696 10072
rect 29656 9722 29684 10066
rect 30760 10062 30788 10406
rect 31036 10266 31064 10610
rect 31116 10600 31168 10606
rect 31116 10542 31168 10548
rect 31024 10260 31076 10266
rect 31024 10202 31076 10208
rect 31128 10130 31156 10542
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 31588 10062 31616 11562
rect 31772 11354 31800 12174
rect 32692 11558 32720 12310
rect 32784 12306 32812 13330
rect 32876 13258 32904 13670
rect 32864 13252 32916 13258
rect 32864 13194 32916 13200
rect 33520 13190 33548 13874
rect 34336 13320 34388 13326
rect 34336 13262 34388 13268
rect 33508 13184 33560 13190
rect 33508 13126 33560 13132
rect 33416 12980 33468 12986
rect 33416 12922 33468 12928
rect 33232 12912 33284 12918
rect 33232 12854 33284 12860
rect 33140 12640 33192 12646
rect 33140 12582 33192 12588
rect 33152 12306 33180 12582
rect 32772 12300 32824 12306
rect 32772 12242 32824 12248
rect 33140 12300 33192 12306
rect 33140 12242 33192 12248
rect 32772 12164 32824 12170
rect 32772 12106 32824 12112
rect 32784 11694 32812 12106
rect 33244 11898 33272 12854
rect 33428 12306 33456 12922
rect 33520 12442 33548 13126
rect 33508 12436 33560 12442
rect 33508 12378 33560 12384
rect 33416 12300 33468 12306
rect 33520 12288 33548 12378
rect 33520 12260 33640 12288
rect 33416 12242 33468 12248
rect 33232 11892 33284 11898
rect 33232 11834 33284 11840
rect 32772 11688 32824 11694
rect 32772 11630 32824 11636
rect 33232 11688 33284 11694
rect 33232 11630 33284 11636
rect 32680 11552 32732 11558
rect 32680 11494 32732 11500
rect 31760 11348 31812 11354
rect 32784 11336 32812 11630
rect 32864 11348 32916 11354
rect 32784 11308 32864 11336
rect 31760 11290 31812 11296
rect 33244 11336 33272 11630
rect 33612 11626 33640 12260
rect 34348 12170 34376 13262
rect 34624 12714 34652 13942
rect 34704 13728 34756 13734
rect 34704 13670 34756 13676
rect 34716 13258 34744 13670
rect 34704 13252 34756 13258
rect 34704 13194 34756 13200
rect 34612 12708 34664 12714
rect 34612 12650 34664 12656
rect 34336 12164 34388 12170
rect 34336 12106 34388 12112
rect 34808 11898 34836 14282
rect 35084 13870 35112 14350
rect 35072 13864 35124 13870
rect 35072 13806 35124 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12102 35388 16050
rect 35440 15428 35492 15434
rect 35440 15370 35492 15376
rect 35452 15042 35480 15370
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 36004 15162 36032 17138
rect 36188 16522 36216 17546
rect 36648 17338 36676 18702
rect 37108 18698 37136 21966
rect 37476 20534 37504 22510
rect 37568 22234 37596 22578
rect 37556 22228 37608 22234
rect 37556 22170 37608 22176
rect 37556 21956 37608 21962
rect 37556 21898 37608 21904
rect 37568 21146 37596 21898
rect 37556 21140 37608 21146
rect 37556 21082 37608 21088
rect 37660 20534 37688 23054
rect 37844 22778 37872 25094
rect 37936 24138 37964 25230
rect 37924 24132 37976 24138
rect 37924 24074 37976 24080
rect 37936 23866 37964 24074
rect 37924 23860 37976 23866
rect 37924 23802 37976 23808
rect 37924 23112 37976 23118
rect 37924 23054 37976 23060
rect 37936 22778 37964 23054
rect 37832 22772 37884 22778
rect 37832 22714 37884 22720
rect 37924 22772 37976 22778
rect 37924 22714 37976 22720
rect 38028 22710 38056 26454
rect 38108 22976 38160 22982
rect 38108 22918 38160 22924
rect 38016 22704 38068 22710
rect 38016 22646 38068 22652
rect 38028 22094 38056 22646
rect 38120 22438 38148 22918
rect 38384 22704 38436 22710
rect 38384 22646 38436 22652
rect 38108 22432 38160 22438
rect 38108 22374 38160 22380
rect 38028 22066 38148 22094
rect 37924 21072 37976 21078
rect 37924 21014 37976 21020
rect 37832 20936 37884 20942
rect 37832 20878 37884 20884
rect 37740 20868 37792 20874
rect 37740 20810 37792 20816
rect 37464 20528 37516 20534
rect 37464 20470 37516 20476
rect 37648 20528 37700 20534
rect 37648 20470 37700 20476
rect 37372 19304 37424 19310
rect 37372 19246 37424 19252
rect 37280 18896 37332 18902
rect 37280 18838 37332 18844
rect 37096 18692 37148 18698
rect 37096 18634 37148 18640
rect 37108 17882 37136 18634
rect 37292 18630 37320 18838
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 37384 18426 37412 19246
rect 37476 18766 37504 20470
rect 37464 18760 37516 18766
rect 37464 18702 37516 18708
rect 37372 18420 37424 18426
rect 37372 18362 37424 18368
rect 37096 17876 37148 17882
rect 37096 17818 37148 17824
rect 37660 17542 37688 20470
rect 37752 18902 37780 20810
rect 37844 20602 37872 20878
rect 37832 20596 37884 20602
rect 37832 20538 37884 20544
rect 37936 19922 37964 21014
rect 38120 20942 38148 22066
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 20942 38240 21286
rect 38396 20942 38424 22646
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 38384 20936 38436 20942
rect 38384 20878 38436 20884
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 38396 19310 38424 20878
rect 38384 19304 38436 19310
rect 38384 19246 38436 19252
rect 37740 18896 37792 18902
rect 37740 18838 37792 18844
rect 37648 17536 37700 17542
rect 37648 17478 37700 17484
rect 36636 17332 36688 17338
rect 36636 17274 36688 17280
rect 36176 16516 36228 16522
rect 36176 16458 36228 16464
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 36636 15360 36688 15366
rect 36636 15302 36688 15308
rect 35992 15156 36044 15162
rect 35992 15098 36044 15104
rect 35452 15014 35572 15042
rect 36648 15026 36676 15302
rect 35440 14952 35492 14958
rect 35440 14894 35492 14900
rect 35452 14618 35480 14894
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 35544 14498 35572 15014
rect 36636 15020 36688 15026
rect 36636 14962 36688 14968
rect 36084 14884 36136 14890
rect 36084 14826 36136 14832
rect 35452 14470 35572 14498
rect 35452 13938 35480 14470
rect 35992 14408 36044 14414
rect 35992 14350 36044 14356
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 36004 14074 36032 14350
rect 36096 14346 36124 14826
rect 37292 14822 37320 15438
rect 38476 15360 38528 15366
rect 38476 15302 38528 15308
rect 37464 15088 37516 15094
rect 38488 15065 38516 15302
rect 37464 15030 37516 15036
rect 38474 15056 38530 15065
rect 36544 14816 36596 14822
rect 36544 14758 36596 14764
rect 37280 14816 37332 14822
rect 37280 14758 37332 14764
rect 36360 14408 36412 14414
rect 36360 14350 36412 14356
rect 36084 14340 36136 14346
rect 36084 14282 36136 14288
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 36372 14006 36400 14350
rect 36360 14000 36412 14006
rect 36360 13942 36412 13948
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35992 13932 36044 13938
rect 35992 13874 36044 13880
rect 36084 13932 36136 13938
rect 36084 13874 36136 13880
rect 35440 13728 35492 13734
rect 35440 13670 35492 13676
rect 35452 12986 35480 13670
rect 36004 13530 36032 13874
rect 35992 13524 36044 13530
rect 35992 13466 36044 13472
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35440 12980 35492 12986
rect 35440 12922 35492 12928
rect 36004 12238 36032 13330
rect 36096 12850 36124 13874
rect 36176 13524 36228 13530
rect 36176 13466 36228 13472
rect 36188 12850 36216 13466
rect 36372 12986 36400 13942
rect 36360 12980 36412 12986
rect 36360 12922 36412 12928
rect 36084 12844 36136 12850
rect 36084 12786 36136 12792
rect 36176 12844 36228 12850
rect 36176 12786 36228 12792
rect 36084 12368 36136 12374
rect 36084 12310 36136 12316
rect 35992 12232 36044 12238
rect 35992 12174 36044 12180
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 35348 11824 35400 11830
rect 35400 11784 35480 11812
rect 35348 11766 35400 11772
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 33600 11620 33652 11626
rect 33600 11562 33652 11568
rect 33612 11354 33640 11562
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 32864 11290 32916 11296
rect 32968 11308 33272 11336
rect 32968 11234 32996 11308
rect 32876 11206 32996 11234
rect 32876 11150 32904 11206
rect 33244 11150 33272 11308
rect 33600 11348 33652 11354
rect 33600 11290 33652 11296
rect 32864 11144 32916 11150
rect 32864 11086 32916 11092
rect 32956 11144 33008 11150
rect 32956 11086 33008 11092
rect 33232 11144 33284 11150
rect 33232 11086 33284 11092
rect 32588 11008 32640 11014
rect 32588 10950 32640 10956
rect 32600 10606 32628 10950
rect 32968 10742 32996 11086
rect 33140 10804 33192 10810
rect 33140 10746 33192 10752
rect 32956 10736 33008 10742
rect 32956 10678 33008 10684
rect 33152 10674 33180 10746
rect 33140 10668 33192 10674
rect 33140 10610 33192 10616
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 33244 10470 33272 11086
rect 33324 11008 33376 11014
rect 33324 10950 33376 10956
rect 33336 10674 33364 10950
rect 33612 10674 33640 11290
rect 33876 11144 33928 11150
rect 33876 11086 33928 11092
rect 33888 10674 33916 11086
rect 33968 10804 34020 10810
rect 33968 10746 34020 10752
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 33600 10668 33652 10674
rect 33600 10610 33652 10616
rect 33876 10668 33928 10674
rect 33876 10610 33928 10616
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32772 10464 32824 10470
rect 32772 10406 32824 10412
rect 32956 10464 33008 10470
rect 32956 10406 33008 10412
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 31576 10056 31628 10062
rect 31576 9998 31628 10004
rect 29644 9716 29696 9722
rect 29644 9658 29696 9664
rect 29748 9586 29776 9998
rect 31484 9988 31536 9994
rect 31484 9930 31536 9936
rect 30932 9920 30984 9926
rect 30932 9862 30984 9868
rect 30944 9636 30972 9862
rect 31496 9722 31524 9930
rect 31668 9920 31720 9926
rect 31668 9862 31720 9868
rect 32128 9920 32180 9926
rect 32128 9862 32180 9868
rect 31680 9722 31708 9862
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 31668 9716 31720 9722
rect 31668 9658 31720 9664
rect 31024 9648 31076 9654
rect 30944 9608 31024 9636
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 28356 9580 28408 9586
rect 28356 9522 28408 9528
rect 29092 9580 29144 9586
rect 29092 9522 29144 9528
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 28184 9178 28212 9522
rect 28368 9178 28396 9522
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28632 8560 28684 8566
rect 28632 8502 28684 8508
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28276 8022 28304 8434
rect 28264 8016 28316 8022
rect 28264 7958 28316 7964
rect 28644 7886 28672 8502
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 27528 7404 27580 7410
rect 27528 7346 27580 7352
rect 27436 7268 27488 7274
rect 27436 7210 27488 7216
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25424 6390 25452 6666
rect 25412 6384 25464 6390
rect 25412 6326 25464 6332
rect 25516 6322 25544 7142
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 26068 6458 26096 6734
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25964 6316 26016 6322
rect 25964 6258 26016 6264
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24676 5636 24728 5642
rect 24676 5578 24728 5584
rect 24780 5386 24808 6190
rect 24872 5574 24900 6258
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5710 25084 6054
rect 25136 5840 25188 5846
rect 25136 5782 25188 5788
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 24308 5364 24360 5370
rect 24780 5358 24900 5386
rect 24308 5306 24360 5312
rect 24872 5302 24900 5358
rect 24860 5296 24912 5302
rect 24860 5238 24912 5244
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23768 4486 23796 4626
rect 23952 4622 23980 5170
rect 24492 5092 24544 5098
rect 24492 5034 24544 5040
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23860 4214 23888 4422
rect 23952 4214 23980 4558
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 23848 4208 23900 4214
rect 23848 4150 23900 4156
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 23756 4004 23808 4010
rect 23756 3946 23808 3952
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23768 3466 23796 3946
rect 24044 3738 24072 4082
rect 24124 4004 24176 4010
rect 24124 3946 24176 3952
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24136 3641 24164 3946
rect 24122 3632 24178 3641
rect 24320 3602 24348 4218
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24122 3567 24178 3576
rect 24308 3596 24360 3602
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23756 3460 23808 3466
rect 23756 3402 23808 3408
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 23032 2990 23060 3402
rect 23768 3126 23796 3402
rect 23756 3120 23808 3126
rect 23756 3062 23808 3068
rect 24136 3058 24164 3567
rect 24308 3538 24360 3544
rect 24320 3097 24348 3538
rect 24306 3088 24362 3097
rect 24124 3052 24176 3058
rect 24306 3023 24308 3032
rect 24124 2994 24176 3000
rect 24360 3023 24362 3032
rect 24308 2994 24360 3000
rect 23020 2984 23072 2990
rect 23020 2926 23072 2932
rect 24412 2854 24440 4082
rect 24504 3534 24532 5034
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24872 4078 24900 4558
rect 25056 4078 25084 5510
rect 25148 5302 25176 5782
rect 25240 5642 25268 6258
rect 25332 5778 25360 6258
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 25228 5636 25280 5642
rect 25228 5578 25280 5584
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 25608 5302 25636 5578
rect 25976 5574 26004 6258
rect 26068 5710 26096 6394
rect 26160 6322 26188 6734
rect 27264 6458 27292 6802
rect 27448 6730 27476 7210
rect 27436 6724 27488 6730
rect 27436 6666 27488 6672
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 27448 6390 27476 6666
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26792 6316 26844 6322
rect 26792 6258 26844 6264
rect 26804 6186 26832 6258
rect 26792 6180 26844 6186
rect 26792 6122 26844 6128
rect 26424 6112 26476 6118
rect 26424 6054 26476 6060
rect 26436 5710 26464 6054
rect 26804 5914 26832 6122
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26424 5704 26476 5710
rect 27344 5704 27396 5710
rect 26424 5646 26476 5652
rect 27264 5664 27344 5692
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 25136 5296 25188 5302
rect 25136 5238 25188 5244
rect 25596 5296 25648 5302
rect 25596 5238 25648 5244
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 25240 4826 25268 5170
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 25332 4146 25360 4558
rect 25424 4282 25452 5102
rect 25976 5098 26004 5510
rect 25964 5092 26016 5098
rect 25964 5034 26016 5040
rect 25780 5024 25832 5030
rect 25780 4966 25832 4972
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 24676 4004 24728 4010
rect 24676 3946 24728 3952
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24688 3482 24716 3946
rect 24872 3670 24900 4014
rect 24860 3664 24912 3670
rect 24766 3632 24822 3641
rect 24860 3606 24912 3612
rect 25332 3602 25360 4082
rect 25424 3738 25452 4218
rect 25792 4214 25820 4966
rect 26240 4752 26292 4758
rect 26292 4700 26372 4706
rect 26240 4694 26372 4700
rect 26252 4678 26372 4694
rect 26436 4690 26464 5646
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26252 4282 26280 4422
rect 26344 4282 26372 4678
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 26700 4616 26752 4622
rect 26884 4616 26936 4622
rect 26752 4576 26832 4604
rect 26700 4558 26752 4564
rect 26608 4480 26660 4486
rect 26608 4422 26660 4428
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 25780 4208 25832 4214
rect 25780 4150 25832 4156
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25412 3732 25464 3738
rect 25412 3674 25464 3680
rect 24766 3567 24768 3576
rect 24820 3567 24822 3576
rect 25320 3596 25372 3602
rect 24768 3538 24820 3544
rect 25320 3538 25372 3544
rect 25700 3534 25728 4082
rect 26620 3942 26648 4422
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26422 3632 26478 3641
rect 26422 3567 26478 3576
rect 26436 3534 26464 3567
rect 25688 3528 25740 3534
rect 24688 3466 25084 3482
rect 25688 3470 25740 3476
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 24688 3460 25096 3466
rect 24688 3454 25044 3460
rect 25044 3402 25096 3408
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 3058 24808 3334
rect 25608 3194 25636 3402
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 26252 3097 26280 3470
rect 26620 3194 26648 3878
rect 26804 3398 26832 4576
rect 26884 4558 26936 4564
rect 26896 4214 26924 4558
rect 26976 4548 27028 4554
rect 27172 4536 27200 5578
rect 27028 4508 27200 4536
rect 26976 4490 27028 4496
rect 26884 4208 26936 4214
rect 26884 4150 26936 4156
rect 26896 3602 26924 4150
rect 27172 4049 27200 4508
rect 27264 4486 27292 5664
rect 27344 5646 27396 5652
rect 27448 4622 27476 6326
rect 27540 5522 27568 7346
rect 27816 7002 27844 7822
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 29104 6798 29132 9318
rect 29748 8974 29776 9522
rect 30944 9382 30972 9608
rect 31024 9590 31076 9596
rect 31024 9512 31076 9518
rect 31024 9454 31076 9460
rect 30932 9376 30984 9382
rect 30932 9318 30984 9324
rect 31036 9178 31064 9454
rect 31024 9172 31076 9178
rect 31024 9114 31076 9120
rect 31300 9036 31352 9042
rect 31300 8978 31352 8984
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 29748 8634 29776 8910
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 30116 8022 30144 8910
rect 31312 8634 31340 8978
rect 31680 8634 31708 9658
rect 32140 9586 32168 9862
rect 32324 9586 32352 10406
rect 32404 10192 32456 10198
rect 32404 10134 32456 10140
rect 32416 9586 32444 10134
rect 32784 9586 32812 10406
rect 32128 9580 32180 9586
rect 32128 9522 32180 9528
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32692 9450 32720 9522
rect 32680 9444 32732 9450
rect 32680 9386 32732 9392
rect 32692 9178 32720 9386
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 31760 8968 31812 8974
rect 31760 8910 31812 8916
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31668 8628 31720 8634
rect 31668 8570 31720 8576
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 31128 8090 31156 8434
rect 31312 8294 31340 8570
rect 31772 8362 31800 8910
rect 31864 8634 31892 8910
rect 31852 8628 31904 8634
rect 31852 8570 31904 8576
rect 31760 8356 31812 8362
rect 31760 8298 31812 8304
rect 31300 8288 31352 8294
rect 31300 8230 31352 8236
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 30104 8016 30156 8022
rect 30104 7958 30156 7964
rect 31772 7886 31800 8298
rect 31392 7880 31444 7886
rect 31312 7840 31392 7868
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 30380 7812 30432 7818
rect 30380 7754 30432 7760
rect 29092 6792 29144 6798
rect 29092 6734 29144 6740
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 27724 5914 27752 6190
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 27540 5494 27660 5522
rect 27632 4826 27660 5494
rect 28172 5160 28224 5166
rect 28172 5102 28224 5108
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 27264 4282 27292 4422
rect 27252 4276 27304 4282
rect 27252 4218 27304 4224
rect 27158 4040 27214 4049
rect 27158 3975 27214 3984
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 27448 3534 27476 4558
rect 27632 4554 27660 4762
rect 27804 4752 27856 4758
rect 27804 4694 27856 4700
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27620 4548 27672 4554
rect 27620 4490 27672 4496
rect 27540 4078 27568 4490
rect 27816 4214 27844 4694
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27804 4208 27856 4214
rect 27804 4150 27856 4156
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27712 4004 27764 4010
rect 27712 3946 27764 3952
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27632 3534 27660 3878
rect 27724 3534 27752 3946
rect 27908 3738 27936 4626
rect 28184 4622 28212 5102
rect 28632 5024 28684 5030
rect 28632 4966 28684 4972
rect 28644 4690 28672 4966
rect 28632 4684 28684 4690
rect 28632 4626 28684 4632
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28080 4480 28132 4486
rect 28080 4422 28132 4428
rect 28092 4162 28120 4422
rect 28184 4282 28212 4558
rect 28644 4282 28672 4626
rect 28724 4548 28776 4554
rect 28724 4490 28776 4496
rect 28172 4276 28224 4282
rect 28172 4218 28224 4224
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 28092 4134 28212 4162
rect 28184 3942 28212 4134
rect 28172 3936 28224 3942
rect 28172 3878 28224 3884
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 26792 3392 26844 3398
rect 26792 3334 26844 3340
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26238 3088 26294 3097
rect 24768 3052 24820 3058
rect 26804 3058 26832 3334
rect 26238 3023 26294 3032
rect 26792 3052 26844 3058
rect 24768 2994 24820 3000
rect 26792 2994 26844 3000
rect 26988 2922 27016 3470
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 27080 3058 27108 3402
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27172 3058 27200 3334
rect 27724 3194 27752 3470
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 28184 2990 28212 3878
rect 28736 3534 28764 4490
rect 29012 4010 29040 6258
rect 29196 5166 29224 7754
rect 30392 7002 30420 7754
rect 30380 6996 30432 7002
rect 30380 6938 30432 6944
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29288 6458 29316 6734
rect 29368 6656 29420 6662
rect 29368 6598 29420 6604
rect 29276 6452 29328 6458
rect 29276 6394 29328 6400
rect 29380 6322 29408 6598
rect 31312 6390 31340 7840
rect 31392 7822 31444 7828
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31944 7744 31996 7750
rect 31944 7686 31996 7692
rect 31956 7342 31984 7686
rect 32968 7410 32996 10406
rect 33416 9376 33468 9382
rect 33416 9318 33468 9324
rect 33428 7410 33456 9318
rect 33980 9110 34008 10746
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 34348 9722 34376 9862
rect 34336 9716 34388 9722
rect 34336 9658 34388 9664
rect 34440 9518 34468 11494
rect 34808 11014 34836 11698
rect 35348 11620 35400 11626
rect 35348 11562 35400 11568
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11008 34848 11014
rect 34796 10950 34848 10956
rect 34704 10804 34756 10810
rect 34704 10746 34756 10752
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 34532 10266 34560 10610
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 34520 10260 34572 10266
rect 34520 10202 34572 10208
rect 34428 9512 34480 9518
rect 34428 9454 34480 9460
rect 33968 9104 34020 9110
rect 33968 9046 34020 9052
rect 33980 8566 34008 9046
rect 34532 9042 34560 10202
rect 34624 10198 34652 10406
rect 34612 10192 34664 10198
rect 34612 10134 34664 10140
rect 34612 10056 34664 10062
rect 34612 9998 34664 10004
rect 34624 9722 34652 9998
rect 34612 9716 34664 9722
rect 34612 9658 34664 9664
rect 34612 9512 34664 9518
rect 34610 9480 34612 9489
rect 34664 9480 34666 9489
rect 34610 9415 34666 9424
rect 34716 9382 34744 10746
rect 34808 10674 34836 10950
rect 35360 10810 35388 11562
rect 35348 10804 35400 10810
rect 35348 10746 35400 10752
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34704 9376 34756 9382
rect 34704 9318 34756 9324
rect 34808 9364 34836 10610
rect 35348 10464 35400 10470
rect 35348 10406 35400 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34980 10260 35032 10266
rect 34980 10202 35032 10208
rect 34992 9586 35020 10202
rect 34980 9580 35032 9586
rect 34980 9522 35032 9528
rect 34992 9450 35020 9522
rect 34980 9444 35032 9450
rect 34980 9386 35032 9392
rect 34888 9376 34940 9382
rect 34808 9336 34888 9364
rect 34520 9036 34572 9042
rect 34520 8978 34572 8984
rect 34716 8974 34744 9318
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34336 8900 34388 8906
rect 34336 8842 34388 8848
rect 33968 8560 34020 8566
rect 33968 8502 34020 8508
rect 34348 8498 34376 8842
rect 34336 8492 34388 8498
rect 34336 8434 34388 8440
rect 34612 8424 34664 8430
rect 34612 8366 34664 8372
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 34440 7954 34468 8230
rect 33784 7948 33836 7954
rect 33784 7890 33836 7896
rect 34428 7948 34480 7954
rect 34428 7890 34480 7896
rect 33508 7744 33560 7750
rect 33508 7686 33560 7692
rect 33520 7410 33548 7686
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 32956 7404 33008 7410
rect 32956 7346 33008 7352
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 33416 7404 33468 7410
rect 33416 7346 33468 7352
rect 33508 7404 33560 7410
rect 33508 7346 33560 7352
rect 33692 7404 33744 7410
rect 33692 7346 33744 7352
rect 31944 7336 31996 7342
rect 31944 7278 31996 7284
rect 31956 6798 31984 7278
rect 31944 6792 31996 6798
rect 31944 6734 31996 6740
rect 32324 6730 32352 7346
rect 32680 7268 32732 7274
rect 32680 7210 32732 7216
rect 32692 6798 32720 7210
rect 32968 6798 32996 7346
rect 33152 6866 33180 7346
rect 33416 7200 33468 7206
rect 33416 7142 33468 7148
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33428 6798 33456 7142
rect 33520 6798 33548 7346
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32956 6792 33008 6798
rect 32956 6734 33008 6740
rect 33416 6792 33468 6798
rect 33416 6734 33468 6740
rect 33508 6792 33560 6798
rect 33508 6734 33560 6740
rect 33704 6730 33732 7346
rect 33796 6798 33824 7890
rect 33784 6792 33836 6798
rect 33784 6734 33836 6740
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 32312 6724 32364 6730
rect 32312 6666 32364 6672
rect 33324 6724 33376 6730
rect 33324 6666 33376 6672
rect 33692 6724 33744 6730
rect 33692 6666 33744 6672
rect 31300 6384 31352 6390
rect 31300 6326 31352 6332
rect 31852 6384 31904 6390
rect 31852 6326 31904 6332
rect 29368 6316 29420 6322
rect 29368 6258 29420 6264
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 31576 6316 31628 6322
rect 31576 6258 31628 6264
rect 30668 5914 30696 6258
rect 31588 6186 31616 6258
rect 31576 6180 31628 6186
rect 31576 6122 31628 6128
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 29736 5636 29788 5642
rect 29736 5578 29788 5584
rect 29828 5636 29880 5642
rect 29828 5578 29880 5584
rect 29748 5370 29776 5578
rect 29840 5370 29868 5578
rect 31588 5370 31616 6122
rect 31864 5710 31892 6326
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 32048 5710 32076 6054
rect 32324 5914 32352 6666
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 32416 6322 32444 6598
rect 33336 6458 33364 6666
rect 33324 6452 33376 6458
rect 33324 6394 33376 6400
rect 32404 6316 32456 6322
rect 32404 6258 32456 6264
rect 32772 6316 32824 6322
rect 32772 6258 32824 6264
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 32312 5908 32364 5914
rect 32312 5850 32364 5856
rect 32416 5710 32444 6258
rect 32784 5710 32812 6258
rect 33152 5914 33180 6258
rect 33324 6248 33376 6254
rect 33324 6190 33376 6196
rect 33140 5908 33192 5914
rect 33140 5850 33192 5856
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 32036 5704 32088 5710
rect 32036 5646 32088 5652
rect 32404 5704 32456 5710
rect 32404 5646 32456 5652
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 32784 5370 32812 5646
rect 33336 5370 33364 6190
rect 33888 5914 33916 6734
rect 34624 6610 34652 8366
rect 34716 8090 34744 8910
rect 34808 8430 34836 9336
rect 34888 9318 34940 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 9178 35388 10406
rect 35452 9994 35480 11784
rect 36096 11778 36124 12310
rect 35728 11762 36124 11778
rect 35716 11756 36124 11762
rect 35768 11750 36124 11756
rect 35716 11698 35768 11704
rect 36096 11354 36124 11750
rect 36188 11694 36216 12786
rect 36268 12776 36320 12782
rect 36268 12718 36320 12724
rect 36280 12442 36308 12718
rect 36268 12436 36320 12442
rect 36268 12378 36320 12384
rect 36176 11688 36228 11694
rect 36176 11630 36228 11636
rect 36188 11354 36216 11630
rect 36280 11354 36308 12378
rect 36556 12374 36584 14758
rect 36728 14408 36780 14414
rect 36728 14350 36780 14356
rect 36636 14340 36688 14346
rect 36636 14282 36688 14288
rect 36648 14074 36676 14282
rect 36636 14068 36688 14074
rect 36636 14010 36688 14016
rect 36740 13394 36768 14350
rect 37476 14346 37504 15030
rect 38474 14991 38530 15000
rect 37464 14340 37516 14346
rect 37464 14282 37516 14288
rect 37372 14272 37424 14278
rect 37372 14214 37424 14220
rect 37384 14074 37412 14214
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 37280 13796 37332 13802
rect 37280 13738 37332 13744
rect 36728 13388 36780 13394
rect 36728 13330 36780 13336
rect 37004 13252 37056 13258
rect 37004 13194 37056 13200
rect 37016 12986 37044 13194
rect 37004 12980 37056 12986
rect 37004 12922 37056 12928
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 36648 12646 36676 12786
rect 37292 12782 37320 13738
rect 37476 13258 37504 14282
rect 37464 13252 37516 13258
rect 37464 13194 37516 13200
rect 37004 12776 37056 12782
rect 37004 12718 37056 12724
rect 37280 12776 37332 12782
rect 37280 12718 37332 12724
rect 36636 12640 36688 12646
rect 36636 12582 36688 12588
rect 37016 12434 37044 12718
rect 37292 12434 37320 12718
rect 37016 12406 37136 12434
rect 37292 12406 37412 12434
rect 36544 12368 36596 12374
rect 36544 12310 36596 12316
rect 37108 12238 37136 12406
rect 36544 12232 36596 12238
rect 37096 12232 37148 12238
rect 36596 12192 36676 12220
rect 36544 12174 36596 12180
rect 36360 12096 36412 12102
rect 36360 12038 36412 12044
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 36372 11762 36400 12038
rect 36464 11830 36492 12038
rect 36452 11824 36504 11830
rect 36452 11766 36504 11772
rect 36360 11756 36412 11762
rect 36360 11698 36412 11704
rect 36084 11348 36136 11354
rect 36084 11290 36136 11296
rect 36176 11348 36228 11354
rect 36176 11290 36228 11296
rect 36268 11348 36320 11354
rect 36268 11290 36320 11296
rect 36268 11144 36320 11150
rect 36268 11086 36320 11092
rect 36084 11076 36136 11082
rect 36084 11018 36136 11024
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 36096 10538 36124 11018
rect 36176 11008 36228 11014
rect 36176 10950 36228 10956
rect 36188 10742 36216 10950
rect 36176 10736 36228 10742
rect 36176 10678 36228 10684
rect 36188 10606 36216 10678
rect 36176 10600 36228 10606
rect 36176 10542 36228 10548
rect 36084 10532 36136 10538
rect 36084 10474 36136 10480
rect 36188 10146 36216 10542
rect 36096 10118 36216 10146
rect 35440 9988 35492 9994
rect 35440 9930 35492 9936
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 35440 9648 35492 9654
rect 35440 9590 35492 9596
rect 35452 9518 35480 9590
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35440 9512 35492 9518
rect 35440 9454 35492 9460
rect 35348 9172 35400 9178
rect 35348 9114 35400 9120
rect 35544 8974 35572 9522
rect 35624 9512 35676 9518
rect 35622 9480 35624 9489
rect 35808 9512 35860 9518
rect 35676 9480 35678 9489
rect 35808 9454 35860 9460
rect 35622 9415 35678 9424
rect 35820 9178 35848 9454
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 35532 8968 35584 8974
rect 35532 8910 35584 8916
rect 35912 8922 35940 9318
rect 35912 8894 36032 8922
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 35268 8634 35296 8774
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 35256 8628 35308 8634
rect 35308 8588 35388 8616
rect 35256 8570 35308 8576
rect 34796 8424 34848 8430
rect 34796 8366 34848 8372
rect 34796 8288 34848 8294
rect 34796 8230 34848 8236
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 34808 7886 34836 8230
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 35256 7880 35308 7886
rect 35360 7868 35388 8588
rect 36004 8498 36032 8894
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 35308 7840 35388 7868
rect 35256 7822 35308 7828
rect 36096 7750 36124 10118
rect 36176 9444 36228 9450
rect 36176 9386 36228 9392
rect 36188 9178 36216 9386
rect 36176 9172 36228 9178
rect 36176 9114 36228 9120
rect 36176 8832 36228 8838
rect 36176 8774 36228 8780
rect 35348 7744 35400 7750
rect 35348 7686 35400 7692
rect 35992 7744 36044 7750
rect 35992 7686 36044 7692
rect 36084 7744 36136 7750
rect 36084 7686 36136 7692
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6798 35388 7686
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 36004 7426 36032 7686
rect 35820 7398 36032 7426
rect 36096 7410 36124 7686
rect 36188 7410 36216 8774
rect 36280 7886 36308 11086
rect 36268 7880 36320 7886
rect 36268 7822 36320 7828
rect 36084 7404 36136 7410
rect 35820 7342 35848 7398
rect 36084 7346 36136 7352
rect 36176 7404 36228 7410
rect 36176 7346 36228 7352
rect 35808 7336 35860 7342
rect 35808 7278 35860 7284
rect 35716 7200 35768 7206
rect 35716 7142 35768 7148
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 35728 6746 35756 7142
rect 35820 6866 35848 7278
rect 36372 6866 36400 11698
rect 36648 11694 36676 12192
rect 37096 12174 37148 12180
rect 36820 12164 36872 12170
rect 36820 12106 36872 12112
rect 36728 11824 36780 11830
rect 36728 11766 36780 11772
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 36544 11552 36596 11558
rect 36544 11494 36596 11500
rect 36452 11008 36504 11014
rect 36452 10950 36504 10956
rect 36464 8974 36492 10950
rect 36556 10674 36584 11494
rect 36648 11150 36676 11630
rect 36636 11144 36688 11150
rect 36636 11086 36688 11092
rect 36544 10668 36596 10674
rect 36544 10610 36596 10616
rect 36556 9586 36584 10610
rect 36648 10062 36676 11086
rect 36740 10810 36768 11766
rect 36728 10804 36780 10810
rect 36728 10746 36780 10752
rect 36832 10470 36860 12106
rect 37004 12096 37056 12102
rect 37004 12038 37056 12044
rect 36912 11552 36964 11558
rect 36912 11494 36964 11500
rect 36924 11218 36952 11494
rect 37016 11218 37044 12038
rect 37108 11354 37136 12174
rect 37384 11558 37412 12406
rect 37476 12306 37504 13194
rect 37832 12640 37884 12646
rect 37832 12582 37884 12588
rect 37464 12300 37516 12306
rect 37464 12242 37516 12248
rect 37372 11552 37424 11558
rect 37372 11494 37424 11500
rect 37096 11348 37148 11354
rect 37096 11290 37148 11296
rect 36912 11212 36964 11218
rect 36912 11154 36964 11160
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 36912 10736 36964 10742
rect 36912 10678 36964 10684
rect 36924 10606 36952 10678
rect 37016 10674 37044 11154
rect 37004 10668 37056 10674
rect 37004 10610 37056 10616
rect 37188 10668 37240 10674
rect 37188 10610 37240 10616
rect 36912 10600 36964 10606
rect 36912 10542 36964 10548
rect 36820 10464 36872 10470
rect 36820 10406 36872 10412
rect 36636 10056 36688 10062
rect 36636 9998 36688 10004
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36648 9042 36676 9998
rect 36832 9926 36860 10406
rect 36820 9920 36872 9926
rect 36820 9862 36872 9868
rect 36832 9586 36860 9862
rect 36924 9722 36952 10542
rect 36912 9716 36964 9722
rect 36912 9658 36964 9664
rect 36924 9586 36952 9658
rect 37200 9654 37228 10610
rect 37280 10464 37332 10470
rect 37280 10406 37332 10412
rect 37292 10130 37320 10406
rect 37384 10146 37412 11494
rect 37476 11082 37504 12242
rect 37844 11626 37872 12582
rect 37832 11620 37884 11626
rect 37832 11562 37884 11568
rect 37464 11076 37516 11082
rect 37464 11018 37516 11024
rect 37844 10538 37872 11562
rect 38384 10600 38436 10606
rect 38384 10542 38436 10548
rect 37832 10532 37884 10538
rect 37832 10474 37884 10480
rect 37280 10124 37332 10130
rect 37384 10118 37504 10146
rect 37280 10066 37332 10072
rect 37372 9988 37424 9994
rect 37372 9930 37424 9936
rect 37188 9648 37240 9654
rect 37188 9590 37240 9596
rect 36820 9580 36872 9586
rect 36820 9522 36872 9528
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 36728 9512 36780 9518
rect 36728 9454 36780 9460
rect 36740 9178 36768 9454
rect 36728 9172 36780 9178
rect 36728 9114 36780 9120
rect 36636 9036 36688 9042
rect 36636 8978 36688 8984
rect 36452 8968 36504 8974
rect 36452 8910 36504 8916
rect 36832 8022 36860 9522
rect 37004 9444 37056 9450
rect 37004 9386 37056 9392
rect 36912 8900 36964 8906
rect 36912 8842 36964 8848
rect 36924 8634 36952 8842
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 36544 8016 36596 8022
rect 36544 7958 36596 7964
rect 36820 8016 36872 8022
rect 36820 7958 36872 7964
rect 36556 7410 36584 7958
rect 37016 7818 37044 9386
rect 37292 8498 37320 9522
rect 37384 8906 37412 9930
rect 37476 9518 37504 10118
rect 38396 9926 38424 10542
rect 38384 9920 38436 9926
rect 38384 9862 38436 9868
rect 37464 9512 37516 9518
rect 37464 9454 37516 9460
rect 37372 8900 37424 8906
rect 37372 8842 37424 8848
rect 37384 8786 37412 8842
rect 37384 8758 37504 8786
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37292 8090 37320 8434
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 37292 7886 37320 8026
rect 37280 7880 37332 7886
rect 37280 7822 37332 7828
rect 37004 7812 37056 7818
rect 37004 7754 37056 7760
rect 37016 7478 37044 7754
rect 37372 7744 37424 7750
rect 37372 7686 37424 7692
rect 37004 7472 37056 7478
rect 37004 7414 37056 7420
rect 36452 7404 36504 7410
rect 36452 7346 36504 7352
rect 36544 7404 36596 7410
rect 36544 7346 36596 7352
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 36360 6860 36412 6866
rect 36360 6802 36412 6808
rect 35728 6718 36032 6746
rect 34532 6582 34652 6610
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 35440 6656 35492 6662
rect 35440 6598 35492 6604
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 34440 5914 34468 6190
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 34428 5908 34480 5914
rect 34428 5850 34480 5856
rect 34532 5710 34560 6582
rect 34808 6322 34836 6598
rect 35452 6390 35480 6598
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 35440 6384 35492 6390
rect 35440 6326 35492 6332
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 34624 5914 34652 6258
rect 35348 6248 35400 6254
rect 35348 6190 35400 6196
rect 34796 6180 34848 6186
rect 34796 6122 34848 6128
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34808 5778 34836 6122
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5772 34848 5778
rect 34796 5714 34848 5720
rect 35360 5710 35388 6190
rect 35452 5914 35480 6326
rect 36004 6322 36032 6718
rect 36464 6458 36492 7346
rect 37384 7002 37412 7686
rect 37372 6996 37424 7002
rect 37372 6938 37424 6944
rect 37476 6730 37504 8758
rect 38476 7948 38528 7954
rect 38476 7890 38528 7896
rect 37924 7880 37976 7886
rect 37924 7822 37976 7828
rect 37936 7546 37964 7822
rect 38384 7744 38436 7750
rect 38384 7686 38436 7692
rect 38396 7585 38424 7686
rect 38382 7576 38438 7585
rect 37924 7540 37976 7546
rect 38382 7511 38438 7520
rect 37924 7482 37976 7488
rect 38488 6866 38516 7890
rect 38476 6860 38528 6866
rect 38476 6802 38528 6808
rect 37464 6724 37516 6730
rect 37464 6666 37516 6672
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 35624 6316 35676 6322
rect 35992 6316 36044 6322
rect 35624 6258 35676 6264
rect 35820 6276 35992 6304
rect 35636 5914 35664 6258
rect 35440 5908 35492 5914
rect 35440 5850 35492 5856
rect 35624 5908 35676 5914
rect 35624 5850 35676 5856
rect 35820 5710 35848 6276
rect 35992 6258 36044 6264
rect 33784 5704 33836 5710
rect 33784 5646 33836 5652
rect 33876 5704 33928 5710
rect 33876 5646 33928 5652
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34704 5704 34756 5710
rect 34704 5646 34756 5652
rect 35072 5704 35124 5710
rect 35072 5646 35124 5652
rect 35348 5704 35400 5710
rect 35348 5646 35400 5652
rect 35808 5704 35860 5710
rect 35808 5646 35860 5652
rect 33796 5370 33824 5646
rect 29736 5364 29788 5370
rect 29736 5306 29788 5312
rect 29828 5364 29880 5370
rect 29828 5306 29880 5312
rect 31576 5364 31628 5370
rect 31576 5306 31628 5312
rect 32772 5364 32824 5370
rect 32772 5306 32824 5312
rect 33324 5364 33376 5370
rect 33324 5306 33376 5312
rect 33784 5364 33836 5370
rect 33784 5306 33836 5312
rect 29368 5228 29420 5234
rect 29368 5170 29420 5176
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 29380 4826 29408 5170
rect 29840 5098 29868 5306
rect 33140 5296 33192 5302
rect 33140 5238 33192 5244
rect 30840 5228 30892 5234
rect 30840 5170 30892 5176
rect 31576 5228 31628 5234
rect 31576 5170 31628 5176
rect 29828 5092 29880 5098
rect 29828 5034 29880 5040
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 30852 4758 30880 5170
rect 30840 4752 30892 4758
rect 30840 4694 30892 4700
rect 31588 4282 31616 5170
rect 31576 4276 31628 4282
rect 31576 4218 31628 4224
rect 30840 4208 30892 4214
rect 30840 4150 30892 4156
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 29092 4072 29144 4078
rect 29090 4040 29092 4049
rect 29184 4072 29236 4078
rect 29144 4040 29146 4049
rect 29000 4004 29052 4010
rect 29184 4014 29236 4020
rect 29090 3975 29146 3984
rect 29000 3946 29052 3952
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28552 2990 28580 3470
rect 29104 2990 29132 3975
rect 29196 3398 29224 4014
rect 29564 3670 29592 4082
rect 29840 3738 29868 4082
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30668 3738 30696 3878
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 30288 3732 30340 3738
rect 30288 3674 30340 3680
rect 30656 3732 30708 3738
rect 30656 3674 30708 3680
rect 29552 3664 29604 3670
rect 29552 3606 29604 3612
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 29748 3534 29776 3606
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 29184 3392 29236 3398
rect 29184 3334 29236 3340
rect 30116 3194 30144 3402
rect 30104 3188 30156 3194
rect 30104 3130 30156 3136
rect 30300 3126 30328 3674
rect 30748 3664 30800 3670
rect 30748 3606 30800 3612
rect 30564 3596 30616 3602
rect 30564 3538 30616 3544
rect 30288 3120 30340 3126
rect 30288 3062 30340 3068
rect 28172 2984 28224 2990
rect 28172 2926 28224 2932
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 26976 2916 27028 2922
rect 26976 2858 27028 2864
rect 30300 2854 30328 3062
rect 30576 2990 30604 3538
rect 30760 3398 30788 3606
rect 30852 3534 30880 4150
rect 31116 4140 31168 4146
rect 31036 4100 31116 4128
rect 30932 4072 30984 4078
rect 30932 4014 30984 4020
rect 30944 3618 30972 4014
rect 31036 3738 31064 4100
rect 31116 4082 31168 4088
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 32036 4140 32088 4146
rect 32036 4082 32088 4088
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 31128 3738 31156 3878
rect 31024 3732 31076 3738
rect 31024 3674 31076 3680
rect 31116 3732 31168 3738
rect 31116 3674 31168 3680
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 30944 3590 31064 3618
rect 31036 3534 31064 3590
rect 30840 3528 30892 3534
rect 30840 3470 30892 3476
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31312 3466 31340 3674
rect 31496 3534 31524 4082
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 31484 3528 31536 3534
rect 31484 3470 31536 3476
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30760 3058 30788 3334
rect 31312 3058 31340 3402
rect 30748 3052 30800 3058
rect 30748 2994 30800 3000
rect 30932 3052 30984 3058
rect 31300 3052 31352 3058
rect 30984 3012 31300 3040
rect 30932 2994 30984 3000
rect 31300 2994 31352 3000
rect 30564 2984 30616 2990
rect 30564 2926 30616 2932
rect 31404 2922 31432 3470
rect 31496 3058 31524 3470
rect 31588 3126 31616 4082
rect 32048 3738 32076 4082
rect 33152 4078 33180 5238
rect 33336 5234 33364 5306
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 33888 5098 33916 5646
rect 34716 5370 34744 5646
rect 35084 5370 35112 5646
rect 34704 5364 34756 5370
rect 34704 5306 34756 5312
rect 35072 5364 35124 5370
rect 35072 5306 35124 5312
rect 35360 5234 35388 5646
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34152 5228 34204 5234
rect 34152 5170 34204 5176
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 33876 5092 33928 5098
rect 33876 5034 33928 5040
rect 33888 4826 33916 5034
rect 34072 4826 34100 5102
rect 34164 4826 34192 5170
rect 33876 4820 33928 4826
rect 33876 4762 33928 4768
rect 34060 4820 34112 4826
rect 34060 4762 34112 4768
rect 34152 4820 34204 4826
rect 34152 4762 34204 4768
rect 33508 4684 33560 4690
rect 33508 4626 33560 4632
rect 33416 4616 33468 4622
rect 33416 4558 33468 4564
rect 33428 4282 33456 4558
rect 33520 4282 33548 4626
rect 34072 4554 34100 4762
rect 34808 4622 34836 5170
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35360 4826 35388 5170
rect 35348 4820 35400 4826
rect 35348 4762 35400 4768
rect 34796 4616 34848 4622
rect 34796 4558 34848 4564
rect 34060 4548 34112 4554
rect 34060 4490 34112 4496
rect 34704 4480 34756 4486
rect 34704 4422 34756 4428
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33508 4276 33560 4282
rect 33508 4218 33560 4224
rect 32312 4072 32364 4078
rect 32312 4014 32364 4020
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 32324 3738 32352 4014
rect 34716 3942 34744 4422
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 32312 3732 32364 3738
rect 32312 3674 32364 3680
rect 31668 3528 31720 3534
rect 31668 3470 31720 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 31576 3120 31628 3126
rect 31576 3062 31628 3068
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 31680 2990 31708 3470
rect 32324 3194 32352 3470
rect 32312 3188 32364 3194
rect 32312 3130 32364 3136
rect 31668 2984 31720 2990
rect 31668 2926 31720 2932
rect 31392 2916 31444 2922
rect 31392 2858 31444 2864
rect 34808 2854 34836 4558
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 38476 3528 38528 3534
rect 38474 3496 38476 3505
rect 38528 3496 38530 3505
rect 38474 3431 38530 3440
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 38476 2984 38528 2990
rect 38476 2926 38528 2932
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 34796 2848 34848 2854
rect 38488 2825 38516 2926
rect 34796 2790 34848 2796
rect 38474 2816 38530 2825
rect 21284 2746 21404 2774
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 21376 2446 21404 2746
rect 34934 2748 35242 2757
rect 38474 2751 38530 2760
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 14844 800 14872 2246
rect 21284 800 21312 2246
rect 23860 800 23888 2382
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 24504 800 24532 2246
rect 27080 800 27108 2246
rect 27724 800 27752 2246
rect 29012 800 29040 2246
rect 29656 800 29684 2382
rect 30300 800 30328 2382
rect 35452 800 35480 2382
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 2382
rect 38476 2304 38528 2310
rect 38476 2246 38528 2252
rect 38488 2145 38516 2246
rect 38474 2136 38530 2145
rect 38474 2071 38530 2080
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 35438 0 35494 800
rect 36082 0 36138 800
<< via2 >>
rect 38566 39480 38622 39536
rect 1306 37460 1362 37496
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1306 37440 1308 37460
rect 1308 37440 1360 37460
rect 1360 37440 1362 37460
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 846 36896 902 36952
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 846 36252 848 36272
rect 848 36252 900 36272
rect 900 36252 902 36272
rect 846 36216 902 36252
rect 846 35572 848 35592
rect 848 35572 900 35592
rect 900 35572 902 35592
rect 846 35536 902 35572
rect 846 34856 902 34912
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 110 33768 166 33824
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 846 30116 902 30152
rect 846 30096 848 30116
rect 848 30096 900 30116
rect 900 30096 902 30116
rect 846 29416 902 29472
rect 846 28736 902 28792
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 1306 25200 1362 25256
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4986 24284 4988 24304
rect 4988 24284 5040 24304
rect 5040 24284 5042 24304
rect 4986 24248 5042 24284
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 7654 24248 7710 24304
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1306 10920 1362 10976
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1306 10260 1362 10296
rect 1306 10240 1308 10260
rect 1308 10240 1360 10260
rect 1360 10240 1362 10260
rect 938 9560 994 9616
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 846 6704 902 6760
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 846 5344 902 5400
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 846 4936 902 4992
rect 846 4256 902 4312
rect 846 3612 848 3632
rect 848 3612 900 3632
rect 900 3612 902 3632
rect 846 3576 902 3612
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 846 2932 848 2952
rect 848 2932 900 2952
rect 900 2932 902 2952
rect 846 2896 902 2932
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 15842 27512 15898 27568
rect 23754 36116 23756 36136
rect 23756 36116 23808 36136
rect 23808 36116 23810 36136
rect 23754 36080 23810 36116
rect 17590 27548 17592 27568
rect 17592 27548 17644 27568
rect 17644 27548 17646 27568
rect 17590 27512 17646 27548
rect 18694 27512 18750 27568
rect 19154 27512 19210 27568
rect 17958 23840 18014 23896
rect 18418 24268 18474 24304
rect 18418 24248 18420 24268
rect 18420 24248 18472 24268
rect 18472 24248 18474 24268
rect 18418 24132 18474 24168
rect 18418 24112 18420 24132
rect 18420 24112 18472 24132
rect 18472 24112 18474 24132
rect 19154 24248 19210 24304
rect 19246 24132 19302 24168
rect 19246 24112 19248 24132
rect 19248 24112 19300 24132
rect 19300 24112 19302 24132
rect 19246 23860 19302 23896
rect 19246 23840 19248 23860
rect 19248 23840 19300 23860
rect 19300 23840 19302 23860
rect 14186 14340 14242 14376
rect 14186 14320 14188 14340
rect 14188 14320 14240 14340
rect 14240 14320 14242 14340
rect 20902 25064 20958 25120
rect 21270 24928 21326 24984
rect 21178 24520 21234 24576
rect 22282 24928 22338 24984
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37922 38800 37978 38856
rect 38290 38120 38346 38176
rect 38198 37460 38254 37496
rect 38198 37440 38200 37460
rect 38200 37440 38252 37460
rect 38252 37440 38254 37460
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 26146 36116 26148 36136
rect 26148 36116 26200 36136
rect 26200 36116 26202 36136
rect 26146 36080 26202 36116
rect 22650 25064 22706 25120
rect 21822 24520 21878 24576
rect 18510 19372 18566 19408
rect 18510 19352 18512 19372
rect 18512 19352 18564 19372
rect 18564 19352 18566 19372
rect 17314 16244 17370 16280
rect 17314 16224 17316 16244
rect 17316 16224 17368 16244
rect 17368 16224 17370 16244
rect 16578 13776 16634 13832
rect 17958 14728 18014 14784
rect 21914 20440 21970 20496
rect 38474 36760 38530 36816
rect 22282 20440 22338 20496
rect 19982 16360 20038 16416
rect 19246 14728 19302 14784
rect 18786 11464 18842 11520
rect 23294 20460 23350 20496
rect 26422 23060 26424 23080
rect 26424 23060 26476 23080
rect 26476 23060 26478 23080
rect 26422 23024 26478 23060
rect 23294 20440 23296 20460
rect 23296 20440 23348 20460
rect 23348 20440 23350 20460
rect 23110 14320 23166 14376
rect 21914 13776 21970 13832
rect 22466 10240 22522 10296
rect 23386 10104 23442 10160
rect 23110 9968 23166 10024
rect 23478 8492 23534 8528
rect 23478 8472 23480 8492
rect 23480 8472 23532 8492
rect 23532 8472 23534 8492
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 38474 36100 38530 36136
rect 38474 36080 38476 36100
rect 38476 36080 38528 36100
rect 38528 36080 38530 36100
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 38474 35436 38476 35456
rect 38476 35436 38528 35456
rect 38528 35436 38530 35456
rect 38474 35400 38530 35436
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 38474 34720 38530 34776
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 38474 34040 38530 34096
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 27526 23432 27582 23488
rect 28446 23060 28448 23080
rect 28448 23060 28500 23080
rect 28500 23060 28502 23080
rect 28446 23024 28502 23060
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 38474 33380 38530 33416
rect 38474 33360 38476 33380
rect 38476 33360 38528 33380
rect 38528 33360 38530 33380
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 38474 31320 38530 31376
rect 38474 30676 38476 30696
rect 38476 30676 38528 30696
rect 38528 30676 38530 30696
rect 38474 30640 38530 30676
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 30010 23432 30066 23488
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 31390 20884 31392 20904
rect 31392 20884 31444 20904
rect 31444 20884 31446 20904
rect 31390 20848 31446 20884
rect 33046 20868 33102 20904
rect 33046 20848 33048 20868
rect 33048 20848 33100 20868
rect 33100 20848 33102 20868
rect 23662 10260 23718 10296
rect 23662 10240 23664 10260
rect 23664 10240 23716 10260
rect 23716 10240 23718 10260
rect 23938 10260 23994 10296
rect 23938 10240 23940 10260
rect 23940 10240 23992 10260
rect 23992 10240 23994 10260
rect 23846 9832 23902 9888
rect 24122 10004 24124 10024
rect 24124 10004 24176 10024
rect 24176 10004 24178 10024
rect 24122 9968 24178 10004
rect 24214 9832 24270 9888
rect 24490 10104 24546 10160
rect 24858 10240 24914 10296
rect 24214 7948 24270 7984
rect 24214 7928 24216 7948
rect 24216 7928 24268 7948
rect 24268 7928 24270 7948
rect 30654 17040 30710 17096
rect 33046 20476 33048 20496
rect 33048 20476 33100 20496
rect 33100 20476 33102 20496
rect 33046 20440 33102 20476
rect 25226 8492 25282 8528
rect 25226 8472 25228 8492
rect 25228 8472 25280 8492
rect 25280 8472 25282 8492
rect 25226 7964 25228 7984
rect 25228 7964 25280 7984
rect 25280 7964 25282 7984
rect 25226 7928 25282 7964
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 38382 27240 38438 27296
rect 35990 20440 36046 20496
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 33414 17060 33470 17096
rect 33414 17040 33416 17060
rect 33416 17040 33468 17060
rect 33468 17040 33470 17060
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35990 19372 36046 19408
rect 35990 19352 35992 19372
rect 35992 19352 36044 19372
rect 36044 19352 36046 19372
rect 36818 19372 36874 19408
rect 36818 19352 36820 19372
rect 36820 19352 36872 19372
rect 36872 19352 36874 19372
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 24122 3576 24178 3632
rect 24306 3052 24362 3088
rect 24306 3032 24308 3052
rect 24308 3032 24360 3052
rect 24360 3032 24362 3052
rect 24766 3596 24822 3632
rect 24766 3576 24768 3596
rect 24768 3576 24820 3596
rect 24820 3576 24822 3596
rect 26422 3576 26478 3632
rect 27158 3984 27214 4040
rect 26238 3032 26294 3088
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34610 9460 34612 9480
rect 34612 9460 34664 9480
rect 34664 9460 34666 9480
rect 34610 9424 34666 9460
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 38474 15000 38530 15056
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 35622 9460 35624 9480
rect 35624 9460 35676 9480
rect 35676 9460 35678 9480
rect 35622 9424 35678 9460
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 38382 7520 38438 7576
rect 29090 4020 29092 4040
rect 29092 4020 29144 4040
rect 29144 4020 29146 4040
rect 29090 3984 29146 4020
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38474 3476 38476 3496
rect 38476 3476 38528 3496
rect 38528 3476 38530 3496
rect 38474 3440 38530 3476
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 38474 2760 38530 2816
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 38474 2080 38530 2136
<< metal3 >>
rect 38561 39538 38627 39541
rect 39200 39538 40000 39568
rect 38561 39536 40000 39538
rect 38561 39480 38566 39536
rect 38622 39480 40000 39536
rect 38561 39478 40000 39480
rect 38561 39475 38627 39478
rect 39200 39448 40000 39478
rect 37917 38858 37983 38861
rect 39200 38858 40000 38888
rect 37917 38856 40000 38858
rect 37917 38800 37922 38856
rect 37978 38800 40000 38856
rect 37917 38798 40000 38800
rect 37917 38795 37983 38798
rect 39200 38768 40000 38798
rect 38285 38178 38351 38181
rect 39200 38178 40000 38208
rect 38285 38176 40000 38178
rect 38285 38120 38290 38176
rect 38346 38120 40000 38176
rect 38285 38118 40000 38120
rect 38285 38115 38351 38118
rect 39200 38088 40000 38118
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 1301 37498 1367 37501
rect 0 37496 1367 37498
rect 0 37440 1306 37496
rect 1362 37440 1367 37496
rect 0 37438 1367 37440
rect 0 37408 800 37438
rect 1301 37435 1367 37438
rect 38193 37498 38259 37501
rect 39200 37498 40000 37528
rect 38193 37496 40000 37498
rect 38193 37440 38198 37496
rect 38254 37440 40000 37496
rect 38193 37438 40000 37440
rect 38193 37435 38259 37438
rect 39200 37408 40000 37438
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 841 36954 907 36957
rect 798 36952 907 36954
rect 798 36896 846 36952
rect 902 36896 907 36952
rect 798 36891 907 36896
rect 798 36848 858 36891
rect 0 36758 858 36848
rect 38469 36818 38535 36821
rect 39200 36818 40000 36848
rect 38469 36816 40000 36818
rect 38469 36760 38474 36816
rect 38530 36760 40000 36816
rect 38469 36758 40000 36760
rect 0 36728 800 36758
rect 38469 36755 38535 36758
rect 39200 36728 40000 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 841 36274 907 36277
rect 798 36272 907 36274
rect 798 36216 846 36272
rect 902 36216 907 36272
rect 798 36211 907 36216
rect 798 36168 858 36211
rect 0 36078 858 36168
rect 23749 36138 23815 36141
rect 26141 36138 26207 36141
rect 23749 36136 26207 36138
rect 23749 36080 23754 36136
rect 23810 36080 26146 36136
rect 26202 36080 26207 36136
rect 23749 36078 26207 36080
rect 0 36048 800 36078
rect 23749 36075 23815 36078
rect 26141 36075 26207 36078
rect 38469 36138 38535 36141
rect 39200 36138 40000 36168
rect 38469 36136 40000 36138
rect 38469 36080 38474 36136
rect 38530 36080 40000 36136
rect 38469 36078 40000 36080
rect 38469 36075 38535 36078
rect 39200 36048 40000 36078
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 841 35594 907 35597
rect 798 35592 907 35594
rect 798 35536 846 35592
rect 902 35536 907 35592
rect 798 35531 907 35536
rect 798 35488 858 35531
rect 0 35398 858 35488
rect 38469 35458 38535 35461
rect 39200 35458 40000 35488
rect 38469 35456 40000 35458
rect 38469 35400 38474 35456
rect 38530 35400 40000 35456
rect 38469 35398 40000 35400
rect 0 35368 800 35398
rect 38469 35395 38535 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 40000 35398
rect 34930 35327 35246 35328
rect 841 34914 907 34917
rect 798 34912 907 34914
rect 798 34856 846 34912
rect 902 34856 907 34912
rect 798 34851 907 34856
rect 798 34808 858 34851
rect 0 34718 858 34808
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 38469 34778 38535 34781
rect 39200 34778 40000 34808
rect 38469 34776 40000 34778
rect 38469 34720 38474 34776
rect 38530 34720 40000 34776
rect 38469 34718 40000 34720
rect 0 34688 800 34718
rect 38469 34715 38535 34718
rect 39200 34688 40000 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 38469 34098 38535 34101
rect 39200 34098 40000 34128
rect 0 34038 1042 34098
rect 0 34008 800 34038
rect 105 33826 171 33829
rect 982 33826 1042 34038
rect 38469 34096 40000 34098
rect 38469 34040 38474 34096
rect 38530 34040 40000 34096
rect 38469 34038 40000 34040
rect 38469 34035 38535 34038
rect 39200 34008 40000 34038
rect 105 33824 1042 33826
rect 105 33768 110 33824
rect 166 33768 1042 33824
rect 105 33766 1042 33768
rect 105 33763 171 33766
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 38469 33418 38535 33421
rect 39200 33418 40000 33448
rect 38469 33416 40000 33418
rect 38469 33360 38474 33416
rect 38530 33360 40000 33416
rect 38469 33358 40000 33360
rect 38469 33355 38535 33358
rect 39200 33328 40000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 38469 31378 38535 31381
rect 39200 31378 40000 31408
rect 38469 31376 40000 31378
rect 38469 31320 38474 31376
rect 38530 31320 40000 31376
rect 38469 31318 40000 31320
rect 38469 31315 38535 31318
rect 39200 31288 40000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 38469 30698 38535 30701
rect 39200 30698 40000 30728
rect 38469 30696 40000 30698
rect 38469 30640 38474 30696
rect 38530 30640 40000 30696
rect 38469 30638 40000 30640
rect 38469 30635 38535 30638
rect 39200 30608 40000 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 841 30154 907 30157
rect 798 30152 907 30154
rect 798 30096 846 30152
rect 902 30096 907 30152
rect 798 30091 907 30096
rect 798 30048 858 30091
rect 0 29958 858 30048
rect 0 29928 800 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 841 29474 907 29477
rect 798 29472 907 29474
rect 798 29416 846 29472
rect 902 29416 907 29472
rect 798 29411 907 29416
rect 798 29368 858 29411
rect 0 29278 858 29368
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 0 29248 800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 841 28794 907 28797
rect 798 28792 907 28794
rect 798 28736 846 28792
rect 902 28736 907 28792
rect 798 28731 907 28736
rect 798 28688 858 28731
rect 0 28598 858 28688
rect 0 28568 800 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 15837 27570 15903 27573
rect 17585 27570 17651 27573
rect 18689 27570 18755 27573
rect 19149 27570 19215 27573
rect 15837 27568 19215 27570
rect 15837 27512 15842 27568
rect 15898 27512 17590 27568
rect 17646 27512 18694 27568
rect 18750 27512 19154 27568
rect 19210 27512 19215 27568
rect 15837 27510 19215 27512
rect 15837 27507 15903 27510
rect 17585 27507 17651 27510
rect 18689 27507 18755 27510
rect 19149 27507 19215 27510
rect 38377 27298 38443 27301
rect 39200 27298 40000 27328
rect 38377 27296 40000 27298
rect 38377 27240 38382 27296
rect 38438 27240 40000 27296
rect 38377 27238 40000 27240
rect 38377 27235 38443 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 39200 27208 40000 27238
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 1301 25258 1367 25261
rect 0 25256 1367 25258
rect 0 25200 1306 25256
rect 1362 25200 1367 25256
rect 0 25198 1367 25200
rect 0 25168 800 25198
rect 1301 25195 1367 25198
rect 20897 25122 20963 25125
rect 22645 25122 22711 25125
rect 20897 25120 22711 25122
rect 20897 25064 20902 25120
rect 20958 25064 22650 25120
rect 22706 25064 22711 25120
rect 20897 25062 22711 25064
rect 20897 25059 20963 25062
rect 22645 25059 22711 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 21265 24986 21331 24989
rect 22277 24986 22343 24989
rect 21265 24984 22343 24986
rect 21265 24928 21270 24984
rect 21326 24928 22282 24984
rect 22338 24928 22343 24984
rect 21265 24926 22343 24928
rect 21265 24923 21331 24926
rect 22277 24923 22343 24926
rect 21173 24578 21239 24581
rect 21817 24578 21883 24581
rect 21173 24576 21883 24578
rect 21173 24520 21178 24576
rect 21234 24520 21822 24576
rect 21878 24520 21883 24576
rect 21173 24518 21883 24520
rect 21173 24515 21239 24518
rect 21817 24515 21883 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 4981 24306 5047 24309
rect 7649 24306 7715 24309
rect 4981 24304 7715 24306
rect 4981 24248 4986 24304
rect 5042 24248 7654 24304
rect 7710 24248 7715 24304
rect 4981 24246 7715 24248
rect 4981 24243 5047 24246
rect 7649 24243 7715 24246
rect 18413 24306 18479 24309
rect 19149 24306 19215 24309
rect 18413 24304 19215 24306
rect 18413 24248 18418 24304
rect 18474 24248 19154 24304
rect 19210 24248 19215 24304
rect 18413 24246 19215 24248
rect 18413 24243 18479 24246
rect 19149 24243 19215 24246
rect 18413 24170 18479 24173
rect 19241 24170 19307 24173
rect 18413 24168 19307 24170
rect 18413 24112 18418 24168
rect 18474 24112 19246 24168
rect 19302 24112 19307 24168
rect 18413 24110 19307 24112
rect 18413 24107 18479 24110
rect 19241 24107 19307 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 17953 23898 18019 23901
rect 19241 23898 19307 23901
rect 17953 23896 19307 23898
rect 17953 23840 17958 23896
rect 18014 23840 19246 23896
rect 19302 23840 19307 23896
rect 17953 23838 19307 23840
rect 17953 23835 18019 23838
rect 19241 23835 19307 23838
rect 27521 23490 27587 23493
rect 30005 23490 30071 23493
rect 27521 23488 30071 23490
rect 27521 23432 27526 23488
rect 27582 23432 30010 23488
rect 30066 23432 30071 23488
rect 27521 23430 30071 23432
rect 27521 23427 27587 23430
rect 30005 23427 30071 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 26417 23082 26483 23085
rect 28441 23082 28507 23085
rect 26417 23080 28507 23082
rect 26417 23024 26422 23080
rect 26478 23024 28446 23080
rect 28502 23024 28507 23080
rect 26417 23022 28507 23024
rect 26417 23019 26483 23022
rect 28441 23019 28507 23022
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 31385 20906 31451 20909
rect 33041 20906 33107 20909
rect 36118 20906 36124 20908
rect 31385 20904 36124 20906
rect 31385 20848 31390 20904
rect 31446 20848 33046 20904
rect 33102 20848 36124 20904
rect 31385 20846 36124 20848
rect 31385 20843 31451 20846
rect 33041 20843 33107 20846
rect 36118 20844 36124 20846
rect 36188 20844 36194 20908
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 21909 20498 21975 20501
rect 22277 20498 22343 20501
rect 23289 20498 23355 20501
rect 21909 20496 23355 20498
rect 21909 20440 21914 20496
rect 21970 20440 22282 20496
rect 22338 20440 23294 20496
rect 23350 20440 23355 20496
rect 21909 20438 23355 20440
rect 21909 20435 21975 20438
rect 22277 20435 22343 20438
rect 23289 20435 23355 20438
rect 33041 20498 33107 20501
rect 35985 20498 36051 20501
rect 33041 20496 36051 20498
rect 33041 20440 33046 20496
rect 33102 20440 35990 20496
rect 36046 20440 36051 20496
rect 33041 20438 36051 20440
rect 33041 20435 33107 20438
rect 35985 20435 36051 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 17902 19348 17908 19412
rect 17972 19410 17978 19412
rect 18505 19410 18571 19413
rect 17972 19408 18571 19410
rect 17972 19352 18510 19408
rect 18566 19352 18571 19408
rect 17972 19350 18571 19352
rect 17972 19348 17978 19350
rect 18505 19347 18571 19350
rect 35985 19410 36051 19413
rect 36118 19410 36124 19412
rect 35985 19408 36124 19410
rect 35985 19352 35990 19408
rect 36046 19352 36124 19408
rect 35985 19350 36124 19352
rect 35985 19347 36051 19350
rect 36118 19348 36124 19350
rect 36188 19410 36194 19412
rect 36813 19410 36879 19413
rect 36188 19408 36879 19410
rect 36188 19352 36818 19408
rect 36874 19352 36879 19408
rect 36188 19350 36879 19352
rect 36188 19348 36194 19350
rect 36813 19347 36879 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 30649 17098 30715 17101
rect 33409 17098 33475 17101
rect 30649 17096 33475 17098
rect 30649 17040 30654 17096
rect 30710 17040 33414 17096
rect 33470 17040 33475 17096
rect 30649 17038 33475 17040
rect 30649 17035 30715 17038
rect 33409 17035 33475 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19374 16356 19380 16420
rect 19444 16418 19450 16420
rect 19977 16418 20043 16421
rect 19444 16416 20043 16418
rect 19444 16360 19982 16416
rect 20038 16360 20043 16416
rect 19444 16358 20043 16360
rect 19444 16356 19450 16358
rect 19977 16355 20043 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 17309 16282 17375 16285
rect 17902 16282 17908 16284
rect 17309 16280 17908 16282
rect 17309 16224 17314 16280
rect 17370 16224 17908 16280
rect 17309 16222 17908 16224
rect 17309 16219 17375 16222
rect 17902 16220 17908 16222
rect 17972 16220 17978 16284
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 38469 15058 38535 15061
rect 39200 15058 40000 15088
rect 38469 15056 40000 15058
rect 38469 15000 38474 15056
rect 38530 15000 40000 15056
rect 38469 14998 40000 15000
rect 38469 14995 38535 14998
rect 39200 14968 40000 14998
rect 17953 14786 18019 14789
rect 19241 14786 19307 14789
rect 17953 14784 19307 14786
rect 17953 14728 17958 14784
rect 18014 14728 19246 14784
rect 19302 14728 19307 14784
rect 17953 14726 19307 14728
rect 17953 14723 18019 14726
rect 19241 14723 19307 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 14181 14378 14247 14381
rect 23105 14378 23171 14381
rect 14181 14376 23171 14378
rect 14181 14320 14186 14376
rect 14242 14320 23110 14376
rect 23166 14320 23171 14376
rect 14181 14318 23171 14320
rect 14181 14315 14247 14318
rect 23105 14315 23171 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 16573 13834 16639 13837
rect 21909 13834 21975 13837
rect 16573 13832 21975 13834
rect 16573 13776 16578 13832
rect 16634 13776 21914 13832
rect 21970 13776 21975 13832
rect 16573 13774 21975 13776
rect 16573 13771 16639 13774
rect 21909 13771 21975 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 18781 11522 18847 11525
rect 19374 11522 19380 11524
rect 18781 11520 19380 11522
rect 18781 11464 18786 11520
rect 18842 11464 19380 11520
rect 18781 11462 19380 11464
rect 18781 11459 18847 11462
rect 19374 11460 19380 11462
rect 19444 11460 19450 11524
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1301 10298 1367 10301
rect 0 10296 1367 10298
rect 0 10240 1306 10296
rect 1362 10240 1367 10296
rect 0 10238 1367 10240
rect 0 10208 800 10238
rect 1301 10235 1367 10238
rect 22461 10298 22527 10301
rect 23657 10298 23723 10301
rect 22461 10296 23723 10298
rect 22461 10240 22466 10296
rect 22522 10240 23662 10296
rect 23718 10240 23723 10296
rect 22461 10238 23723 10240
rect 22461 10235 22527 10238
rect 23657 10235 23723 10238
rect 23933 10298 23999 10301
rect 24853 10298 24919 10301
rect 23933 10296 24919 10298
rect 23933 10240 23938 10296
rect 23994 10240 24858 10296
rect 24914 10240 24919 10296
rect 23933 10238 24919 10240
rect 23933 10235 23999 10238
rect 24853 10235 24919 10238
rect 23381 10162 23447 10165
rect 24485 10162 24551 10165
rect 23381 10160 24551 10162
rect 23381 10104 23386 10160
rect 23442 10104 24490 10160
rect 24546 10104 24551 10160
rect 23381 10102 24551 10104
rect 23381 10099 23447 10102
rect 24485 10099 24551 10102
rect 23105 10026 23171 10029
rect 24117 10026 24183 10029
rect 23105 10024 24183 10026
rect 23105 9968 23110 10024
rect 23166 9968 24122 10024
rect 24178 9968 24183 10024
rect 23105 9966 24183 9968
rect 23105 9963 23171 9966
rect 24117 9963 24183 9966
rect 23841 9890 23907 9893
rect 24209 9890 24275 9893
rect 23841 9888 24275 9890
rect 23841 9832 23846 9888
rect 23902 9832 24214 9888
rect 24270 9832 24275 9888
rect 23841 9830 24275 9832
rect 23841 9827 23907 9830
rect 24209 9827 24275 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 0 9618 800 9648
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 800 9558
rect 933 9555 999 9558
rect 34605 9482 34671 9485
rect 35617 9482 35683 9485
rect 34605 9480 35683 9482
rect 34605 9424 34610 9480
rect 34666 9424 35622 9480
rect 35678 9424 35683 9480
rect 34605 9422 35683 9424
rect 34605 9419 34671 9422
rect 35617 9419 35683 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 23473 8530 23539 8533
rect 25221 8530 25287 8533
rect 23473 8528 25287 8530
rect 23473 8472 23478 8528
rect 23534 8472 25226 8528
rect 25282 8472 25287 8528
rect 23473 8470 25287 8472
rect 23473 8467 23539 8470
rect 25221 8467 25287 8470
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 24209 7986 24275 7989
rect 25221 7986 25287 7989
rect 24209 7984 25287 7986
rect 24209 7928 24214 7984
rect 24270 7928 25226 7984
rect 25282 7928 25287 7984
rect 24209 7926 25287 7928
rect 24209 7923 24275 7926
rect 25221 7923 25287 7926
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 38377 7578 38443 7581
rect 39200 7578 40000 7608
rect 38377 7576 40000 7578
rect 38377 7520 38382 7576
rect 38438 7520 40000 7576
rect 38377 7518 40000 7520
rect 38377 7515 38443 7518
rect 39200 7488 40000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 0 6808 858 6898
rect 798 6765 858 6808
rect 798 6760 907 6765
rect 798 6704 846 6760
rect 902 6704 907 6760
rect 798 6702 907 6704
rect 841 6699 907 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 0 6128 800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5538 800 5568
rect 0 5448 858 5538
rect 798 5405 858 5448
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 798 5400 907 5405
rect 798 5344 846 5400
rect 902 5344 907 5400
rect 798 5342 907 5344
rect 841 5339 907 5342
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 0 4768 800 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 0 4088 800 4118
rect 27153 4042 27219 4045
rect 29085 4042 29151 4045
rect 27153 4040 29151 4042
rect 27153 3984 27158 4040
rect 27214 3984 29090 4040
rect 29146 3984 29151 4040
rect 27153 3982 29151 3984
rect 27153 3979 27219 3982
rect 29085 3979 29151 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 24117 3634 24183 3637
rect 24761 3634 24827 3637
rect 26417 3634 26483 3637
rect 24117 3632 26483 3634
rect 24117 3576 24122 3632
rect 24178 3576 24766 3632
rect 24822 3576 26422 3632
rect 26478 3576 26483 3632
rect 24117 3574 26483 3576
rect 24117 3571 24183 3574
rect 24761 3571 24827 3574
rect 26417 3571 26483 3574
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 38469 3498 38535 3501
rect 39200 3498 40000 3528
rect 38469 3496 40000 3498
rect 38469 3440 38474 3496
rect 38530 3440 40000 3496
rect 38469 3438 40000 3440
rect 0 3408 800 3438
rect 38469 3435 38535 3438
rect 39200 3408 40000 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 24301 3090 24367 3093
rect 26233 3090 26299 3093
rect 24301 3088 26299 3090
rect 24301 3032 24306 3088
rect 24362 3032 26238 3088
rect 26294 3032 26299 3088
rect 24301 3030 26299 3032
rect 24301 3027 24367 3030
rect 26233 3027 26299 3030
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 38469 2818 38535 2821
rect 39200 2818 40000 2848
rect 38469 2816 40000 2818
rect 38469 2760 38474 2816
rect 38530 2760 40000 2816
rect 38469 2758 40000 2760
rect 0 2728 800 2758
rect 38469 2755 38535 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 40000 2758
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 38469 2138 38535 2141
rect 39200 2138 40000 2168
rect 38469 2136 40000 2138
rect 38469 2080 38474 2136
rect 38530 2080 40000 2136
rect 38469 2078 40000 2080
rect 38469 2075 38535 2078
rect 39200 2048 40000 2078
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 36124 20844 36188 20908
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 17908 19348 17972 19412
rect 36124 19348 36188 19412
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19380 16356 19444 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 17908 16220 17972 16284
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 19380 11460 19444 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 17907 19412 17973 19413
rect 17907 19348 17908 19412
rect 17972 19348 17973 19412
rect 17907 19347 17973 19348
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 17910 16285 17970 19347
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 19379 16420 19445 16421
rect 19379 16356 19380 16420
rect 19444 16356 19445 16420
rect 19379 16355 19445 16356
rect 17907 16284 17973 16285
rect 17907 16220 17908 16284
rect 17972 16220 17973 16284
rect 17907 16219 17973 16220
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 19382 11525 19442 16355
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 19379 11524 19445 11525
rect 19379 11460 19380 11524
rect 19444 11460 19445 11524
rect 19379 11459 19445 11460
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 36123 20908 36189 20909
rect 36123 20844 36124 20908
rect 36188 20844 36189 20908
rect 36123 20843 36189 20844
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 36126 19413 36186 20843
rect 36123 19412 36189 19413
rect 36123 19348 36124 19412
rect 36188 19348 36189 19412
rect 36123 19347 36189 19348
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__inv_2  _1278_
timestamp 18001
transform -1 0 15272 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 18001
transform -1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 18001
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1281_
timestamp 18001
transform -1 0 30820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 18001
transform -1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1283_
timestamp 18001
transform -1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 18001
transform -1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 18001
transform -1 0 7452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 18001
transform -1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 18001
transform -1 0 3036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 18001
transform 1 0 33028 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 18001
transform 1 0 28520 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 18001
transform -1 0 25484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 18001
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1292_
timestamp 18001
transform -1 0 27232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 18001
transform 1 0 26312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 18001
transform 1 0 36616 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1295_
timestamp 18001
transform 1 0 29992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1296_
timestamp 18001
transform 1 0 25944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 18001
transform 1 0 25024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 18001
transform 1 0 22632 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1299_
timestamp 18001
transform 1 0 22448 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 18001
transform 1 0 23552 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 18001
transform -1 0 25024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 18001
transform -1 0 16560 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 18001
transform 1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 18001
transform 1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1305_
timestamp 18001
transform -1 0 14996 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1306_
timestamp 18001
transform -1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1307_
timestamp 18001
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1308_
timestamp 18001
transform 1 0 13156 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1309_
timestamp 18001
transform 1 0 14904 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1310_
timestamp 18001
transform -1 0 18032 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1311_
timestamp 18001
transform 1 0 17020 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1312_
timestamp 18001
transform -1 0 17756 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1313_
timestamp 18001
transform 1 0 14812 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1314_
timestamp 18001
transform 1 0 17940 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 18001
transform 1 0 18768 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1316_
timestamp 18001
transform -1 0 21712 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1317_
timestamp 18001
transform 1 0 19688 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1318_
timestamp 18001
transform 1 0 19780 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1319_
timestamp 18001
transform -1 0 19136 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1320_
timestamp 18001
transform -1 0 18032 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1321_
timestamp 18001
transform -1 0 18492 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1322_
timestamp 18001
transform 1 0 18952 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1323_
timestamp 18001
transform -1 0 17020 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1324_
timestamp 18001
transform 1 0 7452 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1325_
timestamp 18001
transform -1 0 8372 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1326_
timestamp 18001
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 18001
transform 1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1328_
timestamp 18001
transform 1 0 7728 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1329_
timestamp 18001
transform -1 0 10120 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1330_
timestamp 18001
transform 1 0 4508 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_1  _1331_
timestamp 18001
transform 1 0 6716 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1332_
timestamp 18001
transform -1 0 7084 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1333_
timestamp 18001
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1334_
timestamp 18001
transform 1 0 7360 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _1335_
timestamp 18001
transform 1 0 8188 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1336_
timestamp 18001
transform -1 0 10396 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1337_
timestamp 18001
transform 1 0 8372 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1338_
timestamp 18001
transform -1 0 10488 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 18001
transform -1 0 11316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1340_
timestamp 18001
transform 1 0 10396 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1341_
timestamp 18001
transform -1 0 12236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1342_
timestamp 18001
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_1  _1343_
timestamp 18001
transform 1 0 8924 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1344_
timestamp 18001
transform 1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1345_
timestamp 18001
transform 1 0 4692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 18001
transform 1 0 9568 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1347_
timestamp 18001
transform 1 0 10580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1348_
timestamp 18001
transform 1 0 3772 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1349_
timestamp 18001
transform 1 0 4600 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1350_
timestamp 18001
transform -1 0 5060 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1351_
timestamp 18001
transform -1 0 4416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1352_
timestamp 18001
transform 1 0 4416 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1353_
timestamp 18001
transform 1 0 4416 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1354_
timestamp 18001
transform 1 0 4784 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 18001
transform 1 0 5612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1356_
timestamp 18001
transform 1 0 1656 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1357_
timestamp 18001
transform -1 0 25944 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1358_
timestamp 18001
transform -1 0 23920 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1359_
timestamp 18001
transform 1 0 25944 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1360_
timestamp 18001
transform 1 0 26220 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1361_
timestamp 18001
transform -1 0 28336 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1362_
timestamp 18001
transform 1 0 28336 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1363_
timestamp 18001
transform 1 0 31280 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 18001
transform 1 0 28704 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1365_
timestamp 18001
transform -1 0 29992 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1366_
timestamp 18001
transform 1 0 28980 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1367_
timestamp 18001
transform -1 0 31556 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1368_
timestamp 18001
transform -1 0 29808 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 18001
transform -1 0 28336 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1370_
timestamp 18001
transform -1 0 26220 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1371_
timestamp 18001
transform -1 0 32476 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1372_
timestamp 18001
transform -1 0 31924 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1373_
timestamp 18001
transform 1 0 30636 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1374_
timestamp 18001
transform -1 0 31188 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1375_
timestamp 18001
transform 1 0 29992 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1376_
timestamp 18001
transform 1 0 30176 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1377_
timestamp 18001
transform -1 0 30820 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1378_
timestamp 18001
transform -1 0 30084 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1379_
timestamp 18001
transform 1 0 30452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1380_
timestamp 18001
transform 1 0 21620 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1381_
timestamp 18001
transform 1 0 22264 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1382_
timestamp 18001
transform -1 0 20424 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1383_
timestamp 18001
transform -1 0 20700 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1384_
timestamp 18001
transform -1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1385_
timestamp 18001
transform -1 0 23736 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1386_
timestamp 18001
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1387_
timestamp 18001
transform 1 0 21804 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1388_
timestamp 18001
transform 1 0 21804 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1389_
timestamp 18001
transform -1 0 23092 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1390_
timestamp 18001
transform -1 0 21160 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1391_
timestamp 18001
transform -1 0 21068 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1392_
timestamp 18001
transform -1 0 21344 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1393_
timestamp 18001
transform 1 0 19412 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1394_
timestamp 18001
transform 1 0 21344 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1395_
timestamp 18001
transform -1 0 20424 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1396_
timestamp 18001
transform 1 0 19412 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1397_
timestamp 18001
transform 1 0 12236 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1398_
timestamp 18001
transform -1 0 12880 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1399_
timestamp 18001
transform -1 0 11408 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1400_
timestamp 18001
transform 1 0 9568 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1401_
timestamp 18001
transform -1 0 11132 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1402_
timestamp 18001
transform 1 0 10672 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1403_
timestamp 18001
transform 1 0 5520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1404_
timestamp 18001
transform 1 0 6440 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1405_
timestamp 18001
transform 1 0 6624 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1406_
timestamp 18001
transform 1 0 4692 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1407_
timestamp 18001
transform 1 0 6716 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1408_
timestamp 18001
transform 1 0 10212 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1409_
timestamp 18001
transform 1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1410_
timestamp 18001
transform -1 0 12144 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 18001
transform -1 0 11408 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1412_
timestamp 18001
transform -1 0 13800 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1413_
timestamp 18001
transform 1 0 13064 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1414_
timestamp 18001
transform 1 0 15824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1415_
timestamp 18001
transform -1 0 15732 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1416_
timestamp 18001
transform -1 0 17296 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1417_
timestamp 18001
transform -1 0 16560 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1418_
timestamp 18001
transform 1 0 18492 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1419_
timestamp 18001
transform -1 0 18400 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1420_
timestamp 18001
transform -1 0 17204 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1421_
timestamp 18001
transform -1 0 16560 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 18001
transform 1 0 18216 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1423_
timestamp 18001
transform 1 0 17756 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1424_
timestamp 18001
transform 1 0 18216 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1425_
timestamp 18001
transform 1 0 18952 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1426_
timestamp 18001
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1427_
timestamp 18001
transform 1 0 18492 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1428_
timestamp 18001
transform 1 0 17296 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1429_
timestamp 18001
transform -1 0 18400 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1430_
timestamp 18001
transform 1 0 16652 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1431_
timestamp 18001
transform -1 0 15824 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1432_
timestamp 18001
transform -1 0 14352 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1433_
timestamp 18001
transform 1 0 14812 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1434_
timestamp 18001
transform 1 0 15732 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1435_
timestamp 18001
transform -1 0 15456 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1436_
timestamp 18001
transform 1 0 14444 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1437_
timestamp 18001
transform 1 0 16008 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1438_
timestamp 18001
transform 1 0 15548 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1439_
timestamp 18001
transform -1 0 16560 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1440_
timestamp 18001
transform -1 0 17664 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1441_
timestamp 18001
transform 1 0 16652 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1442_
timestamp 18001
transform -1 0 16008 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1443_
timestamp 18001
transform -1 0 13616 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1444_
timestamp 18001
transform 1 0 14168 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1445_
timestamp 18001
transform -1 0 13984 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1446_
timestamp 18001
transform 1 0 14168 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1447_
timestamp 18001
transform 1 0 30820 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1448_
timestamp 18001
transform 1 0 30912 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1449_
timestamp 18001
transform -1 0 32016 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1450_
timestamp 18001
transform -1 0 35604 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1451_
timestamp 18001
transform 1 0 35972 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1452_
timestamp 18001
transform 1 0 36432 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1453_
timestamp 18001
transform 1 0 37260 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1454_
timestamp 18001
transform 1 0 37168 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1455_
timestamp 18001
transform -1 0 36800 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1456_
timestamp 18001
transform 1 0 38180 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 18001
transform 1 0 35880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 18001
transform 1 0 37444 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1459_
timestamp 18001
transform 1 0 33580 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 18001
transform -1 0 38364 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1461_
timestamp 18001
transform -1 0 37996 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1462_
timestamp 18001
transform -1 0 37904 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1463_
timestamp 18001
transform -1 0 37720 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1464_
timestamp 18001
transform 1 0 36892 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1465_
timestamp 18001
transform -1 0 36984 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1466_
timestamp 18001
transform -1 0 36524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1467_
timestamp 18001
transform -1 0 36616 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1468_
timestamp 18001
transform -1 0 37168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1469_
timestamp 18001
transform 1 0 35972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1470_
timestamp 18001
transform -1 0 37996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1471_
timestamp 18001
transform 1 0 36524 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1472_
timestamp 18001
transform 1 0 36340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1473_
timestamp 18001
transform 1 0 36248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1474_
timestamp 18001
transform 1 0 35788 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1475_
timestamp 18001
transform 1 0 35512 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1476_
timestamp 18001
transform 1 0 37444 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1477_
timestamp 18001
transform -1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1478_
timestamp 18001
transform -1 0 37812 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1479_
timestamp 18001
transform 1 0 36340 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1480_
timestamp 18001
transform -1 0 36616 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1481_
timestamp 18001
transform -1 0 36340 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1482_
timestamp 18001
transform -1 0 37168 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1483_
timestamp 18001
transform 1 0 36064 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1484_
timestamp 18001
transform -1 0 36064 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1485_
timestamp 18001
transform -1 0 35972 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1486_
timestamp 18001
transform 1 0 35788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1487_
timestamp 18001
transform 1 0 36064 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1488_
timestamp 18001
transform 1 0 36616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1489_
timestamp 18001
transform 1 0 34040 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1490_
timestamp 18001
transform -1 0 34040 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1491_
timestamp 18001
transform 1 0 33304 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1492_
timestamp 18001
transform 1 0 33948 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 18001
transform 1 0 34684 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1494_
timestamp 18001
transform -1 0 34500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1495_
timestamp 18001
transform 1 0 35144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1496_
timestamp 18001
transform -1 0 35604 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1497_
timestamp 18001
transform -1 0 34592 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1498_
timestamp 18001
transform -1 0 35604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1499_
timestamp 18001
transform -1 0 35236 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 18001
transform 1 0 34868 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1501_
timestamp 18001
transform -1 0 35144 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1502_
timestamp 18001
transform -1 0 34684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1503_
timestamp 18001
transform -1 0 33948 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1504_
timestamp 18001
transform 1 0 33856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1505_
timestamp 18001
transform -1 0 33120 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1506_
timestamp 18001
transform 1 0 31372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1507_
timestamp 18001
transform 1 0 31648 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1508_
timestamp 18001
transform 1 0 32108 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 18001
transform -1 0 32476 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1510_
timestamp 18001
transform 1 0 31924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1511_
timestamp 18001
transform -1 0 33396 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1512_
timestamp 18001
transform -1 0 32752 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1513_
timestamp 18001
transform -1 0 33948 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1514_
timestamp 18001
transform -1 0 34408 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1515_
timestamp 18001
transform 1 0 34408 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1516_
timestamp 18001
transform -1 0 34040 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1517_
timestamp 18001
transform 1 0 32844 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1518_
timestamp 18001
transform -1 0 33396 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1519_
timestamp 18001
transform -1 0 30544 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 18001
transform 1 0 29992 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1521_
timestamp 18001
transform -1 0 30728 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1522_
timestamp 18001
transform -1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1523_
timestamp 18001
transform -1 0 32752 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1524_
timestamp 18001
transform -1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1525_
timestamp 18001
transform -1 0 32200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1526_
timestamp 18001
transform 1 0 32936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1527_
timestamp 18001
transform 1 0 32476 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1528_
timestamp 18001
transform -1 0 32844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1529_
timestamp 18001
transform -1 0 31924 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1530_
timestamp 18001
transform 1 0 31556 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1531_
timestamp 18001
transform 1 0 29532 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1532_
timestamp 18001
transform 1 0 28704 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1533_
timestamp 18001
transform -1 0 28704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1534_
timestamp 18001
transform 1 0 28612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1535_
timestamp 18001
transform -1 0 30268 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1536_
timestamp 18001
transform 1 0 29992 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1537_
timestamp 18001
transform 1 0 31464 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1538_
timestamp 18001
transform 1 0 31004 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 18001
transform 1 0 31740 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1540_
timestamp 18001
transform 1 0 30452 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1541_
timestamp 18001
transform 1 0 30176 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1542_
timestamp 18001
transform 1 0 28888 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1543_
timestamp 18001
transform 1 0 28704 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1544_
timestamp 18001
transform -1 0 29532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1545_
timestamp 18001
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1546_
timestamp 18001
transform -1 0 30176 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1547_
timestamp 18001
transform -1 0 28704 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1548_
timestamp 18001
transform 1 0 31372 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1549_
timestamp 18001
transform -1 0 32660 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1550_
timestamp 18001
transform -1 0 33672 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1551_
timestamp 18001
transform -1 0 34960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1552_
timestamp 18001
transform 1 0 35696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1553_
timestamp 18001
transform -1 0 37168 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 18001
transform 1 0 37260 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1555_
timestamp 18001
transform -1 0 37076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1556_
timestamp 18001
transform -1 0 37812 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1557_
timestamp 18001
transform -1 0 38180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1558_
timestamp 18001
transform 1 0 37812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 18001
transform -1 0 37904 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1560_
timestamp 18001
transform -1 0 35236 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1561_
timestamp 18001
transform -1 0 35972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1562_
timestamp 18001
transform -1 0 37720 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1563_
timestamp 18001
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1564_
timestamp 18001
transform 1 0 36800 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1565_
timestamp 18001
transform -1 0 37904 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1566_
timestamp 18001
transform 1 0 37904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1567_
timestamp 18001
transform -1 0 37260 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1568_
timestamp 18001
transform -1 0 36800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1569_
timestamp 18001
transform 1 0 35512 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1570_
timestamp 18001
transform 1 0 35236 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1571_
timestamp 18001
transform 1 0 34868 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1572_
timestamp 18001
transform 1 0 35144 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1573_
timestamp 18001
transform -1 0 36340 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1574_
timestamp 18001
transform 1 0 34132 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1575_
timestamp 18001
transform 1 0 34684 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1576_
timestamp 18001
transform 1 0 31740 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1577_
timestamp 18001
transform -1 0 32936 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1578_
timestamp 18001
transform 1 0 34132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1579_
timestamp 18001
transform 1 0 33580 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1580_
timestamp 18001
transform 1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1581_
timestamp 18001
transform -1 0 31740 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1582_
timestamp 18001
transform 1 0 33672 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1583_
timestamp 18001
transform -1 0 33672 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1584_
timestamp 18001
transform -1 0 33028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1585_
timestamp 18001
transform -1 0 32936 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1586_
timestamp 18001
transform 1 0 30544 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1587_
timestamp 18001
transform 1 0 30544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1588_
timestamp 18001
transform -1 0 32476 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1589_
timestamp 18001
transform -1 0 31280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1590_
timestamp 18001
transform -1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1591_
timestamp 18001
transform 1 0 28980 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1592_
timestamp 18001
transform -1 0 29624 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1593_
timestamp 18001
transform 1 0 27140 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1594_
timestamp 18001
transform 1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1595_
timestamp 18001
transform 1 0 27692 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1596_
timestamp 18001
transform 1 0 28152 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1597_
timestamp 18001
transform 1 0 28060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1598_
timestamp 18001
transform -1 0 28244 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1599_
timestamp 18001
transform -1 0 27508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1600_
timestamp 18001
transform 1 0 26956 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1601_
timestamp 18001
transform -1 0 26864 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1602_
timestamp 18001
transform -1 0 27416 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1603_
timestamp 18001
transform -1 0 28336 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1604_
timestamp 18001
transform -1 0 28244 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _1605_
timestamp 18001
transform -1 0 27600 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1606_
timestamp 18001
transform -1 0 28152 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1607_
timestamp 18001
transform -1 0 28520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1608_
timestamp 18001
transform -1 0 27784 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1609_
timestamp 18001
transform -1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1610_
timestamp 18001
transform -1 0 31188 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1611_
timestamp 18001
transform 1 0 31188 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1612_
timestamp 18001
transform 1 0 32108 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1613_
timestamp 18001
transform 1 0 32752 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1614_
timestamp 18001
transform -1 0 35788 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1615_
timestamp 18001
transform -1 0 36616 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1616_
timestamp 18001
transform -1 0 37076 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1617_
timestamp 18001
transform -1 0 38456 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1618_
timestamp 18001
transform 1 0 36708 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1619_
timestamp 18001
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1620_
timestamp 18001
transform 1 0 32752 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1621_
timestamp 18001
transform -1 0 33028 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1622_
timestamp 18001
transform 1 0 32200 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1623_
timestamp 18001
transform 1 0 37260 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1624_
timestamp 18001
transform -1 0 33764 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1625_
timestamp 18001
transform -1 0 33120 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1626_
timestamp 18001
transform 1 0 32476 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1627_
timestamp 18001
transform -1 0 32476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1628_
timestamp 18001
transform -1 0 25668 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1629_
timestamp 18001
transform -1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1630_
timestamp 18001
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1631_
timestamp 18001
transform -1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1632_
timestamp 18001
transform 1 0 25116 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1633_
timestamp 18001
transform -1 0 25208 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1634_
timestamp 18001
transform -1 0 27048 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1635_
timestamp 18001
transform 1 0 26956 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1636_
timestamp 18001
transform 1 0 25484 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1637_
timestamp 18001
transform -1 0 29992 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1638_
timestamp 18001
transform -1 0 27968 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1639_
timestamp 18001
transform 1 0 29072 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1640_
timestamp 18001
transform -1 0 28520 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1641_
timestamp 18001
transform -1 0 29072 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1642_
timestamp 18001
transform -1 0 28612 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1643_
timestamp 18001
transform -1 0 30912 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1644_
timestamp 18001
transform -1 0 29808 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1645_
timestamp 18001
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1646_
timestamp 18001
transform -1 0 29256 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1647_
timestamp 18001
transform 1 0 28520 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1648_
timestamp 18001
transform -1 0 30452 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1649_
timestamp 18001
transform -1 0 31372 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1650_
timestamp 18001
transform -1 0 30912 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1651_
timestamp 18001
transform -1 0 34316 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1652_
timestamp 18001
transform -1 0 33856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 18001
transform -1 0 34592 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1654_
timestamp 18001
transform 1 0 32752 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1655_
timestamp 18001
transform -1 0 33304 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1656_
timestamp 18001
transform -1 0 34592 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1657_
timestamp 18001
transform 1 0 33488 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1658_
timestamp 18001
transform 1 0 33948 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1659_
timestamp 18001
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1660_
timestamp 18001
transform -1 0 34592 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1661_
timestamp 18001
transform 1 0 35420 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1662_
timestamp 18001
transform -1 0 34224 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1663_
timestamp 18001
transform 1 0 34684 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1664_
timestamp 18001
transform -1 0 34316 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1665_
timestamp 18001
transform 1 0 34316 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1666_
timestamp 18001
transform -1 0 34592 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1667_
timestamp 18001
transform -1 0 34316 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1668_
timestamp 18001
transform 1 0 33580 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1669_
timestamp 18001
transform 1 0 32844 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1670_
timestamp 18001
transform -1 0 33856 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1671_
timestamp 18001
transform -1 0 32568 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1672_
timestamp 18001
transform 1 0 31004 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1673_
timestamp 18001
transform -1 0 30084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1674_
timestamp 18001
transform 1 0 30084 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1675_
timestamp 18001
transform 1 0 31188 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1676_
timestamp 18001
transform -1 0 26680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1677_
timestamp 18001
transform -1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1678_
timestamp 18001
transform 1 0 26496 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1679_
timestamp 18001
transform -1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1680_
timestamp 18001
transform 1 0 26404 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1681_
timestamp 18001
transform -1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1682_
timestamp 18001
transform -1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1683_
timestamp 18001
transform 1 0 31648 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1684_
timestamp 18001
transform -1 0 31188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1685_
timestamp 18001
transform -1 0 31464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1686_
timestamp 18001
transform -1 0 32384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1687_
timestamp 18001
transform 1 0 33028 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1688_
timestamp 18001
transform 1 0 32384 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1689_
timestamp 18001
transform 1 0 27232 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1690_
timestamp 18001
transform -1 0 27140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1691_
timestamp 18001
transform 1 0 27784 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1692_
timestamp 18001
transform 1 0 27876 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1693_
timestamp 18001
transform 1 0 28520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1694_
timestamp 18001
transform -1 0 29624 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1695_
timestamp 18001
transform 1 0 28612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1696_
timestamp 18001
transform 1 0 28336 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1697_
timestamp 18001
transform -1 0 29900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1698_
timestamp 18001
transform -1 0 30176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1699_
timestamp 18001
transform 1 0 30728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1700_
timestamp 18001
transform 1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1701_
timestamp 18001
transform 1 0 31556 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1702_
timestamp 18001
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1703_
timestamp 18001
transform 1 0 32476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1704_
timestamp 18001
transform 1 0 29164 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1705_
timestamp 18001
transform 1 0 29716 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1706_
timestamp 18001
transform 1 0 28796 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1707_
timestamp 18001
transform -1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1708_
timestamp 18001
transform 1 0 27232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1709_
timestamp 18001
transform -1 0 27232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1710_
timestamp 18001
transform -1 0 27784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1711_
timestamp 18001
transform -1 0 28152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1712_
timestamp 18001
transform 1 0 28244 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1713_
timestamp 18001
transform -1 0 29348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1714_
timestamp 18001
transform -1 0 29624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1715_
timestamp 18001
transform 1 0 30452 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1716_
timestamp 18001
transform 1 0 30636 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1717_
timestamp 18001
transform 1 0 31556 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1718_
timestamp 18001
transform -1 0 32384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1719_
timestamp 18001
transform -1 0 32108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1720_
timestamp 18001
transform 1 0 29532 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1721_
timestamp 18001
transform 1 0 29992 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1722_
timestamp 18001
transform 1 0 27324 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1723_
timestamp 18001
transform -1 0 27692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1724_
timestamp 18001
transform -1 0 27416 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1725_
timestamp 18001
transform 1 0 26772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1726_
timestamp 18001
transform -1 0 27600 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1727_
timestamp 18001
transform 1 0 27600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1728_
timestamp 18001
transform -1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1729_
timestamp 18001
transform -1 0 28980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1730_
timestamp 18001
transform 1 0 30176 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1731_
timestamp 18001
transform 1 0 30912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1732_
timestamp 18001
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1733_
timestamp 18001
transform 1 0 30636 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1734_
timestamp 18001
transform 1 0 29532 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1735_
timestamp 18001
transform 1 0 26956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1736_
timestamp 18001
transform -1 0 25668 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1737_
timestamp 18001
transform -1 0 25944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1738_
timestamp 18001
transform 1 0 26220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1739_
timestamp 18001
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1740_
timestamp 18001
transform 1 0 27784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1741_
timestamp 18001
transform 1 0 28336 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1742_
timestamp 18001
transform 1 0 28796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1743_
timestamp 18001
transform 1 0 29992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1744_
timestamp 18001
transform 1 0 29624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1745_
timestamp 18001
transform 1 0 30544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1746_
timestamp 18001
transform -1 0 28520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1747_
timestamp 18001
transform -1 0 28336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1748_
timestamp 18001
transform 1 0 25852 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1749_
timestamp 18001
transform 1 0 22356 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1750_
timestamp 18001
transform 1 0 23368 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1751_
timestamp 18001
transform -1 0 26036 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1752_
timestamp 18001
transform -1 0 26864 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1753_
timestamp 18001
transform 1 0 27600 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp 18001
transform 1 0 28244 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1755_
timestamp 18001
transform 1 0 28704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1756_
timestamp 18001
transform 1 0 28796 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1757_
timestamp 18001
transform 1 0 25944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1758_
timestamp 18001
transform 1 0 27600 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1759_
timestamp 18001
transform 1 0 29256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1760_
timestamp 18001
transform 1 0 29256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1761_
timestamp 18001
transform 1 0 29532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1762_
timestamp 18001
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1763_
timestamp 18001
transform 1 0 29532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1764_
timestamp 18001
transform 1 0 31372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1765_
timestamp 18001
transform 1 0 31096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1766_
timestamp 18001
transform -1 0 32016 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1767_
timestamp 18001
transform 1 0 32108 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1768_
timestamp 18001
transform -1 0 32936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1769_
timestamp 18001
transform -1 0 33948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1770_
timestamp 18001
transform -1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1771_
timestamp 18001
transform -1 0 31280 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1772_
timestamp 18001
transform -1 0 34132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1773_
timestamp 18001
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1774_
timestamp 18001
transform -1 0 35420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1775_
timestamp 18001
transform 1 0 31556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1776_
timestamp 18001
transform -1 0 33028 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1777_
timestamp 18001
transform -1 0 34132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1778_
timestamp 18001
transform -1 0 34592 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1779_
timestamp 18001
transform -1 0 35328 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1780_
timestamp 18001
transform 1 0 35420 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1781_
timestamp 18001
transform 1 0 35144 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1782_
timestamp 18001
transform -1 0 35880 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1783_
timestamp 18001
transform -1 0 35512 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1784_
timestamp 18001
transform -1 0 35328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1785_
timestamp 18001
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1786_
timestamp 18001
transform 1 0 34224 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1787_
timestamp 18001
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1788_
timestamp 18001
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1789_
timestamp 18001
transform -1 0 34500 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1790_
timestamp 18001
transform 1 0 33120 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1791_
timestamp 18001
transform 1 0 33764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1792_
timestamp 18001
transform 1 0 32476 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1793_
timestamp 18001
transform 1 0 32936 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1794_
timestamp 18001
transform 1 0 33856 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1795_
timestamp 18001
transform -1 0 34960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1796_
timestamp 18001
transform 1 0 32108 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1797_
timestamp 18001
transform 1 0 33028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1798_
timestamp 18001
transform 1 0 32844 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1799_
timestamp 18001
transform -1 0 33028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1800_
timestamp 18001
transform -1 0 32936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1801_
timestamp 18001
transform 1 0 31464 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1802_
timestamp 18001
transform -1 0 31924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1803_
timestamp 18001
transform 1 0 32200 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1804_
timestamp 18001
transform 1 0 30912 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1805_
timestamp 18001
transform 1 0 30636 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1806_
timestamp 18001
transform -1 0 32384 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1807_
timestamp 18001
transform 1 0 29992 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1808_
timestamp 18001
transform 1 0 30728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1809_
timestamp 18001
transform 1 0 30636 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1810_
timestamp 18001
transform -1 0 30636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1811_
timestamp 18001
transform 1 0 28980 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1812_
timestamp 18001
transform 1 0 30452 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1813_
timestamp 18001
transform -1 0 23000 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1814_
timestamp 18001
transform 1 0 23920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1815_
timestamp 18001
transform 1 0 25944 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1816_
timestamp 18001
transform 1 0 25944 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1817_
timestamp 18001
transform -1 0 27508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1818_
timestamp 18001
transform 1 0 26956 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1819_
timestamp 18001
transform 1 0 27600 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _1820_
timestamp 18001
transform 1 0 28336 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1821_
timestamp 18001
transform -1 0 30452 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1822_
timestamp 18001
transform 1 0 30452 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1823_
timestamp 18001
transform -1 0 31832 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1824_
timestamp 18001
transform 1 0 32108 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1825_
timestamp 18001
transform -1 0 33488 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1826_
timestamp 18001
transform 1 0 33120 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1827_
timestamp 18001
transform 1 0 33396 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1828_
timestamp 18001
transform -1 0 35236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1829_
timestamp 18001
transform 1 0 34592 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1830_
timestamp 18001
transform -1 0 35972 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1831_
timestamp 18001
transform -1 0 35696 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1832_
timestamp 18001
transform -1 0 36432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1833_
timestamp 18001
transform 1 0 35512 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1834_
timestamp 18001
transform -1 0 34960 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1835_
timestamp 18001
transform -1 0 36984 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1836_
timestamp 18001
transform 1 0 35052 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1837_
timestamp 18001
transform -1 0 35052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1838_
timestamp 18001
transform 1 0 35144 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_1  _1839_
timestamp 18001
transform -1 0 36524 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1840_
timestamp 18001
transform -1 0 36892 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1841_
timestamp 18001
transform -1 0 28244 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1842_
timestamp 18001
transform -1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1843_
timestamp 18001
transform -1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1844_
timestamp 18001
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1845_
timestamp 18001
transform -1 0 26864 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1846_
timestamp 18001
transform 1 0 26588 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1847_
timestamp 18001
transform 1 0 28796 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1848_
timestamp 18001
transform 1 0 28152 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1849_
timestamp 18001
transform -1 0 28796 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1850_
timestamp 18001
transform -1 0 30268 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1851_
timestamp 18001
transform -1 0 30636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1852_
timestamp 18001
transform -1 0 29440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1853_
timestamp 18001
transform 1 0 30360 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1854_
timestamp 18001
transform -1 0 31096 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1855_
timestamp 18001
transform 1 0 30636 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1856_
timestamp 18001
transform 1 0 31096 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1857_
timestamp 18001
transform -1 0 31648 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1858_
timestamp 18001
transform 1 0 31096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1859_
timestamp 18001
transform -1 0 33580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1860_
timestamp 18001
transform -1 0 33212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1861_
timestamp 18001
transform -1 0 33304 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1862_
timestamp 18001
transform 1 0 32292 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1863_
timestamp 18001
transform 1 0 32660 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1864_
timestamp 18001
transform -1 0 36800 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1865_
timestamp 18001
transform 1 0 35512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1866_
timestamp 18001
transform 1 0 36616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1867_
timestamp 18001
transform 1 0 36800 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1868_
timestamp 18001
transform 1 0 37352 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1869_
timestamp 18001
transform 1 0 34408 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1870_
timestamp 18001
transform 1 0 35880 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1871_
timestamp 18001
transform 1 0 33948 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1872_
timestamp 18001
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1873_
timestamp 18001
transform 1 0 37260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1874_
timestamp 18001
transform -1 0 36708 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1875_
timestamp 18001
transform -1 0 37168 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1876_
timestamp 18001
transform -1 0 37904 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1877_
timestamp 18001
transform -1 0 36892 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1878_
timestamp 18001
transform -1 0 37628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1879_
timestamp 18001
transform -1 0 37168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1880_
timestamp 18001
transform -1 0 37168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1881_
timestamp 18001
transform -1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1882_
timestamp 18001
transform 1 0 35696 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1883_
timestamp 18001
transform -1 0 36340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1884_
timestamp 18001
transform -1 0 35604 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1885_
timestamp 18001
transform 1 0 35052 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1886_
timestamp 18001
transform -1 0 11592 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1887_
timestamp 18001
transform -1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1888_
timestamp 18001
transform 1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1889_
timestamp 18001
transform 1 0 8464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1890_
timestamp 18001
transform -1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1891_
timestamp 18001
transform -1 0 7176 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1892_
timestamp 18001
transform -1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1893_
timestamp 18001
transform -1 0 7636 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1894_
timestamp 18001
transform 1 0 8096 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1895_
timestamp 18001
transform -1 0 8832 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1896_
timestamp 18001
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1897_
timestamp 18001
transform 1 0 10212 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1898_
timestamp 18001
transform -1 0 8924 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1899_
timestamp 18001
transform 1 0 9108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1900_
timestamp 18001
transform 1 0 6348 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1901_
timestamp 18001
transform 1 0 7176 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1902_
timestamp 18001
transform 1 0 8096 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1903_
timestamp 18001
transform 1 0 8648 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1904_
timestamp 18001
transform 1 0 9568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1905_
timestamp 18001
transform 1 0 10856 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1906_
timestamp 18001
transform -1 0 10856 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1907_
timestamp 18001
transform 1 0 9844 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1908_
timestamp 18001
transform -1 0 10948 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1909_
timestamp 18001
transform -1 0 9844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1910_
timestamp 18001
transform 1 0 9844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1911_
timestamp 18001
transform -1 0 7912 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1912_
timestamp 18001
transform 1 0 8648 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1913_
timestamp 18001
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1914_
timestamp 18001
transform -1 0 9384 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1915_
timestamp 18001
transform 1 0 7176 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1916_
timestamp 18001
transform -1 0 7176 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1917_
timestamp 18001
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1918_
timestamp 18001
transform -1 0 6164 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1919_
timestamp 18001
transform -1 0 6348 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1920_
timestamp 18001
transform 1 0 5612 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1921_
timestamp 18001
transform 1 0 5612 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1922_
timestamp 18001
transform 1 0 5612 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1923_
timestamp 18001
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1924_
timestamp 18001
transform -1 0 6256 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1925_
timestamp 18001
transform -1 0 5612 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1926_
timestamp 18001
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1927_
timestamp 18001
transform -1 0 7176 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1928_
timestamp 18001
transform 1 0 5612 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1929_
timestamp 18001
transform 1 0 4324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1930_
timestamp 18001
transform 1 0 4784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1931_
timestamp 18001
transform -1 0 4232 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1932_
timestamp 18001
transform 1 0 2944 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1933_
timestamp 18001
transform 1 0 3312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1934_
timestamp 18001
transform -1 0 3680 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1935_
timestamp 18001
transform 1 0 2116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1936_
timestamp 18001
transform -1 0 2392 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1937_
timestamp 18001
transform -1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1938_
timestamp 18001
transform -1 0 3680 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1939_
timestamp 18001
transform -1 0 3496 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1940_
timestamp 18001
transform -1 0 3036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1941_
timestamp 18001
transform -1 0 3496 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1942_
timestamp 18001
transform -1 0 4048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1943_
timestamp 18001
transform -1 0 2576 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1944_
timestamp 18001
transform -1 0 4784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1945_
timestamp 18001
transform 1 0 3220 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1946_
timestamp 18001
transform 1 0 4784 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1947_
timestamp 18001
transform 1 0 4048 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1948_
timestamp 18001
transform 1 0 3220 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1949_
timestamp 18001
transform -1 0 3220 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1950_
timestamp 18001
transform -1 0 5152 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1951_
timestamp 18001
transform -1 0 5428 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1952_
timestamp 18001
transform -1 0 5888 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1953_
timestamp 18001
transform -1 0 4048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1954_
timestamp 18001
transform 1 0 8004 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1955_
timestamp 18001
transform -1 0 7544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1956_
timestamp 18001
transform 1 0 7084 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1957_
timestamp 18001
transform -1 0 8004 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1958_
timestamp 18001
transform 1 0 7360 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1959_
timestamp 18001
transform -1 0 7544 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1960_
timestamp 18001
transform -1 0 7912 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1961_
timestamp 18001
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1962_
timestamp 18001
transform -1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1963_
timestamp 18001
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1964_
timestamp 18001
transform 1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1965_
timestamp 18001
transform -1 0 11316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1966_
timestamp 18001
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1967_
timestamp 18001
transform -1 0 10304 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1968_
timestamp 18001
transform 1 0 11316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1969_
timestamp 18001
transform 1 0 10672 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1970_
timestamp 18001
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1971_
timestamp 18001
transform -1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1972_
timestamp 18001
transform 1 0 11040 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1973_
timestamp 18001
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1974_
timestamp 18001
transform 1 0 9108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1975_
timestamp 18001
transform -1 0 10580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1976_
timestamp 18001
transform 1 0 9936 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1977_
timestamp 18001
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1978_
timestamp 18001
transform -1 0 13156 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1979_
timestamp 18001
transform -1 0 12696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1980_
timestamp 18001
transform 1 0 12604 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1981_
timestamp 18001
transform 1 0 11960 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1982_
timestamp 18001
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1983_
timestamp 18001
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1984_
timestamp 18001
transform -1 0 12328 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1985_
timestamp 18001
transform -1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1986_
timestamp 18001
transform 1 0 11316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1987_
timestamp 18001
transform -1 0 11224 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1988_
timestamp 18001
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1989_
timestamp 18001
transform -1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1990_
timestamp 18001
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1991_
timestamp 18001
transform 1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1992_
timestamp 18001
transform -1 0 8740 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1993_
timestamp 18001
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1994_
timestamp 18001
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1995_
timestamp 18001
transform -1 0 8464 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1996_
timestamp 18001
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1997_
timestamp 18001
transform 1 0 7176 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1998_
timestamp 18001
transform -1 0 8648 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1999_
timestamp 18001
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2000_
timestamp 18001
transform 1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2001_
timestamp 18001
transform 1 0 7544 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2002_
timestamp 18001
transform 1 0 6900 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2003_
timestamp 18001
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2004_
timestamp 18001
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2005_
timestamp 18001
transform 1 0 5612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2006_
timestamp 18001
transform 1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2007_
timestamp 18001
transform -1 0 6808 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2008_
timestamp 18001
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2009_
timestamp 18001
transform 1 0 3220 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2010_
timestamp 18001
transform -1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2011_
timestamp 18001
transform -1 0 4508 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2012_
timestamp 18001
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2013_
timestamp 18001
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2014_
timestamp 18001
transform 1 0 4784 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2015_
timestamp 18001
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2016_
timestamp 18001
transform -1 0 2944 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2017_
timestamp 18001
transform 1 0 5244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2018_
timestamp 18001
transform 1 0 3220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2019_
timestamp 18001
transform 1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2020_
timestamp 18001
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2021_
timestamp 18001
transform -1 0 4324 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2022_
timestamp 18001
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2023_
timestamp 18001
transform 1 0 4692 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2024_
timestamp 18001
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2025_
timestamp 18001
transform -1 0 5888 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2026_
timestamp 18001
transform -1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2027_
timestamp 18001
transform 1 0 7268 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2028_
timestamp 18001
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2029_
timestamp 18001
transform -1 0 8740 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2030_
timestamp 18001
transform -1 0 7728 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2031_
timestamp 18001
transform 1 0 7176 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2032_
timestamp 18001
transform 1 0 2300 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2033_
timestamp 18001
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2034_
timestamp 18001
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2035_
timestamp 18001
transform -1 0 6164 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2036_
timestamp 18001
transform 1 0 7084 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2037_
timestamp 18001
transform 1 0 5612 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2038_
timestamp 18001
transform -1 0 5244 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2039_
timestamp 18001
transform -1 0 5612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2040_
timestamp 18001
transform -1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2041_
timestamp 18001
transform 1 0 2208 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2042_
timestamp 18001
transform -1 0 4232 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2043_
timestamp 18001
transform -1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2044_
timestamp 18001
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2045_
timestamp 18001
transform -1 0 3312 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2046_
timestamp 18001
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2047_
timestamp 18001
transform 1 0 2208 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2048_
timestamp 18001
transform -1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _2049_
timestamp 18001
transform -1 0 2760 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2050_
timestamp 18001
transform -1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2051_
timestamp 18001
transform 1 0 3220 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _2052_
timestamp 18001
transform -1 0 3496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2053_
timestamp 18001
transform 1 0 5336 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2054_
timestamp 18001
transform -1 0 5060 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2055_
timestamp 18001
transform -1 0 5244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2056_
timestamp 18001
transform -1 0 6256 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2057_
timestamp 18001
transform -1 0 3772 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2058_
timestamp 18001
transform 1 0 2944 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2059_
timestamp 18001
transform 1 0 2392 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2060_
timestamp 18001
transform -1 0 2392 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2061_
timestamp 18001
transform -1 0 3680 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2062_
timestamp 18001
transform -1 0 3772 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2063_
timestamp 18001
transform 1 0 2852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2064_
timestamp 18001
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2065_
timestamp 18001
transform 1 0 4048 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2066_
timestamp 18001
transform -1 0 5796 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2067_
timestamp 18001
transform 1 0 4048 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2068_
timestamp 18001
transform -1 0 24196 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2069_
timestamp 18001
transform -1 0 24840 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2070_
timestamp 18001
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2071_
timestamp 18001
transform 1 0 5152 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _2072_
timestamp 18001
transform 1 0 4140 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2073_
timestamp 18001
transform 1 0 3220 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _2074_
timestamp 18001
transform 1 0 3864 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2075_
timestamp 18001
transform -1 0 22356 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2076_
timestamp 18001
transform 1 0 23276 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2077_
timestamp 18001
transform 1 0 22816 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2078_
timestamp 18001
transform -1 0 22816 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2079_
timestamp 18001
transform 1 0 21712 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2080_
timestamp 18001
transform 1 0 22172 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2081_
timestamp 18001
transform -1 0 22172 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2082_
timestamp 18001
transform -1 0 23276 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2083_
timestamp 18001
transform -1 0 24380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2084_
timestamp 18001
transform 1 0 22356 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2085_
timestamp 18001
transform 1 0 21528 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2086_
timestamp 18001
transform 1 0 22172 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2087_
timestamp 18001
transform 1 0 24104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2088_
timestamp 18001
transform -1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2089_
timestamp 18001
transform 1 0 23644 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2090_
timestamp 18001
transform -1 0 25576 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _2091_
timestamp 18001
transform -1 0 24104 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2092_
timestamp 18001
transform 1 0 22080 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2093_
timestamp 18001
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _2094_
timestamp 18001
transform 1 0 25208 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2095_
timestamp 18001
transform -1 0 24840 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2096_
timestamp 18001
transform -1 0 27784 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2097_
timestamp 18001
transform -1 0 27324 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2098_
timestamp 18001
transform -1 0 27508 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2099_
timestamp 18001
transform 1 0 24380 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2100_
timestamp 18001
transform 1 0 23828 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2101_
timestamp 18001
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2102_
timestamp 18001
transform 1 0 23736 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2103_
timestamp 18001
transform -1 0 24104 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2104_
timestamp 18001
transform 1 0 23276 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2105_
timestamp 18001
transform 1 0 24380 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2106_
timestamp 18001
transform 1 0 23828 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2107_
timestamp 18001
transform -1 0 25208 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2108_
timestamp 18001
transform 1 0 25024 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2109_
timestamp 18001
transform 1 0 26036 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2110_
timestamp 18001
transform 1 0 24380 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2111_
timestamp 18001
transform 1 0 25024 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2112_
timestamp 18001
transform 1 0 23368 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2113_
timestamp 18001
transform 1 0 25208 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2114_
timestamp 18001
transform 1 0 24380 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2115_
timestamp 18001
transform 1 0 25208 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2116_
timestamp 18001
transform 1 0 25576 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2117_
timestamp 18001
transform 1 0 23920 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2118_
timestamp 18001
transform 1 0 24932 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2119_
timestamp 18001
transform 1 0 22632 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2120_
timestamp 18001
transform -1 0 28520 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2121_
timestamp 18001
transform 1 0 28244 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _2122_
timestamp 18001
transform -1 0 25944 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2123_
timestamp 18001
transform -1 0 25392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2124_
timestamp 18001
transform 1 0 24748 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2125_
timestamp 18001
transform 1 0 24380 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2126_
timestamp 18001
transform 1 0 23460 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2127_
timestamp 18001
transform -1 0 25944 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2128_
timestamp 18001
transform 1 0 26220 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2129_
timestamp 18001
transform 1 0 27876 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2130_
timestamp 18001
transform -1 0 26772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2131_
timestamp 18001
transform 1 0 27140 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2132_
timestamp 18001
transform -1 0 27140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _2133_
timestamp 18001
transform 1 0 27416 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2134_
timestamp 18001
transform -1 0 28704 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2135_
timestamp 18001
transform -1 0 28244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2136_
timestamp 18001
transform 1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2137_
timestamp 18001
transform 1 0 27508 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2138_
timestamp 18001
transform -1 0 15640 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2139_
timestamp 18001
transform -1 0 16376 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2140_
timestamp 18001
transform 1 0 16008 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2141_
timestamp 18001
transform 1 0 13432 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _2142_
timestamp 18001
transform 1 0 13524 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2143_
timestamp 18001
transform 1 0 15272 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2144_
timestamp 18001
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2145_
timestamp 18001
transform -1 0 14352 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2146_
timestamp 18001
transform -1 0 13432 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2147_
timestamp 18001
transform 1 0 15088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2148_
timestamp 18001
transform 1 0 15456 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _2149_
timestamp 18001
transform 1 0 14260 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2150_
timestamp 18001
transform 1 0 15732 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2151_
timestamp 18001
transform 1 0 17296 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2152_
timestamp 18001
transform -1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2153_
timestamp 18001
transform 1 0 12328 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2154_
timestamp 18001
transform 1 0 14352 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2155_
timestamp 18001
transform 1 0 15640 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2156_
timestamp 18001
transform -1 0 15548 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2157_
timestamp 18001
transform -1 0 13800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2158_
timestamp 18001
transform 1 0 13800 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2159_
timestamp 18001
transform -1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2160_
timestamp 18001
transform -1 0 13892 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2161_
timestamp 18001
transform 1 0 13708 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2162_
timestamp 18001
transform 1 0 12788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2163_
timestamp 18001
transform -1 0 13708 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2164_
timestamp 18001
transform -1 0 15088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2165_
timestamp 18001
transform 1 0 12604 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2166_
timestamp 18001
transform 1 0 14076 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _2167_
timestamp 18001
transform -1 0 14444 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2168_
timestamp 18001
transform 1 0 18400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2169_
timestamp 18001
transform -1 0 19504 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2170_
timestamp 18001
transform 1 0 19412 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2171_
timestamp 18001
transform 1 0 15824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2172_
timestamp 18001
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2173_
timestamp 18001
transform -1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2174_
timestamp 18001
transform -1 0 16652 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2175_
timestamp 18001
transform -1 0 15640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2176_
timestamp 18001
transform -1 0 14720 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2177_
timestamp 18001
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2178_
timestamp 18001
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2179_
timestamp 18001
transform 1 0 17572 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2180_
timestamp 18001
transform 1 0 19504 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2181_
timestamp 18001
transform 1 0 20792 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2182_
timestamp 18001
transform 1 0 17296 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2183_
timestamp 18001
transform -1 0 16008 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _2184_
timestamp 18001
transform 1 0 17480 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2185_
timestamp 18001
transform -1 0 18492 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2186_
timestamp 18001
transform -1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2187_
timestamp 18001
transform 1 0 19872 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2188_
timestamp 18001
transform 1 0 19504 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2189_
timestamp 18001
transform 1 0 18032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2190_
timestamp 18001
transform -1 0 20608 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2191_
timestamp 18001
transform -1 0 21160 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2192_
timestamp 18001
transform 1 0 18124 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2193_
timestamp 18001
transform 1 0 17572 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2194_
timestamp 18001
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2195_
timestamp 18001
transform 1 0 18584 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2196_
timestamp 18001
transform -1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2197_
timestamp 18001
transform 1 0 18124 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2198_
timestamp 18001
transform 1 0 18584 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2199_
timestamp 18001
transform -1 0 19136 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2200_
timestamp 18001
transform 1 0 20884 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2201_
timestamp 18001
transform 1 0 18676 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2202_
timestamp 18001
transform -1 0 21160 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2203_
timestamp 18001
transform 1 0 20608 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2204_
timestamp 18001
transform -1 0 22264 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _2205_
timestamp 18001
transform -1 0 21988 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2206_
timestamp 18001
transform -1 0 19872 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2207_
timestamp 18001
transform 1 0 20148 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2208_
timestamp 18001
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2209_
timestamp 18001
transform -1 0 19136 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _2210_
timestamp 18001
transform -1 0 20608 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2211_
timestamp 18001
transform -1 0 19872 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2212_
timestamp 18001
transform -1 0 19136 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2213_
timestamp 18001
transform 1 0 18216 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2214_
timestamp 18001
transform 1 0 18032 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2215_
timestamp 18001
transform -1 0 20056 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2216_
timestamp 18001
transform 1 0 21344 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2217_
timestamp 18001
transform 1 0 18492 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _2218_
timestamp 18001
transform 1 0 19872 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2219_
timestamp 18001
transform -1 0 21528 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2220_
timestamp 18001
transform 1 0 21160 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2221_
timestamp 18001
transform 1 0 18860 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2222_
timestamp 18001
transform -1 0 20148 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2223_
timestamp 18001
transform 1 0 19228 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2224_
timestamp 18001
transform 1 0 21344 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2225_
timestamp 18001
transform -1 0 20056 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2226_
timestamp 18001
transform -1 0 21252 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2227_
timestamp 18001
transform -1 0 22264 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2228_
timestamp 18001
transform 1 0 21712 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2229_
timestamp 18001
transform -1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2230_
timestamp 18001
transform -1 0 22632 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2231_
timestamp 18001
transform 1 0 21804 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2232_
timestamp 18001
transform 1 0 21804 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2233_
timestamp 18001
transform -1 0 21712 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2234_
timestamp 18001
transform -1 0 21896 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2235_
timestamp 18001
transform 1 0 21804 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2236_
timestamp 18001
transform 1 0 21804 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2237_
timestamp 18001
transform -1 0 22908 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2238_
timestamp 18001
transform -1 0 20608 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2239_
timestamp 18001
transform 1 0 19412 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2240_
timestamp 18001
transform -1 0 19964 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2241_
timestamp 18001
transform -1 0 19688 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2242_
timestamp 18001
transform 1 0 20056 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2243_
timestamp 18001
transform 1 0 20332 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2244_
timestamp 18001
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _2245_
timestamp 18001
transform 1 0 22356 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _2246_
timestamp 18001
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2247_
timestamp 18001
transform -1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2248_
timestamp 18001
transform 1 0 21160 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2249_
timestamp 18001
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2250_
timestamp 18001
transform -1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2251_
timestamp 18001
transform 1 0 21252 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2252_
timestamp 18001
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2253_
timestamp 18001
transform -1 0 23092 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2254_
timestamp 18001
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2255_
timestamp 18001
transform -1 0 20976 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2256_
timestamp 18001
transform 1 0 20148 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2257_
timestamp 18001
transform -1 0 21436 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2258_
timestamp 18001
transform -1 0 22540 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2259_
timestamp 18001
transform 1 0 18768 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2260_
timestamp 18001
transform -1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2261_
timestamp 18001
transform -1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2262_
timestamp 18001
transform 1 0 20792 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2263_
timestamp 18001
transform 1 0 19320 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2264_
timestamp 18001
transform 1 0 21068 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2265_
timestamp 18001
transform 1 0 20332 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2266_
timestamp 18001
transform 1 0 19780 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2267_
timestamp 18001
transform 1 0 19688 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2268_
timestamp 18001
transform -1 0 20608 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2269_
timestamp 18001
transform 1 0 19228 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2270_
timestamp 18001
transform -1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2271_
timestamp 18001
transform 1 0 20332 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2272_
timestamp 18001
transform -1 0 20332 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2273_
timestamp 18001
transform -1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2274_
timestamp 18001
transform -1 0 20148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2275_
timestamp 18001
transform 1 0 19320 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2276_
timestamp 18001
transform 1 0 23644 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2277_
timestamp 18001
transform -1 0 24748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2278_
timestamp 18001
transform -1 0 25668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2279_
timestamp 18001
transform -1 0 24748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2280_
timestamp 18001
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2281_
timestamp 18001
transform -1 0 22448 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2282_
timestamp 18001
transform 1 0 23092 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2283_
timestamp 18001
transform 1 0 22540 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2284_
timestamp 18001
transform 1 0 21804 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2285_
timestamp 18001
transform -1 0 25484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2286_
timestamp 18001
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2287_
timestamp 18001
transform 1 0 23552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2288_
timestamp 18001
transform 1 0 23552 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2289_
timestamp 18001
transform -1 0 24932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2290_
timestamp 18001
transform 1 0 25024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2291_
timestamp 18001
transform 1 0 25760 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2292_
timestamp 18001
transform -1 0 26404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2293_
timestamp 18001
transform -1 0 26128 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2294_
timestamp 18001
transform -1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2295_
timestamp 18001
transform -1 0 24932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2296_
timestamp 18001
transform -1 0 25852 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2297_
timestamp 18001
transform -1 0 25944 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2298_
timestamp 18001
transform 1 0 23644 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2299_
timestamp 18001
transform 1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _2300_
timestamp 18001
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _2301_
timestamp 18001
transform 1 0 22724 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _2302_
timestamp 18001
transform 1 0 22908 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2303_
timestamp 18001
transform -1 0 24564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2304_
timestamp 18001
transform 1 0 24380 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2305_
timestamp 18001
transform 1 0 24656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2306_
timestamp 18001
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2307_
timestamp 18001
transform 1 0 25760 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2308_
timestamp 18001
transform 1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2309_
timestamp 18001
transform -1 0 25576 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2310_
timestamp 18001
transform 1 0 25760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2311_
timestamp 18001
transform 1 0 25116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2312_
timestamp 18001
transform -1 0 23644 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2313_
timestamp 18001
transform 1 0 22172 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2314_
timestamp 18001
transform -1 0 26496 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2315_
timestamp 18001
transform -1 0 25576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2316_
timestamp 18001
transform -1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2317_
timestamp 18001
transform 1 0 22908 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2318_
timestamp 18001
transform 1 0 25392 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2319_
timestamp 18001
transform 1 0 24564 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2320_
timestamp 18001
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2321_
timestamp 18001
transform -1 0 24380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2322_
timestamp 18001
transform 1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2323_
timestamp 18001
transform 1 0 21712 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2324_
timestamp 18001
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _2325_
timestamp 18001
transform 1 0 21804 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2326_
timestamp 18001
transform -1 0 22908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2327_
timestamp 18001
transform -1 0 24656 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2328_
timestamp 18001
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2329_
timestamp 18001
transform -1 0 24380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2330_
timestamp 18001
transform 1 0 25576 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _2331_
timestamp 18001
transform 1 0 24472 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2332_
timestamp 18001
transform -1 0 23092 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2333_
timestamp 18001
transform 1 0 26956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _2334_
timestamp 18001
transform 1 0 24748 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2335_
timestamp 18001
transform 1 0 23644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2336_
timestamp 18001
transform 1 0 21804 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2337_
timestamp 18001
transform 1 0 20700 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2338_
timestamp 18001
transform -1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2339_
timestamp 18001
transform 1 0 22816 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2340_
timestamp 18001
transform 1 0 22172 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2341_
timestamp 18001
transform 1 0 21528 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _2342_
timestamp 18001
transform 1 0 23000 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2343_
timestamp 18001
transform 1 0 22816 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2344_
timestamp 18001
transform -1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2345_
timestamp 18001
transform -1 0 22816 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2346_
timestamp 18001
transform 1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2347_
timestamp 18001
transform 1 0 23552 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2348_
timestamp 18001
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2349_
timestamp 18001
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2350_
timestamp 18001
transform 1 0 23920 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2351_
timestamp 18001
transform 1 0 22080 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2352_
timestamp 18001
transform 1 0 21160 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2353_
timestamp 18001
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2354_
timestamp 18001
transform -1 0 23644 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2355_
timestamp 18001
transform 1 0 22172 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2356_
timestamp 18001
transform 1 0 23920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2357_
timestamp 18001
transform 1 0 25024 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2358_
timestamp 18001
transform -1 0 24104 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2359_
timestamp 18001
transform 1 0 24380 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2360_
timestamp 18001
transform -1 0 9844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2361_
timestamp 18001
transform 1 0 9200 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2362_
timestamp 18001
transform -1 0 10672 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2363_
timestamp 18001
transform -1 0 11316 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2364_
timestamp 18001
transform -1 0 11684 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2365_
timestamp 18001
transform 1 0 11040 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2366_
timestamp 18001
transform -1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2367_
timestamp 18001
transform 1 0 11500 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2368_
timestamp 18001
transform 1 0 12420 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2369_
timestamp 18001
transform 1 0 10580 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2370_
timestamp 18001
transform -1 0 10488 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2371_
timestamp 18001
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2372_
timestamp 18001
transform 1 0 10120 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2373_
timestamp 18001
transform 1 0 8372 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2374_
timestamp 18001
transform 1 0 9660 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2375_
timestamp 18001
transform -1 0 7360 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2376_
timestamp 18001
transform -1 0 8004 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2377_
timestamp 18001
transform -1 0 7268 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2378_
timestamp 18001
transform -1 0 6900 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2379_
timestamp 18001
transform 1 0 7176 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2380_
timestamp 18001
transform 1 0 7084 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2381_
timestamp 18001
transform 1 0 7452 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2382_
timestamp 18001
transform 1 0 7084 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2383_
timestamp 18001
transform -1 0 6992 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2384_
timestamp 18001
transform 1 0 6256 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2385_
timestamp 18001
transform 1 0 4968 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2386_
timestamp 18001
transform -1 0 5612 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2387_
timestamp 18001
transform 1 0 4416 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2388_
timestamp 18001
transform 1 0 3864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2389_
timestamp 18001
transform -1 0 5336 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2390_
timestamp 18001
transform 1 0 3772 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2391_
timestamp 18001
transform -1 0 4968 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2392_
timestamp 18001
transform -1 0 3680 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2393_
timestamp 18001
transform -1 0 4600 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2394_
timestamp 18001
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2395_
timestamp 18001
transform -1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2396_
timestamp 18001
transform -1 0 3496 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2397_
timestamp 18001
transform -1 0 5888 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2398_
timestamp 18001
transform -1 0 5060 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2399_
timestamp 18001
transform -1 0 4324 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2400_
timestamp 18001
transform -1 0 5888 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2401_
timestamp 18001
transform 1 0 4416 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2402_
timestamp 18001
transform 1 0 5152 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2403_
timestamp 18001
transform 1 0 6624 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2404_
timestamp 18001
transform 1 0 7268 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2405_
timestamp 18001
transform -1 0 9016 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2406_
timestamp 18001
transform -1 0 8004 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2407_
timestamp 18001
transform 1 0 7452 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2408_
timestamp 18001
transform 1 0 12972 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2409_
timestamp 18001
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2410_
timestamp 18001
transform 1 0 15364 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2411_
timestamp 18001
transform 1 0 16652 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2412_
timestamp 18001
transform 1 0 17572 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2413_
timestamp 18001
transform 1 0 15732 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2414_
timestamp 18001
transform 1 0 23368 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _2415_
timestamp 18001
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2416_
timestamp 18001
transform -1 0 25668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2417_
timestamp 18001
transform 1 0 23828 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2418_
timestamp 18001
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _2419_
timestamp 18001
transform 1 0 22908 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2420_
timestamp 18001
transform 1 0 22172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2421_
timestamp 18001
transform 1 0 23276 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2422_
timestamp 18001
transform -1 0 24012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2423_
timestamp 18001
transform 1 0 24012 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _2424_
timestamp 18001
transform 1 0 24840 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _2425_
timestamp 18001
transform 1 0 24472 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _2426_
timestamp 18001
transform 1 0 24472 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2427_
timestamp 18001
transform -1 0 25760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2428_
timestamp 18001
transform 1 0 24932 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2429_
timestamp 18001
transform 1 0 25116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2430_
timestamp 18001
transform -1 0 24472 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2431_
timestamp 18001
transform 1 0 24472 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _2432_
timestamp 18001
transform -1 0 25392 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2433_
timestamp 18001
transform -1 0 26036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2434_
timestamp 18001
transform -1 0 27324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2435_
timestamp 18001
transform 1 0 26588 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _2436_
timestamp 18001
transform 1 0 25944 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2437_
timestamp 18001
transform -1 0 29256 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2438_
timestamp 18001
transform 1 0 28428 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2439_
timestamp 18001
transform 1 0 27600 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2440_
timestamp 18001
transform 1 0 27508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2441_
timestamp 18001
transform 1 0 28980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2442_
timestamp 18001
transform 1 0 29808 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2443_
timestamp 18001
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2444_
timestamp 18001
transform 1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2445_
timestamp 18001
transform -1 0 26036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2446_
timestamp 18001
transform -1 0 26588 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2447_
timestamp 18001
transform 1 0 26680 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2448_
timestamp 18001
transform 1 0 28704 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2449_
timestamp 18001
transform -1 0 27508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2450_
timestamp 18001
transform 1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2451_
timestamp 18001
transform -1 0 30268 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2452_
timestamp 18001
transform -1 0 29532 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _2453_
timestamp 18001
transform 1 0 32476 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2454_
timestamp 18001
transform 1 0 32016 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2455_
timestamp 18001
transform -1 0 33396 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2456_
timestamp 18001
transform -1 0 32660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2457_
timestamp 18001
transform 1 0 29808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2458_
timestamp 18001
transform -1 0 32936 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2459_
timestamp 18001
transform 1 0 31004 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2460_
timestamp 18001
transform -1 0 33856 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2461_
timestamp 18001
transform -1 0 31004 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2462_
timestamp 18001
transform -1 0 30268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2463_
timestamp 18001
transform 1 0 31556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2464_
timestamp 18001
transform -1 0 35144 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2465_
timestamp 18001
transform -1 0 34592 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2466_
timestamp 18001
transform 1 0 32384 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2467_
timestamp 18001
transform 1 0 33028 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2468_
timestamp 18001
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2469_
timestamp 18001
transform -1 0 31924 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2470_
timestamp 18001
transform 1 0 29532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2471_
timestamp 18001
transform 1 0 29900 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2472_
timestamp 18001
transform -1 0 26864 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2473_
timestamp 18001
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2474_
timestamp 18001
transform 1 0 27784 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2475_
timestamp 18001
transform -1 0 28612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2476_
timestamp 18001
transform 1 0 28796 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2477_
timestamp 18001
transform 1 0 29808 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2478_
timestamp 18001
transform -1 0 33764 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2479_
timestamp 18001
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2480_
timestamp 18001
transform -1 0 34592 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_4  _2481_
timestamp 18001
transform 1 0 33580 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__o211ai_4  _2482_
timestamp 18001
transform -1 0 33396 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2483_
timestamp 18001
transform 1 0 26312 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 18001
transform 1 0 24656 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2485_
timestamp 18001
transform -1 0 27876 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2486_
timestamp 18001
transform 1 0 26956 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2487_
timestamp 18001
transform 1 0 27508 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2488_
timestamp 18001
transform 1 0 31372 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2489_
timestamp 18001
transform 1 0 27968 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2490_
timestamp 18001
transform 1 0 29072 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2491_
timestamp 18001
transform -1 0 29440 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2492_
timestamp 18001
transform 1 0 27876 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _2493_
timestamp 18001
transform 1 0 28060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2494_
timestamp 18001
transform -1 0 31464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2495_
timestamp 18001
transform 1 0 29992 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _2496_
timestamp 18001
transform 1 0 30360 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2497_
timestamp 18001
transform 1 0 31832 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _2498_
timestamp 18001
transform 1 0 32660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2499_
timestamp 18001
transform -1 0 33580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2500_
timestamp 18001
transform -1 0 34592 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2501_
timestamp 18001
transform -1 0 35512 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2502_
timestamp 18001
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2503_
timestamp 18001
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 18001
transform 1 0 23000 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2505_
timestamp 18001
transform -1 0 27876 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2506_
timestamp 18001
transform 1 0 27048 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2507_
timestamp 18001
transform 1 0 12788 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2508_
timestamp 18001
transform 1 0 13800 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2509_
timestamp 18001
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2510_
timestamp 18001
transform 1 0 14168 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2511_
timestamp 18001
transform 1 0 14996 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2512_
timestamp 18001
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2513_
timestamp 18001
transform 1 0 14720 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2514_
timestamp 18001
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2515_
timestamp 18001
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2516_
timestamp 18001
transform -1 0 15548 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2517_
timestamp 18001
transform -1 0 11408 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2518_
timestamp 18001
transform 1 0 12696 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2519_
timestamp 18001
transform -1 0 13984 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2520_
timestamp 18001
transform 1 0 13156 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _2521_
timestamp 18001
transform 1 0 15824 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2522_
timestamp 18001
transform -1 0 17848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _2523_
timestamp 18001
transform -1 0 18308 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _2524_
timestamp 18001
transform -1 0 12880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _2525_
timestamp 18001
transform 1 0 13432 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2526_
timestamp 18001
transform 1 0 16836 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2527_
timestamp 18001
transform 1 0 15916 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2528_
timestamp 18001
transform 1 0 16836 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2529_
timestamp 18001
transform 1 0 19228 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2530_
timestamp 18001
transform -1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2531_
timestamp 18001
transform -1 0 17664 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2532_
timestamp 18001
transform 1 0 16284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2533_
timestamp 18001
transform -1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2534_
timestamp 18001
transform 1 0 18492 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2535_
timestamp 18001
transform 1 0 14812 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2536_
timestamp 18001
transform 1 0 15640 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2537_
timestamp 18001
transform -1 0 16928 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 18001
transform 1 0 17296 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2539_
timestamp 18001
transform 1 0 17940 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 18001
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2541_
timestamp 18001
transform 1 0 17388 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 18001
transform 1 0 17572 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2543_
timestamp 18001
transform -1 0 15456 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2544_
timestamp 18001
transform -1 0 13156 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2545_
timestamp 18001
transform 1 0 12328 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2546_
timestamp 18001
transform 1 0 11960 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2547_
timestamp 18001
transform 1 0 13156 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2548_
timestamp 18001
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2549_
timestamp 18001
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2550_
timestamp 18001
transform -1 0 15364 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2551_
timestamp 18001
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2552_
timestamp 18001
transform -1 0 11408 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2553_
timestamp 18001
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2554_
timestamp 18001
transform 1 0 9568 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2555_
timestamp 18001
transform 1 0 9936 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2556_
timestamp 18001
transform -1 0 10028 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2557_
timestamp 18001
transform 1 0 11868 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2558_
timestamp 18001
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2559_
timestamp 18001
transform -1 0 13984 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2560_
timestamp 18001
transform -1 0 12328 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2561_
timestamp 18001
transform 1 0 9936 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2562_
timestamp 18001
transform 1 0 10028 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2563_
timestamp 18001
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2564_
timestamp 18001
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2565_
timestamp 18001
transform -1 0 13984 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2566_
timestamp 18001
transform 1 0 15272 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 18001
transform 1 0 15456 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2568_
timestamp 18001
transform 1 0 16376 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2569_
timestamp 18001
transform -1 0 17664 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2570_
timestamp 18001
transform 1 0 14720 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2571_
timestamp 18001
transform 1 0 13156 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2572_
timestamp 18001
transform 1 0 11776 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2573_
timestamp 18001
transform 1 0 10580 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2574_
timestamp 18001
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2575_
timestamp 18001
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2576_
timestamp 18001
transform -1 0 16468 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2577_
timestamp 18001
transform 1 0 14996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2578_
timestamp 18001
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2579_
timestamp 18001
transform 1 0 13340 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2580_
timestamp 18001
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2581_
timestamp 18001
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2582_
timestamp 18001
transform 1 0 12420 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2583_
timestamp 18001
transform -1 0 12420 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2584_
timestamp 18001
transform -1 0 13340 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2585_
timestamp 18001
transform 1 0 12788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2586_
timestamp 18001
transform -1 0 13248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2587_
timestamp 18001
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2588_
timestamp 18001
transform -1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2589_
timestamp 18001
transform 1 0 12696 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2590_
timestamp 18001
transform -1 0 13432 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2591_
timestamp 18001
transform -1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2592_
timestamp 18001
transform 1 0 18400 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2593_
timestamp 18001
transform 1 0 19228 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2594_
timestamp 18001
transform 1 0 16560 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2595_
timestamp 18001
transform 1 0 15364 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _2596_
timestamp 18001
transform 1 0 14812 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2597_
timestamp 18001
transform 1 0 13340 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2598_
timestamp 18001
transform -1 0 13800 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2599_
timestamp 18001
transform 1 0 13340 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2600_
timestamp 18001
transform -1 0 13156 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2601_
timestamp 18001
transform -1 0 13800 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2602_
timestamp 18001
transform -1 0 14720 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2603_
timestamp 18001
transform 1 0 17940 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2604_
timestamp 18001
transform 1 0 18308 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _2605_
timestamp 18001
transform -1 0 17020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2606_
timestamp 18001
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2607_
timestamp 18001
transform 1 0 15088 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2608_
timestamp 18001
transform 1 0 14996 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2609_
timestamp 18001
transform -1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2610_
timestamp 18001
transform 1 0 17296 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2611_
timestamp 18001
transform 1 0 17388 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _2612_
timestamp 18001
transform 1 0 15732 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 18001
transform -1 0 19136 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2614_
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 18001
transform 1 0 19872 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2616_
timestamp 18001
transform 1 0 21896 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2617_
timestamp 18001
transform 1 0 20424 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2618_
timestamp 18001
transform 1 0 19872 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2619_
timestamp 18001
transform 1 0 19228 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2620_
timestamp 18001
transform 1 0 27600 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2621_
timestamp 18001
transform -1 0 31280 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2622_
timestamp 18001
transform -1 0 33764 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2623_
timestamp 18001
transform 1 0 30452 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2624_
timestamp 18001
transform -1 0 32660 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2625_
timestamp 18001
transform -1 0 31096 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2626_
timestamp 18001
transform 1 0 22172 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2627_
timestamp 18001
transform -1 0 26312 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2628_
timestamp 18001
transform 1 0 21804 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2629_
timestamp 18001
transform 1 0 22540 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2630_
timestamp 18001
transform 1 0 24104 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2631_
timestamp 18001
transform -1 0 25668 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2632_
timestamp 18001
transform 1 0 24196 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2633_
timestamp 18001
transform -1 0 27324 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2634_
timestamp 18001
transform -1 0 27692 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2635_
timestamp 18001
transform -1 0 27876 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2636_
timestamp 18001
transform -1 0 27876 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2637_
timestamp 18001
transform -1 0 26864 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2638_
timestamp 18001
transform -1 0 26220 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2639_
timestamp 18001
transform 1 0 24840 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2640_
timestamp 18001
transform -1 0 24932 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2641_
timestamp 18001
transform 1 0 22356 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2642_
timestamp 18001
transform 1 0 24840 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 18001
transform 1 0 27324 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2644_
timestamp 18001
transform -1 0 30084 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2645_
timestamp 18001
transform 1 0 27416 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2646_
timestamp 18001
transform 1 0 21068 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2647_
timestamp 18001
transform 1 0 21712 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2648_
timestamp 18001
transform 1 0 18860 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2649_
timestamp 18001
transform 1 0 22816 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2650_
timestamp 18001
transform 1 0 23000 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2651_
timestamp 18001
transform 1 0 22080 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2652_
timestamp 18001
transform 1 0 22540 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2653_
timestamp 18001
transform -1 0 21436 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2654_
timestamp 18001
transform 1 0 21160 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2655_
timestamp 18001
transform 1 0 17204 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2656_
timestamp 18001
transform -1 0 22356 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2657_
timestamp 18001
transform 1 0 19228 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2658_
timestamp 18001
transform -1 0 21896 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2659_
timestamp 18001
transform 1 0 19320 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 18001
transform 1 0 18584 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2661_
timestamp 18001
transform 1 0 22080 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2662_
timestamp 18001
transform 1 0 10764 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2663_
timestamp 18001
transform 1 0 11316 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2664_
timestamp 18001
transform 1 0 12144 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2665_
timestamp 18001
transform -1 0 15824 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2666_
timestamp 18001
transform 1 0 15916 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2667_
timestamp 18001
transform -1 0 19228 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2668_
timestamp 18001
transform -1 0 20516 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2669_
timestamp 18001
transform -1 0 21068 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2670_
timestamp 18001
transform 1 0 16652 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2671_
timestamp 18001
transform 1 0 14352 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2672_
timestamp 18001
transform 1 0 13064 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2673_
timestamp 18001
transform 1 0 15456 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2674_
timestamp 18001
transform -1 0 19136 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2675_
timestamp 18001
transform 1 0 12328 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2676_
timestamp 18001
transform 1 0 13064 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2677_
timestamp 18001
transform 1 0 24380 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2678_
timestamp 18001
transform 1 0 22908 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2679_
timestamp 18001
transform 1 0 24472 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2680_
timestamp 18001
transform 1 0 26128 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2681_
timestamp 18001
transform 1 0 28060 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2682_
timestamp 18001
transform 1 0 28612 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 18001
transform 1 0 27968 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 18001
transform 1 0 27968 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 18001
transform 1 0 30176 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 18001
transform -1 0 35512 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2687_
timestamp 18001
transform -1 0 34316 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 18001
transform 1 0 34684 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2689_
timestamp 18001
transform 1 0 34868 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2690_
timestamp 18001
transform 1 0 35328 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2691_
timestamp 18001
transform 1 0 34868 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 18001
transform 1 0 33212 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 18001
transform 1 0 31740 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 18001
transform 1 0 30360 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _2695__125
timestamp 18001
transform -1 0 30176 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 18001
transform 1 0 29624 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _2696__124
timestamp 18001
transform -1 0 30728 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 18001
transform 1 0 30084 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2697_
timestamp 18001
transform 1 0 26956 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2698_
timestamp 18001
transform 1 0 26864 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2699_
timestamp 18001
transform 1 0 26956 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 18001
transform -1 0 30636 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2701_
timestamp 18001
transform 1 0 29532 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 18001
transform 1 0 31464 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2703_
timestamp 18001
transform 1 0 30544 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2704_
timestamp 18001
transform 1 0 32476 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2705_
timestamp 18001
transform 1 0 32752 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2706_
timestamp 18001
transform 1 0 36616 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2707_
timestamp 18001
transform 1 0 36432 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2708_
timestamp 18001
transform 1 0 34684 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2709_
timestamp 18001
transform 1 0 36616 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2710_
timestamp 18001
transform 1 0 36616 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2711_
timestamp 18001
transform 1 0 36708 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2712_
timestamp 18001
transform 1 0 36708 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2713_
timestamp 18001
transform 1 0 34684 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2714_
timestamp 18001
transform 1 0 34776 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _2715__123
timestamp 18001
transform -1 0 33120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2715_
timestamp 18001
transform 1 0 32568 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _2716__122
timestamp 18001
transform 1 0 32568 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2716_
timestamp 18001
transform 1 0 32844 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2717_
timestamp 18001
transform 1 0 6532 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2718_
timestamp 18001
transform -1 0 8832 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2719_
timestamp 18001
transform -1 0 9476 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2720_
timestamp 18001
transform 1 0 6624 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2721_
timestamp 18001
transform 1 0 6348 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2722_
timestamp 18001
transform -1 0 9752 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2723_
timestamp 18001
transform -1 0 10580 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 18001
transform 1 0 8924 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 18001
transform 1 0 10212 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 18001
transform 1 0 10212 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2727_
timestamp 18001
transform 1 0 9384 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2728_
timestamp 18001
transform 1 0 7544 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2729_
timestamp 18001
transform 1 0 6440 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2730_
timestamp 18001
transform 1 0 4600 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2731_
timestamp 18001
transform 1 0 4416 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2732_
timestamp 18001
transform 1 0 5612 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2733_
timestamp 18001
transform 1 0 6716 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2734_
timestamp 18001
transform 1 0 3864 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2735_
timestamp 18001
transform 1 0 2024 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2736_
timestamp 18001
transform 1 0 1380 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2737_
timestamp 18001
transform 1 0 1380 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2738_
timestamp 18001
transform 1 0 3772 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2739_
timestamp 18001
transform -1 0 5336 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2740_
timestamp 18001
transform 1 0 1380 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2741_
timestamp 18001
transform 1 0 1840 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2742_
timestamp 18001
transform -1 0 4048 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2743_
timestamp 18001
transform 1 0 4416 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2744_
timestamp 18001
transform 1 0 4784 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2745_
timestamp 18001
transform 1 0 7544 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2746_
timestamp 18001
transform 1 0 6808 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2747_
timestamp 18001
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _2748_
timestamp 18001
transform 1 0 19412 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _2749_
timestamp 18001
transform 1 0 19596 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2750_
timestamp 18001
transform 1 0 19688 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2751_
timestamp 18001
transform 1 0 19780 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2752_
timestamp 18001
transform 1 0 21068 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2753_
timestamp 18001
transform 1 0 22172 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2754_
timestamp 18001
transform 1 0 24472 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2755_
timestamp 18001
transform 1 0 22264 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2756_
timestamp 18001
transform 1 0 6624 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2757_
timestamp 18001
transform 1 0 6164 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2758_
timestamp 18001
transform 1 0 7820 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2759_
timestamp 18001
transform 1 0 6532 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2760_
timestamp 18001
transform 1 0 9016 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2761_
timestamp 18001
transform 1 0 9108 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2762_
timestamp 18001
transform 1 0 9568 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2763_
timestamp 18001
transform 1 0 10488 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2764_
timestamp 18001
transform 1 0 12144 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2765_
timestamp 18001
transform -1 0 15916 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2766_
timestamp 18001
transform -1 0 13984 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2767_
timestamp 18001
transform 1 0 11500 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2768_
timestamp 18001
transform -1 0 11408 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2769_
timestamp 18001
transform -1 0 9568 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2770_
timestamp 18001
transform 1 0 6900 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2771_
timestamp 18001
transform 1 0 6164 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2772_
timestamp 18001
transform 1 0 8924 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2773_
timestamp 18001
transform 1 0 6532 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2774_
timestamp 18001
transform 1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2775_
timestamp 18001
transform 1 0 5336 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2776_
timestamp 18001
transform 1 0 3864 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2777_
timestamp 18001
transform 1 0 3220 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2778_
timestamp 18001
transform 1 0 1840 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2779_
timestamp 18001
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2780_
timestamp 18001
transform -1 0 5796 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2781_
timestamp 18001
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2782_
timestamp 18001
transform 1 0 4968 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2783_
timestamp 18001
transform 1 0 5060 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2784_
timestamp 18001
transform 1 0 7728 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2785_
timestamp 18001
transform 1 0 6348 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2786_
timestamp 18001
transform 1 0 8924 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2787_
timestamp 18001
transform 1 0 9292 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2788_
timestamp 18001
transform 1 0 11132 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2789_
timestamp 18001
transform 1 0 9844 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2790_
timestamp 18001
transform -1 0 13616 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2791_
timestamp 18001
transform 1 0 9568 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2792_
timestamp 18001
transform -1 0 11040 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2793_
timestamp 18001
transform -1 0 9568 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2794_
timestamp 18001
transform 1 0 5704 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2795_
timestamp 18001
transform -1 0 9384 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2796_
timestamp 18001
transform -1 0 9568 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2797_
timestamp 18001
transform 1 0 4968 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2798_
timestamp 18001
transform 1 0 3312 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2799_
timestamp 18001
transform 1 0 1840 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2800_
timestamp 18001
transform 1 0 3864 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2801_
timestamp 18001
transform 1 0 2208 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 18001
transform 1 0 2576 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2803_
timestamp 18001
transform 1 0 4324 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 18001
transform 1 0 4416 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2805_
timestamp 18001
transform 1 0 6808 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2806_
timestamp 18001
transform 1 0 6532 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2807_
timestamp 18001
transform -1 0 10212 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2808_
timestamp 18001
transform 1 0 19228 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2809_
timestamp 18001
transform 1 0 12052 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2810_
timestamp 18001
transform 1 0 11040 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2811_
timestamp 18001
transform -1 0 15824 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2812_
timestamp 18001
transform -1 0 17296 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2813_
timestamp 18001
transform 1 0 17020 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2814_
timestamp 18001
transform 1 0 15088 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2815_
timestamp 18001
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _2816_
timestamp 18001
transform 1 0 24380 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2817_
timestamp 18001
transform 1 0 29992 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2818_
timestamp 18001
transform 1 0 27232 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2819_
timestamp 18001
transform 1 0 30084 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2820_
timestamp 18001
transform 1 0 32752 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2821_
timestamp 18001
transform 1 0 34592 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2822_
timestamp 18001
transform 1 0 35420 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2823_
timestamp 18001
transform 1 0 24932 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2824_
timestamp 18001
transform 1 0 21252 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2825_
timestamp 18001
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2826_
timestamp 18001
transform 1 0 26956 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2827_
timestamp 18001
transform 1 0 16652 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2828_
timestamp 18001
transform 1 0 19504 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2829_
timestamp 18001
transform 1 0 19412 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2830_
timestamp 18001
transform 1 0 14076 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2831_
timestamp 18001
transform 1 0 14444 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2832_
timestamp 18001
transform 1 0 16652 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2833_
timestamp 18001
transform 1 0 16928 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2834_
timestamp 18001
transform 1 0 17572 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2835_
timestamp 18001
transform 1 0 17756 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2836_
timestamp 18001
transform 1 0 16652 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2837_
timestamp 18001
transform -1 0 17572 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2838_
timestamp 18001
transform -1 0 16008 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2839_
timestamp 18001
transform -1 0 13616 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2840_
timestamp 18001
transform 1 0 10488 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2841_
timestamp 18001
transform 1 0 11316 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2842_
timestamp 18001
transform 1 0 11592 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2843_
timestamp 18001
transform 1 0 12512 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2844_
timestamp 18001
transform 1 0 14076 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2845_
timestamp 18001
transform -1 0 15824 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2846_
timestamp 18001
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2847_
timestamp 18001
transform 1 0 10764 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2848_
timestamp 18001
transform 1 0 9200 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2849_
timestamp 18001
transform 1 0 8740 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2850_
timestamp 18001
transform 1 0 8096 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2851_
timestamp 18001
transform 1 0 9384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2852_
timestamp 18001
transform -1 0 11868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2853_
timestamp 18001
transform 1 0 12696 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2854_
timestamp 18001
transform 1 0 13616 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2855_
timestamp 18001
transform -1 0 12604 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2856_
timestamp 18001
transform 1 0 9476 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2857_
timestamp 18001
transform 1 0 9108 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2858_
timestamp 18001
transform 1 0 9016 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2859_
timestamp 18001
transform 1 0 10856 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2860_
timestamp 18001
transform 1 0 14076 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2861_
timestamp 18001
transform 1 0 14720 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2862_
timestamp 18001
transform 1 0 14720 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2863_
timestamp 18001
transform 1 0 15732 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2864_
timestamp 18001
transform -1 0 19044 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2865_
timestamp 18001
transform 1 0 14168 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2866_
timestamp 18001
transform 1 0 12144 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2867_
timestamp 18001
transform -1 0 12144 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2868_
timestamp 18001
transform 1 0 10396 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2869_
timestamp 18001
transform 1 0 19044 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2870_
timestamp 18001
transform 1 0 19228 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2871_
timestamp 18001
transform 1 0 17940 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2872_
timestamp 18001
transform 1 0 2484 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2873_
timestamp 18001
transform 1 0 3772 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2874_
timestamp 18001
transform -1 0 6256 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2875_
timestamp 18001
transform 1 0 5888 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2876_
timestamp 18001
transform 1 0 4324 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2877_
timestamp 18001
transform 1 0 2484 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2878_
timestamp 18001
transform 1 0 1748 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2879_
timestamp 18001
transform 1 0 1380 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2880_
timestamp 18001
transform 1 0 1380 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2881_
timestamp 18001
transform 1 0 3496 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2882_
timestamp 18001
transform -1 0 6992 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2883_
timestamp 18001
transform -1 0 6900 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2884_
timestamp 18001
transform 1 0 1472 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2885_
timestamp 18001
transform 1 0 1380 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2886_
timestamp 18001
transform 1 0 2208 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2887_
timestamp 18001
transform -1 0 5704 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2888_
timestamp 18001
transform -1 0 6348 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2889_
timestamp 18001
transform 1 0 6624 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2890_
timestamp 18001
transform 1 0 17020 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _2956_
timestamp 18001
transform 1 0 2392 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2957_
timestamp 18001
transform -1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2958_
timestamp 18001
transform -1 0 38180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2959_
timestamp 18001
transform -1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2960_
timestamp 18001
transform 1 0 24196 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2961_
timestamp 18001
transform -1 0 25760 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2962_
timestamp 18001
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__X
timestamp 18001
transform -1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2089__A1
timestamp 18001
transform 1 0 24288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2090__S
timestamp 18001
transform 1 0 25024 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2092__S
timestamp 18001
transform -1 0 22080 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2502__S
timestamp 18001
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2657__RESET_B
timestamp 18001
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2670__RESET_B
timestamp 18001
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2707__CLK
timestamp 18001
transform 1 0 36248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2812__RESET_B
timestamp 18001
transform 1 0 14996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2814__RESET_B
timestamp 18001
transform 1 0 14904 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2854__RESET_B
timestamp 18001
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2863__RESET_B
timestamp 18001
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2870__RESET_B
timestamp 18001
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2871__RESET_B
timestamp 18001
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2889__Q
timestamp 18001
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform -1 0 21712 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform 1 0 23644 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_A
timestamp 18001
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_X
timestamp 18001
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_A
timestamp 18001
transform 1 0 12420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_X
timestamp 18001
transform 1 0 12604 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_A
timestamp 18001
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_X
timestamp 18001
transform 1 0 31556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_A
timestamp 18001
transform 1 0 29808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_X
timestamp 18001
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_clk_A
timestamp 18001
transform 1 0 7360 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_clk_A
timestamp 18001
transform 1 0 5060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_clk_A
timestamp 18001
transform -1 0 11776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_clk_A
timestamp 18001
transform -1 0 14720 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_clk_A
timestamp 18001
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_clk_A
timestamp 18001
transform 1 0 5244 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_clk_A
timestamp 18001
transform 1 0 5336 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_clk_A
timestamp 18001
transform 1 0 7912 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_clk_A
timestamp 18001
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_clk_A
timestamp 18001
transform 1 0 11408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_clk_A
timestamp 18001
transform 1 0 18676 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_clk_A
timestamp 18001
transform 1 0 14168 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_clk_A
timestamp 18001
transform 1 0 22816 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_clk_A
timestamp 18001
transform 1 0 26404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_clk_A
timestamp 18001
transform 1 0 23736 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_clk_A
timestamp 18001
transform 1 0 30820 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_clk_A
timestamp 18001
transform 1 0 32936 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_clk_A
timestamp 18001
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_clk_A
timestamp 18001
transform 1 0 28244 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_clk_A
timestamp 18001
transform -1 0 27232 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_clk_A
timestamp 18001
transform 1 0 32384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_clk_A
timestamp 18001
transform 1 0 35604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_clk_A
timestamp 18001
transform 1 0 23920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_clk_A
timestamp 18001
transform 1 0 23644 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_clk_A
timestamp 18001
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_clk_A
timestamp 18001
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_clk_A
timestamp 18001
transform 1 0 17572 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_28_clk_A
timestamp 18001
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_29_clk_A
timestamp 18001
transform -1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 18001
transform 1 0 12512 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp 18001
transform 1 0 30084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload2_A
timestamp 18001
transform 1 0 30360 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout35_A
timestamp 18001
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout56_A
timestamp 18001
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout58_A
timestamp 18001
transform -1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout59_A
timestamp 18001
transform 1 0 11500 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout60_A
timestamp 18001
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout61_A
timestamp 18001
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout61_X
timestamp 18001
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout67_A
timestamp 18001
transform 1 0 4048 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout68_A
timestamp 18001
transform 1 0 12696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout69_A
timestamp 18001
transform 1 0 18400 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout70_A
timestamp 18001
transform 1 0 12880 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout71_A
timestamp 18001
transform -1 0 12144 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout71_X
timestamp 18001
transform 1 0 12512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout72_A
timestamp 18001
transform 1 0 4324 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout72_X
timestamp 18001
transform 1 0 4968 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_A
timestamp 18001
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout78_A
timestamp 18001
transform 1 0 29900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout79_A
timestamp 18001
transform 1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout80_A
timestamp 18001
transform 1 0 25852 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout83_A
timestamp 18001
transform 1 0 21344 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout86_A
timestamp 18001
transform -1 0 30728 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout87_A
timestamp 18001
transform -1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout87_X
timestamp 18001
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 1840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 14904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 1840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform 1 0 21804 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 18001
transform -1 0 12972 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 18001
transform -1 0 12420 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 18001
transform 1 0 29716 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 18001
transform 1 0 29992 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_0_clk
timestamp 18001
transform 1 0 6348 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_1_clk
timestamp 18001
transform -1 0 5060 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_2_clk
timestamp 18001
transform 1 0 9936 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_3_clk
timestamp 18001
transform 1 0 14720 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_4_clk
timestamp 18001
transform 1 0 9844 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_5_clk
timestamp 18001
transform -1 0 5244 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_6_clk
timestamp 18001
transform 1 0 4324 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_7_clk
timestamp 18001
transform 1 0 6348 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_8_clk
timestamp 18001
transform -1 0 5428 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_9_clk
timestamp 18001
transform 1 0 11592 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_10_clk
timestamp 18001
transform 1 0 18860 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_11_clk
timestamp 18001
transform 1 0 14352 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_12_clk
timestamp 18001
transform -1 0 22172 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_13_clk
timestamp 18001
transform 1 0 24932 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_14_clk
timestamp 18001
transform 1 0 22356 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_15_clk
timestamp 18001
transform 1 0 29532 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_16_clk
timestamp 18001
transform -1 0 34132 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_17_clk
timestamp 18001
transform 1 0 34592 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_18_clk
timestamp 18001
transform 1 0 26956 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_19_clk
timestamp 18001
transform 1 0 26036 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_20_clk
timestamp 18001
transform 1 0 33120 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_21_clk
timestamp 18001
transform 1 0 35788 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_23_clk
timestamp 18001
transform -1 0 23920 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_24_clk
timestamp 18001
transform -1 0 23644 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_25_clk
timestamp 18001
transform 1 0 19228 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_26_clk
timestamp 18001
transform 1 0 16376 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_27_clk
timestamp 18001
transform 1 0 17756 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_28_clk
timestamp 18001
transform 1 0 10396 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_29_clk
timestamp 18001
transform 1 0 4232 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 18001
transform 1 0 11500 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_6  clkload1
timestamp 18001
transform 1 0 29440 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload2
timestamp 18001
transform 1 0 28520 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload3
timestamp 18001
transform 1 0 3772 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  clkload4
timestamp 18001
transform 1 0 9936 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload5
timestamp 18001
transform 1 0 18492 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  clkload6
timestamp 18001
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_6  clkload7
timestamp 18001
transform 1 0 17756 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  clkload8
timestamp 18001
transform 1 0 10764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload9
timestamp 18001
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload10
timestamp 18001
transform 1 0 14352 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_6  clkload11
timestamp 18001
transform 1 0 9844 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload12
timestamp 18001
transform 1 0 5060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload13
timestamp 18001
transform 1 0 5336 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload14
timestamp 18001
transform 1 0 6348 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload15
timestamp 18001
transform 1 0 5428 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload16
timestamp 18001
transform 1 0 19228 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload17
timestamp 18001
transform 1 0 14904 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload18
timestamp 18001
transform 1 0 26036 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload19
timestamp 18001
transform 1 0 35788 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload20
timestamp 18001
transform -1 0 23460 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload21
timestamp 18001
transform 1 0 22632 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload22
timestamp 18001
transform 1 0 22172 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  clkload23
timestamp 18001
transform 1 0 22356 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  clkload24
timestamp 18001
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  clkload25
timestamp 18001
transform 1 0 33120 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload26
timestamp 18001
transform 1 0 34592 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload27
timestamp 18001
transform 1 0 26220 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 18001
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 18001
transform 1 0 12788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 18001
transform -1 0 10856 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 18001
transform 1 0 14996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 18001
transform -1 0 18492 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 18001
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 18001
transform 1 0 27140 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 18001
transform -1 0 31924 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout22
timestamp 18001
transform 1 0 33948 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 18001
transform 1 0 35604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 18001
transform 1 0 35144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 18001
transform -1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 18001
transform -1 0 15456 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 18001
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout33
timestamp 18001
transform -1 0 14260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 18001
transform 1 0 18400 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 18001
transform 1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout36
timestamp 18001
transform 1 0 36984 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 18001
transform 1 0 36616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 18001
transform -1 0 33764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 18001
transform -1 0 32016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout40
timestamp 18001
transform 1 0 34592 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 18001
transform -1 0 29808 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 18001
transform 1 0 25852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 18001
transform 1 0 15824 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 18001
transform -1 0 25852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 18001
transform 1 0 26956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 18001
transform -1 0 24472 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 18001
transform 1 0 23368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 18001
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 18001
transform 1 0 25300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 18001
transform -1 0 4324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 18001
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 18001
transform 1 0 3128 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 18001
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 18001
transform 1 0 8004 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 18001
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout56
timestamp 18001
transform -1 0 4416 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 18001
transform 1 0 12512 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 18001
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 18001
transform 1 0 11684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 18001
transform -1 0 18768 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 18001
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 18001
transform 1 0 4784 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 18001
transform -1 0 3680 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp 18001
transform -1 0 3680 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 18001
transform -1 0 9200 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 18001
transform -1 0 4140 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp 18001
transform 1 0 3680 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 18001
transform -1 0 12144 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 18001
transform 1 0 17388 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 18001
transform 1 0 12328 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 18001
transform 1 0 12144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 18001
transform -1 0 4692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout73
timestamp 18001
transform -1 0 21068 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 18001
transform 1 0 27508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 18001
transform -1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 18001
transform -1 0 35236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout77
timestamp 18001
transform 1 0 29532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 18001
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout79
timestamp 18001
transform -1 0 20792 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout80
timestamp 18001
transform -1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 18001
transform -1 0 20976 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout82
timestamp 18001
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout83
timestamp 18001
transform -1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout84
timestamp 18001
transform -1 0 30360 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout85
timestamp 18001
transform 1 0 29532 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout86
timestamp 18001
transform 1 0 29992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp 18001
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 18001
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 18001
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 18001
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 18001
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93
timestamp 1636986456
transform 1 0 9660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 18001
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 18001
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636986456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636986456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 18001
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_141
timestamp 18001
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 18001
transform 1 0 14628 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636986456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 18001
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636986456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636986456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 18001
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636986456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 18001
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_217
timestamp 18001
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636986456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_237
timestamp 18001
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_245
timestamp 18001
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 18001
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 18001
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_258
timestamp 1636986456
transform 1 0 24840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 18001
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 18001
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 18001
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 18001
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_293
timestamp 18001
transform 1 0 28060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_301
timestamp 18001
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 18001
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 18001
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 18001
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636986456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 18001
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636986456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636986456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 18001
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 18001
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 18001
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 18001
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 18001
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 18001
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_401
timestamp 18001
transform 1 0 37996 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6
timestamp 1636986456
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_18
timestamp 18001
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_22
timestamp 18001
transform 1 0 3128 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_50
timestamp 18001
transform 1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 18001
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp 18001
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_133
timestamp 1636986456
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1636986456
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 18001
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 18001
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 18001
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_249
timestamp 18001
transform 1 0 24012 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_253
timestamp 18001
transform 1 0 24380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 18001
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_284
timestamp 18001
transform 1 0 27232 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_290
timestamp 18001
transform 1 0 27784 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_298
timestamp 1636986456
transform 1 0 28520 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 18001
transform 1 0 29624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 18001
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_321
timestamp 18001
transform 1 0 30636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 18001
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 18001
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_401
timestamp 18001
transform 1 0 37996 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6
timestamp 1636986456
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 18001
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 18001
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_45
timestamp 18001
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_107
timestamp 18001
transform 1 0 10948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 18001
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 18001
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 18001
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 18001
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 18001
transform 1 0 27968 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 18001
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 18001
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_320
timestamp 18001
transform 1 0 30544 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_340
timestamp 1636986456
transform 1 0 32384 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_352
timestamp 1636986456
transform 1 0 33488 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_401
timestamp 18001
transform 1 0 37996 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 18001
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 18001
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_47
timestamp 18001
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 18001
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_63
timestamp 18001
transform 1 0 6900 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_74
timestamp 18001
transform 1 0 7912 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 18001
transform 1 0 8464 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_84
timestamp 1636986456
transform 1 0 8832 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 18001
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_103
timestamp 18001
transform 1 0 10580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 18001
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_116
timestamp 18001
transform 1 0 11776 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_122
timestamp 18001
transform 1 0 12328 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_126
timestamp 1636986456
transform 1 0 12696 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_138
timestamp 1636986456
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_150
timestamp 1636986456
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 18001
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_225
timestamp 18001
transform 1 0 21804 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_266
timestamp 18001
transform 1 0 25576 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_295
timestamp 18001
transform 1 0 28244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_301
timestamp 18001
transform 1 0 28796 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_313
timestamp 18001
transform 1 0 29900 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_321
timestamp 18001
transform 1 0 30636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 18001
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_337
timestamp 18001
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_353
timestamp 1636986456
transform 1 0 33580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_365
timestamp 1636986456
transform 1 0 34684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_377
timestamp 1636986456
transform 1 0 35788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp 18001
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 18001
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6
timestamp 1636986456
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 18001
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 18001
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 18001
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 18001
transform 1 0 6348 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 18001
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_94
timestamp 18001
transform 1 0 9752 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 18001
transform 1 0 10304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_110
timestamp 18001
transform 1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp 18001
transform 1 0 11960 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636986456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_220
timestamp 1636986456
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_236
timestamp 18001
transform 1 0 22816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_246
timestamp 18001
transform 1 0 23736 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp 18001
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_277
timestamp 18001
transform 1 0 26588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_283
timestamp 18001
transform 1 0 27140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 18001
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_295
timestamp 18001
transform 1 0 28244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 18001
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 18001
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_345
timestamp 18001
transform 1 0 32844 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_373
timestamp 1636986456
transform 1 0 35420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_385
timestamp 1636986456
transform 1 0 36524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_397
timestamp 18001
transform 1 0 37628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 18001
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6
timestamp 1636986456
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_18
timestamp 18001
transform 1 0 2760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_22
timestamp 18001
transform 1 0 3128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 18001
transform 1 0 6808 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_71
timestamp 1636986456
transform 1 0 7636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 18001
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 18001
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_135
timestamp 1636986456
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_147
timestamp 1636986456
transform 1 0 14628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_159
timestamp 18001
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 18001
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 18001
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_201
timestamp 18001
transform 1 0 19596 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_239
timestamp 1636986456
transform 1 0 23092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_251
timestamp 18001
transform 1 0 24196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 18001
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 18001
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636986456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 18001
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 18001
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_320
timestamp 18001
transform 1 0 30544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_328
timestamp 18001
transform 1 0 31280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_344
timestamp 18001
transform 1 0 32752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_357
timestamp 18001
transform 1 0 33948 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636986456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 18001
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 18001
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 18001
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 18001
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp 18001
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 18001
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_62
timestamp 18001
transform 1 0 6808 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 18001
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 18001
transform 1 0 11776 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_124
timestamp 18001
transform 1 0 12512 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_161
timestamp 1636986456
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_173
timestamp 1636986456
transform 1 0 17020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_185
timestamp 18001
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 18001
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636986456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 18001
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_217
timestamp 18001
transform 1 0 21068 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_227
timestamp 18001
transform 1 0 21988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 18001
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 18001
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp 18001
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_276
timestamp 18001
transform 1 0 26496 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636986456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 18001
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 18001
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 18001
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_316
timestamp 1636986456
transform 1 0 30176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_328
timestamp 18001
transform 1 0 31280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_337
timestamp 18001
transform 1 0 32108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_345
timestamp 18001
transform 1 0 32844 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_353
timestamp 18001
transform 1 0 33580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_358
timestamp 18001
transform 1 0 34040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_368
timestamp 18001
transform 1 0 34960 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_376
timestamp 1636986456
transform 1 0 35696 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_388
timestamp 1636986456
transform 1 0 36800 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_400
timestamp 18001
transform 1 0 37904 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 18001
transform 1 0 38456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6
timestamp 18001
transform 1 0 1656 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_12
timestamp 18001
transform 1 0 2208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_28
timestamp 18001
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 18001
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 18001
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 18001
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 18001
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_86
timestamp 18001
transform 1 0 9016 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 18001
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 18001
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 18001
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_134
timestamp 1636986456
transform 1 0 13432 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_146
timestamp 1636986456
transform 1 0 14536 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 18001
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 18001
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636986456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_188
timestamp 1636986456
transform 1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_200
timestamp 1636986456
transform 1 0 19504 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1636986456
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 18001
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_266
timestamp 18001
transform 1 0 25576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_273
timestamp 18001
transform 1 0 26220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 18001
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_294
timestamp 18001
transform 1 0 28152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_310
timestamp 18001
transform 1 0 29624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_318
timestamp 18001
transform 1 0 30360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_330
timestamp 18001
transform 1 0 31464 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_351
timestamp 1636986456
transform 1 0 33396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_363
timestamp 18001
transform 1 0 34500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_372
timestamp 18001
transform 1 0 35328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_381
timestamp 18001
transform 1 0 36156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_389
timestamp 18001
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636986456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 18001
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 18001
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 18001
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_117
timestamp 18001
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_149
timestamp 1636986456
transform 1 0 14812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_161
timestamp 1636986456
transform 1 0 15916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_173
timestamp 18001
transform 1 0 17020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 18001
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 18001
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 18001
transform 1 0 19596 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_222
timestamp 1636986456
transform 1 0 21528 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_237
timestamp 1636986456
transform 1 0 22908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 18001
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 18001
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_259
timestamp 18001
transform 1 0 24932 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_275
timestamp 18001
transform 1 0 26404 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_283
timestamp 18001
transform 1 0 27140 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_292
timestamp 1636986456
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 18001
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_319
timestamp 1636986456
transform 1 0 30452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_331
timestamp 18001
transform 1 0 31556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_342
timestamp 18001
transform 1 0 32568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_346
timestamp 18001
transform 1 0 32936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_350
timestamp 18001
transform 1 0 33304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 18001
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 18001
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_371
timestamp 18001
transform 1 0 35236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_378
timestamp 18001
transform 1 0 35880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_6
timestamp 18001
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_14
timestamp 18001
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 18001
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1636986456
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636986456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 18001
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_80
timestamp 1636986456
transform 1 0 8464 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_92
timestamp 18001
transform 1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_115
timestamp 1636986456
transform 1 0 11684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_127
timestamp 1636986456
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_139
timestamp 18001
transform 1 0 13892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 18001
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_189
timestamp 1636986456
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_201
timestamp 1636986456
transform 1 0 19596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 18001
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_241
timestamp 18001
transform 1 0 23276 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_264
timestamp 1636986456
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 18001
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_289
timestamp 1636986456
transform 1 0 27692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_301
timestamp 1636986456
transform 1 0 28796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_313
timestamp 1636986456
transform 1 0 29900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_325
timestamp 18001
transform 1 0 31004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 18001
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_347
timestamp 18001
transform 1 0 33028 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_357
timestamp 1636986456
transform 1 0 33948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_369
timestamp 18001
transform 1 0 35052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_379
timestamp 18001
transform 1 0 35972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 18001
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636986456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 18001
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 18001
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_63
timestamp 18001
transform 1 0 6900 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 18001
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 18001
transform 1 0 9200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_92
timestamp 18001
transform 1 0 9568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 18001
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_122
timestamp 1636986456
transform 1 0 12328 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 18001
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 18001
transform 1 0 15916 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 18001
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636986456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_209
timestamp 18001
transform 1 0 20332 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_217
timestamp 18001
transform 1 0 21068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_242
timestamp 18001
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 18001
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_264
timestamp 1636986456
transform 1 0 25392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_276
timestamp 18001
transform 1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 18001
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 18001
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_336
timestamp 1636986456
transform 1 0 32016 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_348
timestamp 18001
transform 1 0 33120 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 18001
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_368
timestamp 18001
transform 1 0 34960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_378
timestamp 18001
transform 1 0 35880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_384
timestamp 18001
transform 1 0 36432 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 18001
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_34
timestamp 18001
transform 1 0 4232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 18001
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 18001
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_121
timestamp 18001
transform 1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 18001
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_148
timestamp 18001
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 18001
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 18001
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 18001
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_185
timestamp 1636986456
transform 1 0 18124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_197
timestamp 18001
transform 1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 18001
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_238
timestamp 18001
transform 1 0 23000 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_256
timestamp 18001
transform 1 0 24656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 18001
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 18001
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_288
timestamp 18001
transform 1 0 27600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_292
timestamp 18001
transform 1 0 27968 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_306
timestamp 1636986456
transform 1 0 29256 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_318
timestamp 18001
transform 1 0 30360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 18001
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1636986456
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_349
timestamp 18001
transform 1 0 33212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_355
timestamp 18001
transform 1 0 33764 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_372
timestamp 1636986456
transform 1 0 35328 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_384
timestamp 18001
transform 1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 18001
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1636986456
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 18001
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636986456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636986456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_53
timestamp 18001
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 18001
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 18001
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_102
timestamp 1636986456
transform 1 0 10488 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 18001
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 18001
transform 1 0 14352 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_155
timestamp 18001
transform 1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_174
timestamp 18001
transform 1 0 17112 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_182
timestamp 18001
transform 1 0 17848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 18001
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636986456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1636986456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 18001
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_227
timestamp 1636986456
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_239
timestamp 1636986456
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 18001
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 18001
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_259
timestamp 18001
transform 1 0 24932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_267
timestamp 18001
transform 1 0 25668 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1636986456
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_288
timestamp 18001
transform 1 0 27600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_298
timestamp 18001
transform 1 0 28520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 18001
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_309
timestamp 18001
transform 1 0 29532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_319
timestamp 18001
transform 1 0 30452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_325
timestamp 18001
transform 1 0 31004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_331
timestamp 18001
transform 1 0 31556 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_335
timestamp 1636986456
transform 1 0 31924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_347
timestamp 1636986456
transform 1 0 33028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 18001
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 18001
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_372
timestamp 18001
transform 1 0 35328 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_380
timestamp 18001
transform 1 0 36064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_385
timestamp 18001
transform 1 0 36524 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636986456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 18001
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 18001
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 18001
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 18001
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_72
timestamp 18001
transform 1 0 7728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_81
timestamp 18001
transform 1 0 8556 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 18001
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 18001
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 18001
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_127
timestamp 18001
transform 1 0 12788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_154
timestamp 18001
transform 1 0 15272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 18001
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 18001
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 18001
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 18001
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_243
timestamp 18001
transform 1 0 23460 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_248
timestamp 1636986456
transform 1 0 23920 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_263
timestamp 18001
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 18001
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 18001
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1636986456
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_296
timestamp 18001
transform 1 0 28336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_304
timestamp 18001
transform 1 0 29072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_312
timestamp 1636986456
transform 1 0 29808 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_333
timestamp 18001
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_352
timestamp 18001
transform 1 0 33488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_360
timestamp 18001
transform 1 0 34224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1636986456
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 18001
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1636986456
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 18001
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636986456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 18001
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 18001
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 18001
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_156
timestamp 18001
transform 1 0 15456 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_164
timestamp 18001
transform 1 0 16192 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp 18001
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 18001
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636986456
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 18001
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_236
timestamp 18001
transform 1 0 22816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 18001
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_276
timestamp 1636986456
transform 1 0 26496 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_294
timestamp 18001
transform 1 0 28152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 18001
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 18001
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_316
timestamp 18001
transform 1 0 30176 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_320
timestamp 18001
transform 1 0 30544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_325
timestamp 18001
transform 1 0 31004 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_340
timestamp 1636986456
transform 1 0 32384 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_352
timestamp 18001
transform 1 0 33488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_356
timestamp 18001
transform 1 0 33856 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_385
timestamp 18001
transform 1 0 36524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 18001
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_35
timestamp 18001
transform 1 0 4324 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1636986456
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 18001
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 18001
transform 1 0 8832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_121
timestamp 18001
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_130
timestamp 18001
transform 1 0 13064 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_141
timestamp 18001
transform 1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_153
timestamp 1636986456
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 18001
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 18001
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 18001
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 18001
transform 1 0 17388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_201
timestamp 18001
transform 1 0 19596 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 18001
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 18001
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_260
timestamp 18001
transform 1 0 25024 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_271
timestamp 18001
transform 1 0 26036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_293
timestamp 18001
transform 1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_309
timestamp 18001
transform 1 0 29532 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_313
timestamp 18001
transform 1 0 29900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 18001
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_337
timestamp 18001
transform 1 0 32108 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_368
timestamp 1636986456
transform 1 0 34960 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_397
timestamp 18001
transform 1 0 37628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_8
timestamp 18001
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_12
timestamp 18001
transform 1 0 2208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_49
timestamp 18001
transform 1 0 5612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 18001
transform 1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_70
timestamp 18001
transform 1 0 7544 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 18001
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636986456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 18001
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 18001
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 18001
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 18001
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_161
timestamp 18001
transform 1 0 15916 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 18001
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636986456
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_209
timestamp 18001
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_231
timestamp 1636986456
transform 1 0 22356 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_243
timestamp 18001
transform 1 0 23460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 18001
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_259
timestamp 18001
transform 1 0 24932 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_267
timestamp 18001
transform 1 0 25668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_277
timestamp 18001
transform 1 0 26588 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_285
timestamp 18001
transform 1 0 27324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_301
timestamp 18001
transform 1 0 28796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 18001
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_324
timestamp 1636986456
transform 1 0 30912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_336
timestamp 18001
transform 1 0 32016 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_353
timestamp 18001
transform 1 0 33580 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 18001
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 18001
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_369
timestamp 18001
transform 1 0 35052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_385
timestamp 18001
transform 1 0 36524 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636986456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_15
timestamp 18001
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 18001
transform 1 0 3036 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_70
timestamp 18001
transform 1 0 7544 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636986456
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_105
timestamp 18001
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_115
timestamp 18001
transform 1 0 11684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_139
timestamp 1636986456
transform 1 0 13892 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_151
timestamp 1636986456
transform 1 0 14996 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_163
timestamp 18001
transform 1 0 16100 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 18001
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 18001
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 18001
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_232
timestamp 18001
transform 1 0 22448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 18001
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 18001
transform 1 0 23460 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_247
timestamp 18001
transform 1 0 23828 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_255
timestamp 18001
transform 1 0 24564 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_259
timestamp 18001
transform 1 0 24932 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_267
timestamp 18001
transform 1 0 25668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 18001
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_287
timestamp 1636986456
transform 1 0 27508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_299
timestamp 1636986456
transform 1 0 28612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_311
timestamp 18001
transform 1 0 29716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_319
timestamp 18001
transform 1 0 30452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_328
timestamp 18001
transform 1 0 31280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_337
timestamp 18001
transform 1 0 32108 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_350
timestamp 1636986456
transform 1 0 33304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_362
timestamp 18001
transform 1 0 34408 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_368
timestamp 18001
transform 1 0 34960 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 18001
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_400
timestamp 18001
transform 1 0 37904 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_406
timestamp 18001
transform 1 0 38456 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_15
timestamp 18001
transform 1 0 2484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_23
timestamp 18001
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_37
timestamp 18001
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 18001
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_101
timestamp 1636986456
transform 1 0 10396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 18001
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 18001
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_156
timestamp 18001
transform 1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_188
timestamp 18001
transform 1 0 18400 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_192
timestamp 18001
transform 1 0 18768 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 18001
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_218
timestamp 18001
transform 1 0 21160 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_224
timestamp 18001
transform 1 0 21712 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_232
timestamp 18001
transform 1 0 22448 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_243
timestamp 18001
transform 1 0 23460 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 18001
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_269
timestamp 18001
transform 1 0 25852 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_282
timestamp 1636986456
transform 1 0 27048 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_315
timestamp 18001
transform 1 0 30084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_334
timestamp 18001
transform 1 0 31832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_338
timestamp 18001
transform 1 0 32200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_371
timestamp 18001
transform 1 0 35236 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_390
timestamp 1636986456
transform 1 0 36984 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 18001
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 18001
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636986456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_44
timestamp 1636986456
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 18001
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 18001
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 18001
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 18001
transform 1 0 12236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_133
timestamp 18001
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 18001
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 18001
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 18001
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_197
timestamp 18001
transform 1 0 19228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 18001
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636986456
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_237
timestamp 18001
transform 1 0 22908 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_243
timestamp 18001
transform 1 0 23460 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_252
timestamp 1636986456
transform 1 0 24288 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_264
timestamp 18001
transform 1 0 25392 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_272
timestamp 18001
transform 1 0 26128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 18001
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_337
timestamp 18001
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_350
timestamp 1636986456
transform 1 0 33304 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_362
timestamp 1636986456
transform 1 0 34408 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_374
timestamp 18001
transform 1 0 35512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_383
timestamp 18001
transform 1 0 36340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_397
timestamp 18001
transform 1 0 37628 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 18001
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 18001
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 18001
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_19
timestamp 18001
transform 1 0 2852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_34
timestamp 18001
transform 1 0 4232 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_55
timestamp 18001
transform 1 0 6164 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_63
timestamp 18001
transform 1 0 6900 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_69
timestamp 18001
transform 1 0 7452 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 18001
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 18001
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_132
timestamp 18001
transform 1 0 13248 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 18001
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 18001
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_155
timestamp 18001
transform 1 0 15364 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_180
timestamp 18001
transform 1 0 17664 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_188
timestamp 18001
transform 1 0 18400 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 18001
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_201
timestamp 18001
transform 1 0 19596 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 18001
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 18001
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_225
timestamp 18001
transform 1 0 21804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_237
timestamp 18001
transform 1 0 22908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 18001
transform 1 0 25668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_275
timestamp 18001
transform 1 0 26404 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_280
timestamp 18001
transform 1 0 26864 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_286
timestamp 18001
transform 1 0 27416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_291
timestamp 18001
transform 1 0 27876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 18001
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 18001
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_315
timestamp 18001
transform 1 0 30084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_319
timestamp 18001
transform 1 0 30452 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_385
timestamp 18001
transform 1 0 36524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 18001
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_33
timestamp 18001
transform 1 0 4140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_39
timestamp 18001
transform 1 0 4692 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 18001
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_70
timestamp 18001
transform 1 0 7544 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_105
timestamp 18001
transform 1 0 10764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 18001
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 18001
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 18001
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_176
timestamp 18001
transform 1 0 17296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 18001
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 18001
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_262
timestamp 1636986456
transform 1 0 25208 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 18001
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_281
timestamp 18001
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_286
timestamp 18001
transform 1 0 27416 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_297
timestamp 1636986456
transform 1 0 28428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_309
timestamp 18001
transform 1 0 29532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_328
timestamp 18001
transform 1 0 31280 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 18001
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 18001
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_353
timestamp 18001
transform 1 0 33580 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_362
timestamp 18001
transform 1 0 34408 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_383
timestamp 18001
transform 1 0 36340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_387
timestamp 18001
transform 1 0 36708 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_393
timestamp 18001
transform 1 0 37260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_404
timestamp 18001
transform 1 0 38272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 18001
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 18001
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 18001
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 18001
transform 1 0 4048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_51
timestamp 18001
transform 1 0 5796 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_72
timestamp 1636986456
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 18001
transform 1 0 9108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 18001
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_143
timestamp 18001
transform 1 0 14260 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 18001
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_156
timestamp 18001
transform 1 0 15456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_164
timestamp 18001
transform 1 0 16192 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 18001
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_205
timestamp 18001
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_226
timestamp 18001
transform 1 0 21896 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 18001
transform 1 0 25576 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_274
timestamp 18001
transform 1 0 26312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_301
timestamp 18001
transform 1 0 28796 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_350
timestamp 1636986456
transform 1 0 33304 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 18001
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_375
timestamp 18001
transform 1 0 35604 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_31
timestamp 18001
transform 1 0 3956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_39
timestamp 18001
transform 1 0 4692 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_46
timestamp 18001
transform 1 0 5336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 18001
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 18001
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_154
timestamp 1636986456
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 18001
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 18001
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 18001
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_212
timestamp 1636986456
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 18001
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 18001
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_302
timestamp 1636986456
transform 1 0 28888 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_314
timestamp 18001
transform 1 0 29992 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_317
timestamp 18001
transform 1 0 30268 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_323
timestamp 1636986456
transform 1 0 30820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 18001
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 18001
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_365
timestamp 18001
transform 1 0 34684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 18001
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1636986456
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 18001
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636986456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_18
timestamp 18001
transform 1 0 2760 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 18001
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 18001
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 18001
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_45
timestamp 1636986456
transform 1 0 5244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_57
timestamp 1636986456
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1636986456
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 18001
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 18001
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 18001
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_102
timestamp 18001
transform 1 0 10488 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_173
timestamp 18001
transform 1 0 17020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_208
timestamp 18001
transform 1 0 20240 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_231
timestamp 18001
transform 1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_241
timestamp 18001
transform 1 0 23276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_247
timestamp 18001
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 18001
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_271
timestamp 18001
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_279
timestamp 18001
transform 1 0 26772 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_295
timestamp 1636986456
transform 1 0 28244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 18001
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_333
timestamp 18001
transform 1 0 31740 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_341
timestamp 18001
transform 1 0 32476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 18001
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_365
timestamp 18001
transform 1 0 34684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_369
timestamp 18001
transform 1 0 35052 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_374
timestamp 1636986456
transform 1 0 35512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_394
timestamp 18001
transform 1 0 37352 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_402
timestamp 18001
transform 1 0 38088 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 18001
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_11
timestamp 18001
transform 1 0 2116 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_18
timestamp 18001
transform 1 0 2760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 18001
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 18001
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 18001
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 18001
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 18001
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636986456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 18001
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 18001
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 18001
transform 1 0 15180 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 18001
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_177
timestamp 18001
transform 1 0 17388 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_199
timestamp 18001
transform 1 0 19412 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636986456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_237
timestamp 18001
transform 1 0 22908 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_247
timestamp 1636986456
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 18001
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 18001
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_301
timestamp 18001
transform 1 0 28796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_337
timestamp 18001
transform 1 0 32108 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_359
timestamp 1636986456
transform 1 0 34132 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_371
timestamp 1636986456
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_383
timestamp 18001
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 18001
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1636986456
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 18001
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 18001
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_43
timestamp 18001
transform 1 0 5060 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 18001
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_116
timestamp 18001
transform 1 0 11776 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_124
timestamp 18001
transform 1 0 12512 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 18001
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 18001
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 18001
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_149
timestamp 18001
transform 1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_166
timestamp 18001
transform 1 0 16376 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_174
timestamp 18001
transform 1 0 17112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 18001
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_220
timestamp 18001
transform 1 0 21344 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 18001
transform 1 0 22080 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 18001
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 18001
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 18001
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_264
timestamp 18001
transform 1 0 25392 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_270
timestamp 18001
transform 1 0 25944 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 18001
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_309
timestamp 18001
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_317
timestamp 18001
transform 1 0 30268 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_330
timestamp 18001
transform 1 0 31464 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_343
timestamp 18001
transform 1 0 32660 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1636986456
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1636986456
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1636986456
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 18001
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 18001
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_11
timestamp 18001
transform 1 0 2116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 18001
transform 1 0 3588 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_44
timestamp 18001
transform 1 0 5152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 18001
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 18001
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 18001
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 18001
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_122
timestamp 18001
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 18001
transform 1 0 13248 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_136
timestamp 18001
transform 1 0 13616 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_143
timestamp 18001
transform 1 0 14260 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_154
timestamp 1636986456
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 18001
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636986456
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_181
timestamp 18001
transform 1 0 17756 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_187
timestamp 18001
transform 1 0 18308 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_199
timestamp 18001
transform 1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 18001
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 18001
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 18001
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 18001
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_240
timestamp 18001
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_244
timestamp 18001
transform 1 0 23552 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_267
timestamp 18001
transform 1 0 25668 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 18001
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_290
timestamp 18001
transform 1 0 27784 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_298
timestamp 18001
transform 1 0 28520 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_309
timestamp 18001
transform 1 0 29532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_330
timestamp 18001
transform 1 0 31464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_356
timestamp 18001
transform 1 0 33856 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_384
timestamp 18001
transform 1 0 36432 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1636986456
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 18001
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 18001
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp 18001
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 18001
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 18001
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_63
timestamp 18001
transform 1 0 6900 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 18001
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_126
timestamp 18001
transform 1 0 12696 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_130
timestamp 18001
transform 1 0 13064 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_161
timestamp 18001
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 18001
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_204
timestamp 1636986456
transform 1 0 19872 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_216
timestamp 18001
transform 1 0 20976 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 18001
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_262
timestamp 18001
transform 1 0 25208 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_285
timestamp 18001
transform 1 0 27324 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 18001
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 18001
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_313
timestamp 18001
transform 1 0 29900 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_326
timestamp 18001
transform 1 0 31096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_355
timestamp 18001
transform 1 0 33764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_365
timestamp 18001
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_394
timestamp 1636986456
transform 1 0 37352 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 18001
transform 1 0 38456 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 18001
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_38
timestamp 18001
transform 1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636986456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_79
timestamp 18001
transform 1 0 8372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_91
timestamp 18001
transform 1 0 9476 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 18001
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_121
timestamp 18001
transform 1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 18001
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 18001
transform 1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_206
timestamp 1636986456
transform 1 0 20056 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 18001
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 18001
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_234
timestamp 18001
transform 1 0 22632 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_242
timestamp 18001
transform 1 0 23368 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_247
timestamp 18001
transform 1 0 23828 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_254
timestamp 18001
transform 1 0 24472 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_258
timestamp 18001
transform 1 0 24840 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1636986456
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 18001
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp 18001
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_299
timestamp 18001
transform 1 0 28612 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_306
timestamp 18001
transform 1 0 29256 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_321
timestamp 18001
transform 1 0 30636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_325
timestamp 18001
transform 1 0 31004 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 18001
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1636986456
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_374
timestamp 1636986456
transform 1 0 35512 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 18001
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1636986456
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 18001
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636986456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_15
timestamp 18001
transform 1 0 2484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 18001
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_43
timestamp 1636986456
transform 1 0 5060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_55
timestamp 18001
transform 1 0 6164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 18001
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 18001
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 18001
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_107
timestamp 1636986456
transform 1 0 10948 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_119
timestamp 18001
transform 1 0 12052 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 18001
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_144
timestamp 18001
transform 1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_148
timestamp 18001
transform 1 0 14720 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 18001
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 18001
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 18001
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 18001
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 18001
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_257
timestamp 18001
transform 1 0 24748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_268
timestamp 18001
transform 1 0 25760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_276
timestamp 18001
transform 1 0 26496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_291
timestamp 18001
transform 1 0 27876 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_312
timestamp 1636986456
transform 1 0 29808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_324
timestamp 18001
transform 1 0 30912 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_328
timestamp 18001
transform 1 0 31280 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_370
timestamp 18001
transform 1 0 35144 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_394
timestamp 1636986456
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 18001
transform 1 0 38456 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 18001
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_14
timestamp 18001
transform 1 0 2392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_29
timestamp 18001
transform 1 0 3772 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 18001
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 18001
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636986456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_72
timestamp 1636986456
transform 1 0 7728 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_84
timestamp 18001
transform 1 0 8832 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_90
timestamp 18001
transform 1 0 9384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 18001
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 18001
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_172
timestamp 1636986456
transform 1 0 16928 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 18001
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_188
timestamp 18001
transform 1 0 18400 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_196
timestamp 18001
transform 1 0 19136 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_221
timestamp 18001
transform 1 0 21436 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_253
timestamp 18001
transform 1 0 24380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_264
timestamp 18001
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 18001
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 18001
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_298
timestamp 18001
transform 1 0 28520 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_311
timestamp 18001
transform 1 0 29716 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_318
timestamp 1636986456
transform 1 0 30360 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 18001
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_340
timestamp 18001
transform 1 0 32384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_346
timestamp 18001
transform 1 0 32936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_358
timestamp 18001
transform 1 0 34040 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_367
timestamp 18001
transform 1 0 34868 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_373
timestamp 18001
transform 1 0 35420 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1636986456
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 18001
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 18001
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 18001
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 18001
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_125
timestamp 18001
transform 1 0 12604 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 18001
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_182
timestamp 1636986456
transform 1 0 17848 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 18001
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_204
timestamp 1636986456
transform 1 0 19872 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_216
timestamp 18001
transform 1 0 20976 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 18001
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 18001
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636986456
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 18001
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_269
timestamp 18001
transform 1 0 25852 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_277
timestamp 18001
transform 1 0 26588 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_285
timestamp 18001
transform 1 0 27324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_294
timestamp 18001
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 18001
transform 1 0 28520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_302
timestamp 18001
transform 1 0 28888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_335
timestamp 18001
transform 1 0 31924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_339
timestamp 18001
transform 1 0 32292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_343
timestamp 18001
transform 1 0 32660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_351
timestamp 18001
transform 1 0 33396 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 18001
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1636986456
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_377
timestamp 18001
transform 1 0 35788 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_390
timestamp 1636986456
transform 1 0 36984 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 18001
transform 1 0 38088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 18001
transform 1 0 38456 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 18001
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_11
timestamp 18001
transform 1 0 2116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 18001
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 18001
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_94
timestamp 1636986456
transform 1 0 9752 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 18001
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 18001
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_122
timestamp 18001
transform 1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_215
timestamp 18001
transform 1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_264
timestamp 18001
transform 1 0 25392 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_271
timestamp 18001
transform 1 0 26036 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_287
timestamp 18001
transform 1 0 27508 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_294
timestamp 1636986456
transform 1 0 28152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_306
timestamp 18001
transform 1 0 29256 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_312
timestamp 18001
transform 1 0 29808 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1636986456
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 18001
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 18001
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1636986456
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_349
timestamp 18001
transform 1 0 33212 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_363
timestamp 18001
transform 1 0 34500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_371
timestamp 18001
transform 1 0 35236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 18001
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_400
timestamp 18001
transform 1 0 37904 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 18001
transform 1 0 38456 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636986456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_15
timestamp 18001
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 18001
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_50
timestamp 1636986456
transform 1 0 5704 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_62
timestamp 18001
transform 1 0 6808 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 18001
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636986456
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 18001
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_121
timestamp 18001
transform 1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 18001
transform 1 0 12604 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 18001
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_165
timestamp 18001
transform 1 0 16284 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_192
timestamp 18001
transform 1 0 18768 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 18001
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_221
timestamp 18001
transform 1 0 21436 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_242
timestamp 18001
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 18001
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_288
timestamp 18001
transform 1 0 27600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 18001
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_317
timestamp 1636986456
transform 1 0 30268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_348
timestamp 18001
transform 1 0 33120 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 18001
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1636986456
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_389
timestamp 18001
transform 1 0 36892 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_393
timestamp 18001
transform 1 0 37260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 18001
transform 1 0 38456 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636986456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636986456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp 18001
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_34
timestamp 18001
transform 1 0 4232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 18001
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_60
timestamp 1636986456
transform 1 0 6624 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_72
timestamp 18001
transform 1 0 7728 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 18001
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_140
timestamp 18001
transform 1 0 13984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_162
timestamp 18001
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 18001
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_188
timestamp 1636986456
transform 1 0 18400 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_200
timestamp 18001
transform 1 0 19504 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 18001
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_235
timestamp 1636986456
transform 1 0 22724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_247
timestamp 18001
transform 1 0 23828 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 18001
transform 1 0 24564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_273
timestamp 18001
transform 1 0 26220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 18001
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_284
timestamp 1636986456
transform 1 0 27232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_296
timestamp 18001
transform 1 0 28336 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_305
timestamp 18001
transform 1 0 29164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_309
timestamp 18001
transform 1 0 29532 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_313
timestamp 18001
transform 1 0 29900 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_319
timestamp 1636986456
transform 1 0 30452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 18001
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 18001
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_344
timestamp 1636986456
transform 1 0 32752 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_359
timestamp 18001
transform 1 0 34132 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1636986456
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 18001
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 18001
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1636986456
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 18001
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636986456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_15
timestamp 18001
transform 1 0 2484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 18001
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 18001
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 18001
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_47
timestamp 18001
transform 1 0 5428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_69
timestamp 18001
transform 1 0 7452 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_75
timestamp 18001
transform 1 0 8004 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 18001
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_93
timestamp 18001
transform 1 0 9660 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 18001
transform 1 0 10212 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 18001
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 18001
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 18001
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 18001
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_203
timestamp 18001
transform 1 0 19780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_212
timestamp 18001
transform 1 0 20608 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_226
timestamp 18001
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 18001
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636986456
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636986456
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_277
timestamp 18001
transform 1 0 26588 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_284
timestamp 18001
transform 1 0 27232 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_292
timestamp 18001
transform 1 0 27968 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_296
timestamp 18001
transform 1 0 28336 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_300
timestamp 18001
transform 1 0 28704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_309
timestamp 18001
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_320
timestamp 1636986456
transform 1 0 30544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 18001
transform 1 0 31648 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_344
timestamp 18001
transform 1 0 32752 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_350
timestamp 18001
transform 1 0 33304 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_358
timestamp 18001
transform 1 0 34040 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_375
timestamp 18001
transform 1 0 35604 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_383
timestamp 18001
transform 1 0 36340 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_390
timestamp 18001
transform 1 0 36984 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_400
timestamp 18001
transform 1 0 37904 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 18001
transform 1 0 38456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 18001
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_9
timestamp 18001
transform 1 0 1932 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_60
timestamp 18001
transform 1 0 6624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 18001
transform 1 0 8556 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_87
timestamp 1636986456
transform 1 0 9108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_99
timestamp 1636986456
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 18001
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 18001
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_136
timestamp 1636986456
transform 1 0 13616 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_148
timestamp 1636986456
transform 1 0 14720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 18001
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636986456
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636986456
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 18001
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_205
timestamp 18001
transform 1 0 19964 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_210
timestamp 18001
transform 1 0 20424 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 18001
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 18001
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_234
timestamp 18001
transform 1 0 22632 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_260
timestamp 18001
transform 1 0 25024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_265
timestamp 18001
transform 1 0 25484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 18001
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_295
timestamp 18001
transform 1 0 28244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_310
timestamp 18001
transform 1 0 29624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_326
timestamp 18001
transform 1 0 31096 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 18001
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_340
timestamp 18001
transform 1 0 32384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_357
timestamp 18001
transform 1 0 33948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_361
timestamp 18001
transform 1 0 34316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_365
timestamp 18001
transform 1 0 34684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_375
timestamp 18001
transform 1 0 35604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 18001
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_393
timestamp 18001
transform 1 0 37260 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 18001
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 18001
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_14
timestamp 18001
transform 1 0 2392 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 18001
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 18001
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 18001
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_56
timestamp 18001
transform 1 0 6256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_66
timestamp 1636986456
transform 1 0 7176 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_105
timestamp 1636986456
transform 1 0 10764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_117
timestamp 18001
transform 1 0 11868 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_120
timestamp 1636986456
transform 1 0 12144 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 18001
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636986456
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_153
timestamp 18001
transform 1 0 15180 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_168
timestamp 1636986456
transform 1 0 16560 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_180
timestamp 18001
transform 1 0 17664 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_188
timestamp 18001
transform 1 0 18400 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_197
timestamp 18001
transform 1 0 19228 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_212
timestamp 18001
transform 1 0 20608 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_238
timestamp 18001
transform 1 0 23000 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_246
timestamp 18001
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_276
timestamp 18001
transform 1 0 26496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 18001
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 18001
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_316
timestamp 1636986456
transform 1 0 30176 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_328
timestamp 18001
transform 1 0 31280 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_338
timestamp 18001
transform 1 0 32200 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_351
timestamp 1636986456
transform 1 0 33396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 18001
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1636986456
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_377
timestamp 18001
transform 1 0 35788 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 18001
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_28
timestamp 18001
transform 1 0 3680 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_34
timestamp 1636986456
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_46
timestamp 18001
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 18001
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636986456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 18001
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 18001
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_89
timestamp 18001
transform 1 0 9292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 18001
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_115
timestamp 1636986456
transform 1 0 11684 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_127
timestamp 18001
transform 1 0 12788 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_133
timestamp 18001
transform 1 0 13340 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_140
timestamp 18001
transform 1 0 13984 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_152
timestamp 1636986456
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 18001
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 18001
transform 1 0 16928 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_187
timestamp 18001
transform 1 0 18308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_196
timestamp 18001
transform 1 0 19136 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_212
timestamp 18001
transform 1 0 20608 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 18001
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_230
timestamp 1636986456
transform 1 0 22264 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_242
timestamp 18001
transform 1 0 23368 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_267
timestamp 18001
transform 1 0 25668 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_297
timestamp 18001
transform 1 0 28428 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 18001
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_322
timestamp 18001
transform 1 0 30728 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_330
timestamp 18001
transform 1 0 31464 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 18001
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 18001
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_349
timestamp 18001
transform 1 0 33212 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_365
timestamp 18001
transform 1 0 34684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_372
timestamp 18001
transform 1 0 35328 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_380
timestamp 18001
transform 1 0 36064 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_385
timestamp 18001
transform 1 0 36524 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_401
timestamp 18001
transform 1 0 37996 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636986456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_15
timestamp 18001
transform 1 0 2484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_19
timestamp 18001
transform 1 0 2852 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 18001
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_43
timestamp 18001
transform 1 0 5060 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_74
timestamp 18001
transform 1 0 7912 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 18001
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 18001
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 18001
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_98
timestamp 18001
transform 1 0 10120 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_119
timestamp 18001
transform 1 0 12052 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 18001
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_162
timestamp 18001
transform 1 0 16008 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_173
timestamp 18001
transform 1 0 17020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_181
timestamp 18001
transform 1 0 17756 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_185
timestamp 18001
transform 1 0 18124 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 18001
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_208
timestamp 1636986456
transform 1 0 20240 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_227
timestamp 18001
transform 1 0 21988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_235
timestamp 18001
transform 1 0 22724 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 18001
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 18001
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_290
timestamp 18001
transform 1 0 27784 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 18001
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_319
timestamp 18001
transform 1 0 30452 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_336
timestamp 18001
transform 1 0 32016 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_345
timestamp 18001
transform 1 0 32844 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_353
timestamp 18001
transform 1 0 33580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 18001
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_365
timestamp 18001
transform 1 0 34684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_385
timestamp 18001
transform 1 0 36524 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_398
timestamp 18001
transform 1 0 37720 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 18001
transform 1 0 38456 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_25
timestamp 18001
transform 1 0 3404 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_34
timestamp 18001
transform 1 0 4232 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_72
timestamp 18001
transform 1 0 7728 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_76
timestamp 18001
transform 1 0 8096 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 18001
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_121
timestamp 18001
transform 1 0 12236 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_134
timestamp 18001
transform 1 0 13432 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_149
timestamp 18001
transform 1 0 14812 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_161
timestamp 18001
transform 1 0 15916 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 18001
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636986456
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 18001
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_197
timestamp 1636986456
transform 1 0 19228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_209
timestamp 18001
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_217
timestamp 18001
transform 1 0 21068 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 18001
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_237
timestamp 18001
transform 1 0 22908 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 18001
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_288
timestamp 1636986456
transform 1 0 27600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_300
timestamp 18001
transform 1 0 28704 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_310
timestamp 18001
transform 1 0 29624 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_318
timestamp 18001
transform 1 0 30360 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 18001
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_347
timestamp 18001
transform 1 0 33028 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_358
timestamp 18001
transform 1 0 34040 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_368
timestamp 18001
transform 1 0 34960 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_380
timestamp 18001
transform 1 0 36064 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_386
timestamp 18001
transform 1 0 36616 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 18001
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1636986456
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 18001
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_57
timestamp 18001
transform 1 0 6348 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_66
timestamp 18001
transform 1 0 7176 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 18001
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 18001
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 18001
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_102
timestamp 18001
transform 1 0 10488 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 18001
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 18001
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_149
timestamp 18001
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_166
timestamp 1636986456
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_178
timestamp 18001
transform 1 0 17480 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 18001
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 18001
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 18001
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_203
timestamp 18001
transform 1 0 19780 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_212
timestamp 18001
transform 1 0 20608 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 18001
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 18001
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 18001
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 18001
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_262
timestamp 18001
transform 1 0 25208 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 18001
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 18001
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 18001
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_318
timestamp 18001
transform 1 0 30360 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_346
timestamp 18001
transform 1 0 32936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 18001
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 18001
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_370
timestamp 1636986456
transform 1 0 35144 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_382
timestamp 18001
transform 1 0 36248 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 18001
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636986456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_15
timestamp 18001
transform 1 0 2484 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_26
timestamp 1636986456
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_38
timestamp 18001
transform 1 0 4600 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_46
timestamp 18001
transform 1 0 5336 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 18001
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_65
timestamp 18001
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_90
timestamp 18001
transform 1 0 9384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 18001
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 18001
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_121
timestamp 18001
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 18001
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_149
timestamp 18001
transform 1 0 14812 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 18001
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 18001
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_177
timestamp 18001
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_184
timestamp 18001
transform 1 0 18032 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_206
timestamp 18001
transform 1 0 20056 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 18001
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_233
timestamp 18001
transform 1 0 22540 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_265
timestamp 1636986456
transform 1 0 25484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 18001
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 18001
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_287
timestamp 18001
transform 1 0 27508 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_292
timestamp 18001
transform 1 0 27968 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_356
timestamp 18001
transform 1 0 33856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_362
timestamp 18001
transform 1 0 34408 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_368
timestamp 18001
transform 1 0 34960 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_383
timestamp 18001
transform 1 0 36340 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 18001
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 18001
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_400
timestamp 18001
transform 1 0 37904 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 18001
transform 1 0 38456 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636986456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_15
timestamp 18001
transform 1 0 2484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 18001
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_32
timestamp 18001
transform 1 0 4048 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 18001
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_98
timestamp 18001
transform 1 0 10120 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_119
timestamp 18001
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_127
timestamp 18001
transform 1 0 12788 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_133
timestamp 18001
transform 1 0 13340 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_149
timestamp 18001
transform 1 0 14812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_153
timestamp 18001
transform 1 0 15180 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_157
timestamp 18001
transform 1 0 15548 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_168
timestamp 18001
transform 1 0 16560 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_184
timestamp 18001
transform 1 0 18032 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 18001
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 18001
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_217
timestamp 1636986456
transform 1 0 21068 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_229
timestamp 1636986456
transform 1 0 22172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_241
timestamp 18001
transform 1 0 23276 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_262
timestamp 18001
transform 1 0 25208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 18001
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_322
timestamp 18001
transform 1 0 30728 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_328
timestamp 1636986456
transform 1 0 31280 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_340
timestamp 1636986456
transform 1 0 32384 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_352
timestamp 1636986456
transform 1 0 33488 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 18001
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_375
timestamp 18001
transform 1 0 35604 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_386
timestamp 18001
transform 1 0 36616 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_394
timestamp 18001
transform 1 0 37352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 18001
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_16
timestamp 18001
transform 1 0 2576 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636986456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_69
timestamp 18001
transform 1 0 7452 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 18001
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_121
timestamp 18001
transform 1 0 12236 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_131
timestamp 18001
transform 1 0 13156 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_137
timestamp 18001
transform 1 0 13708 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_144
timestamp 18001
transform 1 0 14352 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_155
timestamp 18001
transform 1 0 15364 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 18001
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636986456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636986456
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_198
timestamp 18001
transform 1 0 19320 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_207
timestamp 1636986456
transform 1 0 20148 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 18001
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_228
timestamp 18001
transform 1 0 22080 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_242
timestamp 18001
transform 1 0 23368 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 18001
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_319
timestamp 18001
transform 1 0 30452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 18001
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_337
timestamp 18001
transform 1 0 32108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_346
timestamp 18001
transform 1 0 32936 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_381
timestamp 18001
transform 1 0 36156 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 18001
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_393
timestamp 18001
transform 1 0 37260 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_48
timestamp 1636986456
transform 1 0 5520 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_60
timestamp 18001
transform 1 0 6624 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_66
timestamp 18001
transform 1 0 7176 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_70
timestamp 1636986456
transform 1 0 7544 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 18001
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636986456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_97
timestamp 18001
transform 1 0 10028 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_105
timestamp 18001
transform 1 0 10764 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 18001
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 18001
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_150
timestamp 18001
transform 1 0 14904 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_176
timestamp 18001
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_183
timestamp 18001
transform 1 0 17940 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_187
timestamp 18001
transform 1 0 18308 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_197
timestamp 18001
transform 1 0 19228 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_211
timestamp 18001
transform 1 0 20516 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_244
timestamp 18001
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_258
timestamp 18001
transform 1 0 24840 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_289
timestamp 18001
transform 1 0 27692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 18001
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 18001
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_317
timestamp 18001
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_338
timestamp 18001
transform 1 0 32200 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_350
timestamp 1636986456
transform 1 0 33304 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 18001
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_365
timestamp 18001
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_369
timestamp 18001
transform 1 0 35052 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_373
timestamp 1636986456
transform 1 0 35420 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_385
timestamp 18001
transform 1 0 36524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_389
timestamp 18001
transform 1 0 36892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 18001
transform 1 0 38456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 18001
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_7
timestamp 18001
transform 1 0 1748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 18001
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 18001
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_90
timestamp 18001
transform 1 0 9384 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_98
timestamp 18001
transform 1 0 10120 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_104
timestamp 18001
transform 1 0 10672 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 18001
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 18001
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_178
timestamp 18001
transform 1 0 17480 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_188
timestamp 1636986456
transform 1 0 18400 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_209
timestamp 18001
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_213
timestamp 18001
transform 1 0 20700 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 18001
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_230
timestamp 18001
transform 1 0 22264 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_249
timestamp 18001
transform 1 0 24012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 18001
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_289
timestamp 18001
transform 1 0 27692 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_318
timestamp 18001
transform 1 0 30360 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_325
timestamp 18001
transform 1 0 31004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_329
timestamp 18001
transform 1 0 31372 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_337
timestamp 18001
transform 1 0 32108 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_364
timestamp 1636986456
transform 1 0 34592 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_376
timestamp 1636986456
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 18001
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_404
timestamp 18001
transform 1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_15
timestamp 18001
transform 1 0 2484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_19
timestamp 18001
transform 1 0 2852 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 18001
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 18001
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 18001
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_141
timestamp 18001
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_164
timestamp 18001
transform 1 0 16192 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_172
timestamp 18001
transform 1 0 16928 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1636986456
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1636986456
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_221
timestamp 18001
transform 1 0 21436 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_227
timestamp 18001
transform 1 0 21988 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_239
timestamp 18001
transform 1 0 23092 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 18001
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_270
timestamp 18001
transform 1 0 25944 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 18001
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_329
timestamp 1636986456
transform 1 0 31372 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_341
timestamp 18001
transform 1 0 32476 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_350
timestamp 18001
transform 1 0 33304 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_361
timestamp 18001
transform 1 0 34316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_365
timestamp 18001
transform 1 0 34684 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_386
timestamp 18001
transform 1 0 36616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 18001
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_6
timestamp 18001
transform 1 0 1656 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_35
timestamp 18001
transform 1 0 4324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 18001
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_61
timestamp 18001
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 18001
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_126
timestamp 18001
transform 1 0 12696 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 18001
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 18001
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1636986456
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 18001
transform 1 0 17756 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_189
timestamp 18001
transform 1 0 18492 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 18001
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 18001
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_241
timestamp 18001
transform 1 0 23276 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 18001
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_289
timestamp 18001
transform 1 0 27692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_312
timestamp 18001
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_337
timestamp 18001
transform 1 0 32108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_348
timestamp 18001
transform 1 0 33120 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_375
timestamp 18001
transform 1 0 35604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_383
timestamp 18001
transform 1 0 36340 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_400
timestamp 18001
transform 1 0 37904 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 18001
transform 1 0 38456 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_6
timestamp 1636986456
transform 1 0 1656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_18
timestamp 18001
transform 1 0 2760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_44
timestamp 18001
transform 1 0 5152 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_54
timestamp 18001
transform 1 0 6072 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_105
timestamp 18001
transform 1 0 10764 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_115
timestamp 18001
transform 1 0 11684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 18001
transform 1 0 12236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_130
timestamp 18001
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 18001
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_141
timestamp 18001
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_152
timestamp 18001
transform 1 0 15088 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_181
timestamp 18001
transform 1 0 17756 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_189
timestamp 18001
transform 1 0 18492 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 18001
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_197
timestamp 18001
transform 1 0 19228 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_221
timestamp 18001
transform 1 0 21436 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_240
timestamp 18001
transform 1 0 23184 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 18001
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_261
timestamp 18001
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_291
timestamp 18001
transform 1 0 27876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_297
timestamp 18001
transform 1 0 28428 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 18001
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_329
timestamp 1636986456
transform 1 0 31372 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_341
timestamp 18001
transform 1 0 32476 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_351
timestamp 18001
transform 1 0 33396 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_385
timestamp 18001
transform 1 0 36524 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_391
timestamp 1636986456
transform 1 0 37076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 18001
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_6
timestamp 1636986456
transform 1 0 1656 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_18
timestamp 18001
transform 1 0 2760 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_26
timestamp 18001
transform 1 0 3496 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_33
timestamp 18001
transform 1 0 4140 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_41
timestamp 18001
transform 1 0 4876 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 18001
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 18001
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_64
timestamp 18001
transform 1 0 6992 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_90
timestamp 18001
transform 1 0 9384 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_95
timestamp 18001
transform 1 0 9844 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_107
timestamp 18001
transform 1 0 10948 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 18001
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 18001
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_121
timestamp 18001
transform 1 0 12236 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_148
timestamp 18001
transform 1 0 14720 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_196
timestamp 18001
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_202
timestamp 18001
transform 1 0 19688 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_206
timestamp 18001
transform 1 0 20056 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_216
timestamp 18001
transform 1 0 20976 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_232
timestamp 18001
transform 1 0 22448 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_240
timestamp 18001
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 18001
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_289
timestamp 1636986456
transform 1 0 27692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_301
timestamp 18001
transform 1 0 28796 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 18001
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_337
timestamp 18001
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_347
timestamp 1636986456
transform 1 0 33028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_359
timestamp 18001
transform 1 0 34132 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_380
timestamp 1636986456
transform 1 0 36064 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1636986456
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 18001
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636986456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636986456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_29
timestamp 18001
transform 1 0 3772 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_33
timestamp 18001
transform 1 0 4140 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_39
timestamp 18001
transform 1 0 4692 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_62
timestamp 18001
transform 1 0 6808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_74
timestamp 18001
transform 1 0 7912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 18001
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 18001
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 18001
transform 1 0 9660 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_128
timestamp 18001
transform 1 0 12880 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_132
timestamp 18001
transform 1 0 13248 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_141
timestamp 18001
transform 1 0 14076 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_148
timestamp 18001
transform 1 0 14720 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_168
timestamp 18001
transform 1 0 16560 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 18001
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1636986456
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_209
timestamp 18001
transform 1 0 20332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_233
timestamp 18001
transform 1 0 22540 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_238
timestamp 18001
transform 1 0 23000 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_273
timestamp 18001
transform 1 0 26220 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_282
timestamp 1636986456
transform 1 0 27048 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_294
timestamp 1636986456
transform 1 0 28152 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 18001
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_309
timestamp 18001
transform 1 0 29532 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_330
timestamp 18001
transform 1 0 31464 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_336
timestamp 18001
transform 1 0 32016 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_393
timestamp 18001
transform 1 0 37260 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_401
timestamp 18001
transform 1 0 37996 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636986456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_15
timestamp 18001
transform 1 0 2484 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_23
timestamp 18001
transform 1 0 3220 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 18001
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_64
timestamp 18001
transform 1 0 6992 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_92
timestamp 1636986456
transform 1 0 9568 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 18001
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_120
timestamp 18001
transform 1 0 12144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_128
timestamp 18001
transform 1 0 12880 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_150
timestamp 18001
transform 1 0 14904 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_156
timestamp 18001
transform 1 0 15456 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 18001
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_169
timestamp 18001
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_180
timestamp 18001
transform 1 0 17664 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_211
timestamp 1636986456
transform 1 0 20516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 18001
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_258
timestamp 18001
transform 1 0 24840 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 18001
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_305
timestamp 18001
transform 1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_316
timestamp 18001
transform 1 0 30176 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_322
timestamp 1636986456
transform 1 0 30728 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 18001
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_337
timestamp 18001
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_341
timestamp 18001
transform 1 0 32476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_347
timestamp 18001
transform 1 0 33028 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_355
timestamp 18001
transform 1 0 33764 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 18001
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1636986456
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 18001
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 18001
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_7
timestamp 18001
transform 1 0 1748 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 18001
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_46
timestamp 18001
transform 1 0 5336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_63
timestamp 18001
transform 1 0 6900 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_78
timestamp 18001
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1636986456
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_97
timestamp 18001
transform 1 0 10028 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_102
timestamp 18001
transform 1 0 10488 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_126
timestamp 1636986456
transform 1 0 12696 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 18001
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 18001
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_164
timestamp 18001
transform 1 0 16192 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_172
timestamp 18001
transform 1 0 16928 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_183
timestamp 18001
transform 1 0 17940 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_217
timestamp 18001
transform 1 0 21068 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 18001
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_261
timestamp 18001
transform 1 0 25116 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_271
timestamp 18001
transform 1 0 26036 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_275
timestamp 18001
transform 1 0 26404 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_300
timestamp 18001
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_309
timestamp 18001
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_317
timestamp 18001
transform 1 0 30268 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_338
timestamp 18001
transform 1 0 32200 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_350
timestamp 1636986456
transform 1 0 33304 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 18001
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 18001
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_373
timestamp 18001
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_382
timestamp 1636986456
transform 1 0 36248 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_394
timestamp 18001
transform 1 0 37352 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_402
timestamp 18001
transform 1 0 38088 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636986456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636986456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_27
timestamp 18001
transform 1 0 3588 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_48
timestamp 18001
transform 1 0 5520 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_57
timestamp 18001
transform 1 0 6348 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_67
timestamp 1636986456
transform 1 0 7268 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_79
timestamp 1636986456
transform 1 0 8372 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_91
timestamp 18001
transform 1 0 9476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_113
timestamp 18001
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_136
timestamp 18001
transform 1 0 13616 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_140
timestamp 18001
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_164
timestamp 18001
transform 1 0 16192 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_199
timestamp 1636986456
transform 1 0 19412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_211
timestamp 1636986456
transform 1 0 20516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 18001
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 18001
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_258
timestamp 18001
transform 1 0 24840 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_270
timestamp 18001
transform 1 0 25944 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 18001
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 18001
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_315
timestamp 18001
transform 1 0 30084 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_323
timestamp 18001
transform 1 0 30820 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 18001
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_342
timestamp 18001
transform 1 0 32568 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_365
timestamp 1636986456
transform 1 0 34684 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_377
timestamp 1636986456
transform 1 0 35788 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_389
timestamp 18001
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1636986456
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 18001
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_15
timestamp 18001
transform 1 0 2484 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_23
timestamp 18001
transform 1 0 3220 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_29
timestamp 18001
transform 1 0 3772 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_75
timestamp 18001
transform 1 0 8004 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 18001
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_125
timestamp 1636986456
transform 1 0 12604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 18001
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_141
timestamp 18001
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_155
timestamp 18001
transform 1 0 15364 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_167
timestamp 18001
transform 1 0 16468 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 18001
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_210
timestamp 1636986456
transform 1 0 20424 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_222
timestamp 18001
transform 1 0 21528 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_230
timestamp 18001
transform 1 0 22264 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_242
timestamp 18001
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 18001
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_285
timestamp 18001
transform 1 0 27324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_293
timestamp 18001
transform 1 0 28060 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_325
timestamp 18001
transform 1 0 31004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 18001
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_388
timestamp 1636986456
transform 1 0 36800 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_400
timestamp 18001
transform 1 0 37904 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 18001
transform 1 0 38456 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_3
timestamp 18001
transform 1 0 1380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_11
timestamp 18001
transform 1 0 2116 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_32
timestamp 18001
transform 1 0 4048 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_42
timestamp 18001
transform 1 0 4968 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 18001
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_57
timestamp 18001
transform 1 0 6348 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_68
timestamp 18001
transform 1 0 7360 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_92
timestamp 18001
transform 1 0 9568 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1636986456
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1636986456
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1636986456
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_149
timestamp 18001
transform 1 0 14812 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 18001
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1636986456
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_181
timestamp 18001
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_189
timestamp 18001
transform 1 0 18492 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_248
timestamp 18001
transform 1 0 23920 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_256
timestamp 18001
transform 1 0 24656 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 18001
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_281
timestamp 18001
transform 1 0 26956 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 18001
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1636986456
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_377
timestamp 1636986456
transform 1 0 35788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_389
timestamp 18001
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 18001
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_401
timestamp 18001
transform 1 0 37996 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_15
timestamp 18001
transform 1 0 2484 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_21
timestamp 18001
transform 1 0 3036 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 18001
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_52
timestamp 18001
transform 1 0 5888 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_60
timestamp 18001
transform 1 0 6624 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_66
timestamp 1636986456
transform 1 0 7176 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_78
timestamp 18001
transform 1 0 8280 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_85
timestamp 18001
transform 1 0 8924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_108
timestamp 18001
transform 1 0 11040 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 18001
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_141
timestamp 18001
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_149
timestamp 18001
transform 1 0 14812 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_155
timestamp 18001
transform 1 0 15364 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 18001
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_246
timestamp 18001
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 18001
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1636986456
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_277
timestamp 18001
transform 1 0 26588 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_285
timestamp 18001
transform 1 0 27324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 18001
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 18001
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_343
timestamp 18001
transform 1 0 32660 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_347
timestamp 18001
transform 1 0 33028 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 18001
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 18001
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1636986456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1636986456
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1636986456
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 18001
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_15
timestamp 18001
transform 1 0 2484 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636986456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1636986456
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_81
timestamp 18001
transform 1 0 8556 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_89
timestamp 18001
transform 1 0 9292 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_97
timestamp 18001
transform 1 0 10028 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_163
timestamp 18001
transform 1 0 16100 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_176
timestamp 18001
transform 1 0 17296 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_197
timestamp 18001
transform 1 0 19228 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 18001
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_259
timestamp 18001
transform 1 0 24932 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 18001
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 18001
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1636986456
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_293
timestamp 18001
transform 1 0 28060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_305
timestamp 18001
transform 1 0 29164 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 18001
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_341
timestamp 18001
transform 1 0 32476 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_345
timestamp 18001
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_359
timestamp 1636986456
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_371
timestamp 1636986456
transform 1 0 35236 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_383
timestamp 18001
transform 1 0 36340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 18001
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 18001
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_401
timestamp 18001
transform 1 0 37996 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_6
timestamp 1636986456
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_18
timestamp 18001
transform 1 0 2760 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 18001
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_29
timestamp 18001
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_55
timestamp 18001
transform 1 0 6164 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_59
timestamp 18001
transform 1 0 6532 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1636986456
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_97
timestamp 18001
transform 1 0 10028 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_133
timestamp 18001
transform 1 0 13340 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 18001
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_149
timestamp 18001
transform 1 0 14812 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_159
timestamp 18001
transform 1 0 15732 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_169
timestamp 18001
transform 1 0 16652 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_177
timestamp 18001
transform 1 0 17388 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_188
timestamp 18001
transform 1 0 18400 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1636986456
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_209
timestamp 18001
transform 1 0 20332 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_230
timestamp 18001
transform 1 0 22264 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_238
timestamp 18001
transform 1 0 23000 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_268
timestamp 1636986456
transform 1 0 25760 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_280
timestamp 18001
transform 1 0 26864 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_290
timestamp 18001
transform 1 0 27784 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_296
timestamp 1636986456
transform 1 0 28336 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_312
timestamp 18001
transform 1 0 29808 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_319
timestamp 18001
transform 1 0 30452 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_355
timestamp 18001
transform 1 0 33764 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 18001
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1636986456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1636986456
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1636986456
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_401
timestamp 18001
transform 1 0 37996 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_6
timestamp 1636986456
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_18
timestamp 1636986456
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_46
timestamp 18001
transform 1 0 5336 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 18001
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_99
timestamp 1636986456
transform 1 0 10212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 18001
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1636986456
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_125
timestamp 18001
transform 1 0 12604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_129
timestamp 18001
transform 1 0 12972 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_134
timestamp 1636986456
transform 1 0 13432 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_146
timestamp 1636986456
transform 1 0 14536 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_158
timestamp 18001
transform 1 0 15640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 18001
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1636986456
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1636986456
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 18001
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_210
timestamp 18001
transform 1 0 20424 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 18001
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1636986456
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_237
timestamp 18001
transform 1 0 22908 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_270
timestamp 18001
transform 1 0 25944 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 18001
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_301
timestamp 18001
transform 1 0 28796 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 18001
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1636986456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1636986456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1636986456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1636986456
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 18001
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 18001
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 18001
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_401
timestamp 18001
transform 1 0 37996 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_6
timestamp 1636986456
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_18
timestamp 18001
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 18001
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_29
timestamp 18001
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_35
timestamp 18001
transform 1 0 4324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_43
timestamp 18001
transform 1 0 5060 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 18001
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_93
timestamp 1636986456
transform 1 0 9660 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_105
timestamp 1636986456
transform 1 0 10764 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_117
timestamp 1636986456
transform 1 0 11868 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_129
timestamp 18001
transform 1 0 12972 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 18001
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1636986456
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1636986456
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1636986456
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1636986456
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 18001
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 18001
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_237
timestamp 18001
transform 1 0 22908 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_256
timestamp 18001
transform 1 0 24656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_266
timestamp 18001
transform 1 0 25576 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_275
timestamp 18001
transform 1 0 26404 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_283
timestamp 18001
transform 1 0 27140 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_299
timestamp 18001
transform 1 0 28612 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_317
timestamp 18001
transform 1 0 30268 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_339
timestamp 1636986456
transform 1 0 32292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_351
timestamp 1636986456
transform 1 0 33396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 18001
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1636986456
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1636986456
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1636986456
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_401
timestamp 18001
transform 1 0 37996 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_27
timestamp 18001
transform 1 0 3588 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_35
timestamp 18001
transform 1 0 4324 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 18001
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_61
timestamp 18001
transform 1 0 6716 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_86
timestamp 1636986456
transform 1 0 9016 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_98
timestamp 1636986456
transform 1 0 10120 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 18001
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1636986456
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1636986456
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1636986456
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1636986456
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 18001
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 18001
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1636986456
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1636986456
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_193
timestamp 18001
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_225
timestamp 18001
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_254
timestamp 18001
transform 1 0 24472 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 18001
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_284
timestamp 18001
transform 1 0 27232 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_328
timestamp 18001
transform 1 0 31280 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1636986456
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1636986456
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1636986456
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1636986456
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 18001
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 18001
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 18001
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_9
timestamp 1636986456
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_21
timestamp 18001
transform 1 0 3036 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 18001
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 18001
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_57
timestamp 1636986456
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_69
timestamp 18001
transform 1 0 7452 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 18001
transform 1 0 8372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 18001
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1636986456
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1636986456
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 18001
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1636986456
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1636986456
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 18001
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1636986456
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1636986456
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 18001
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1636986456
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_181
timestamp 1636986456
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 18001
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1636986456
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_209
timestamp 18001
transform 1 0 20332 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_217
timestamp 18001
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 18001
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1636986456
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_237
timestamp 18001
transform 1 0 22908 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_245
timestamp 18001
transform 1 0 23644 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1636986456
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_268
timestamp 18001
transform 1 0 25760 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_273
timestamp 18001
transform 1 0 26220 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 18001
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 18001
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 18001
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_300
timestamp 18001
transform 1 0 28704 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 18001
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 18001
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 18001
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 18001
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_328
timestamp 18001
transform 1 0 31280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 18001
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 18001
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_342
timestamp 18001
transform 1 0 32568 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_349
timestamp 18001
transform 1 0 33212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_356
timestamp 18001
transform 1 0 33856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 18001
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 18001
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 18001
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 18001
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_384
timestamp 18001
transform 1 0 36432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 18001
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_393
timestamp 18001
transform 1 0 37260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_397
timestamp 18001
transform 1 0 37628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 18001
transform -1 0 8832 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 18001
transform -1 0 18952 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 18001
transform -1 0 3680 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 18001
transform -1 0 8648 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 18001
transform -1 0 7636 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 18001
transform -1 0 25024 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 18001
transform -1 0 24104 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 18001
transform -1 0 25116 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 18001
transform -1 0 25116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 18001
transform -1 0 24104 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 18001
transform 1 0 10580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 18001
transform -1 0 10580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 18001
transform -1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 18001
transform -1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 18001
transform -1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 18001
transform -1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 18001
transform 1 0 5060 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 18001
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 18001
transform -1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 18001
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 18001
transform -1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 18001
transform -1 0 8740 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 18001
transform -1 0 8740 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 18001
transform -1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 18001
transform 1 0 25300 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 18001
transform 1 0 26312 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 18001
transform -1 0 9936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 18001
transform -1 0 9384 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 18001
transform 1 0 8464 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 18001
transform -1 0 5152 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 18001
transform -1 0 10948 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 18001
transform -1 0 30268 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 18001
transform -1 0 8832 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 18001
transform -1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 18001
transform -1 0 23368 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 18001
transform -1 0 8372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 18001
transform -1 0 13340 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 18001
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 18001
transform 1 0 9476 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 18001
transform -1 0 25484 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 18001
transform -1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 18001
transform -1 0 3404 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 18001
transform -1 0 3680 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 18001
transform -1 0 3496 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 18001
transform 1 0 31188 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 18001
transform -1 0 8372 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 18001
transform -1 0 19412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 18001
transform -1 0 15732 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 18001
transform -1 0 4600 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 18001
transform -1 0 15088 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 18001
transform -1 0 8280 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 18001
transform -1 0 5888 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 18001
transform 1 0 3956 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 18001
transform -1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 18001
transform -1 0 5888 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 18001
transform -1 0 6256 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 18001
transform -1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 18001
transform -1 0 21344 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 18001
transform -1 0 4692 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 18001
transform -1 0 6072 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 18001
transform -1 0 9660 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 18001
transform -1 0 8740 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 18001
transform -1 0 7544 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 18001
transform -1 0 28428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 18001
transform -1 0 28060 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 18001
transform -1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 18001
transform -1 0 26772 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 18001
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 18001
transform -1 0 38548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 18001
transform -1 0 27692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 18001
transform 1 0 23460 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 18001
transform -1 0 7360 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 18001
transform -1 0 36248 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 18001
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 18001
transform -1 0 11684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 18001
transform -1 0 26680 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 18001
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 18001
transform -1 0 6624 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 18001
transform -1 0 21436 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 18001
transform -1 0 21896 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 18001
transform -1 0 7268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 18001
transform -1 0 16836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 18001
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 18001
transform -1 0 35788 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 18001
transform -1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 18001
transform 1 0 4048 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 18001
transform 1 0 3956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 18001
transform -1 0 28428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 18001
transform 1 0 26956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 18001
transform -1 0 27692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 18001
transform -1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 18001
transform -1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 18001
transform -1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 18001
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 18001
transform -1 0 26404 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 18001
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 18001
transform -1 0 6716 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 18001
transform -1 0 16468 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 18001
transform -1 0 12236 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 18001
transform -1 0 25576 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 18001
transform -1 0 12420 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 18001
transform -1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 18001
transform -1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 18001
transform -1 0 13984 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 18001
transform 1 0 4048 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 18001
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 18001
transform -1 0 11316 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 18001
transform 1 0 9844 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 18001
transform -1 0 12236 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 18001
transform -1 0 9660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 18001
transform -1 0 6808 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 18001
transform -1 0 3956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 18001
transform -1 0 7084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 18001
transform -1 0 4232 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 18001
transform -1 0 5980 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 18001
transform -1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 18001
transform -1 0 8648 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 18001
transform 1 0 12420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 18001
transform -1 0 7084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 18001
transform -1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 18001
transform -1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 18001
transform -1 0 18400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 18001
transform -1 0 4784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 18001
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 18001
transform -1 0 23828 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 18001
transform 1 0 10212 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 18001
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 18001
transform -1 0 4416 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 18001
transform -1 0 3680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 18001
transform -1 0 28888 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 18001
transform -1 0 38272 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 18001
transform -1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 18001
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 18001
transform -1 0 12328 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 18001
transform -1 0 4784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 18001
transform 1 0 17756 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 18001
transform -1 0 31832 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 18001
transform 1 0 29716 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 18001
transform -1 0 14812 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 18001
transform -1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 18001
transform 1 0 32292 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 18001
transform -1 0 29256 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 18001
transform -1 0 3680 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 18001
transform -1 0 12420 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 18001
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 18001
transform -1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 18001
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 18001
transform 1 0 9936 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 18001
transform -1 0 17940 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 18001
transform 1 0 15916 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 18001
transform -1 0 34408 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 18001
transform -1 0 9844 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 18001
transform -1 0 12236 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 18001
transform -1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 18001
transform -1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 18001
transform -1 0 14720 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 18001
transform -1 0 8740 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 18001
transform -1 0 15272 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 18001
transform -1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 18001
transform -1 0 17388 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 18001
transform -1 0 37352 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 18001
transform -1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 18001
transform -1 0 14168 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 18001
transform -1 0 18676 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 18001
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 18001
transform -1 0 25208 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 18001
transform -1 0 13616 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 18001
transform -1 0 12236 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 18001
transform -1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 18001
transform 1 0 4232 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 18001
transform 1 0 12880 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 18001
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 18001
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 18001
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap15
timestamp 18001
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap16
timestamp 18001
transform -1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap17
timestamp 18001
transform -1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap29
timestamp 18001
transform -1 0 16928 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 18001
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 18001
transform -1 0 24288 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 18001
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 18001
transform -1 0 26864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 18001
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 18001
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 18001
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_144
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_145
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_146
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_147
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_148
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_149
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_150
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_151
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_152
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_153
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_154
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_155
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_156
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_157
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_158
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_159
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_160
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_161
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_162
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_163
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_164
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_165
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_166
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_167
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_168
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_169
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_170
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_171
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_172
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_173
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_174
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_175
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_176
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_177
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_178
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_179
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_180
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_181
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_182
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_183
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_184
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_185
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_186
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_187
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_188
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_189
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_190
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_191
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_192
timestamp 18001
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_193
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_194
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_195
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_196
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_197
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_198
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_199
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_200
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_201
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_202
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_203
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_204
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_205
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_206
timestamp 18001
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_207
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_208
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_209
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_210
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_211
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_212
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_213
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_214
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_215
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_216
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_217
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_218
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_219
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_220
timestamp 18001
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_221
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_222
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_223
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_224
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_225
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_226
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_227
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_228
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_229
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_230
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_231
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_232
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_233
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_234
timestamp 18001
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_235
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_236
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_237
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_238
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_239
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_240
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_241
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_242
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_243
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_244
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_245
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_246
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_247
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_248
timestamp 18001
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_249
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_250
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_251
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_252
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_253
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_254
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_255
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_256
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_257
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_258
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_259
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_260
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_261
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_262
timestamp 18001
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_263
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_264
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_265
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_266
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_267
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_268
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_269
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_270
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_271
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_272
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_273
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_274
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_275
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_276
timestamp 18001
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_277
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_278
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_279
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_280
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_281
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_282
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_283
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_284
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_285
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_286
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_287
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_288
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_289
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_290
timestamp 18001
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_291
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_292
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_293
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_294
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_295
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_296
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_297
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_298
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_299
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_300
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_301
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_302
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_303
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_304
timestamp 18001
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_305
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_306
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_307
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_308
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_309
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_310
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_311
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_312
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_313
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_314
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_315
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_316
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_317
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_318
timestamp 18001
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_319
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_320
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_321
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_322
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_323
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_324
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_325
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_326
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_327
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_328
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_329
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_330
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_331
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_332
timestamp 18001
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_333
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_334
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_335
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_336
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_337
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_338
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_339
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_340
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_341
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_342
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_343
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_344
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_345
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_346
timestamp 18001
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_347
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_348
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_349
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_350
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_351
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_352
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_353
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_354
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_355
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_356
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_357
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_358
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_359
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_360
timestamp 18001
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_361
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_362
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_363
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_364
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_365
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_366
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_367
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_368
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_369
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_370
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_371
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_372
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_373
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_374
timestamp 18001
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_375
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_376
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_377
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_378
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_379
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_380
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_381
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_382
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_383
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_384
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_385
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_386
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_387
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_388
timestamp 18001
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_389
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_390
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_391
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_392
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_393
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_394
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_395
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_396
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_397
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_398
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_399
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_400
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_401
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_402
timestamp 18001
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_403
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_404
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_405
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_406
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_407
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_408
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_409
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_410
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_411
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_412
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_413
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_414
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_415
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_416
timestamp 18001
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_417
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_418
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_419
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_420
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_421
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_422
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_423
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_424
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_425
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_426
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_427
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_428
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_429
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_430
timestamp 18001
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_431
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_432
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_433
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_434
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_435
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_436
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_437
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_438
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_439
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_440
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_441
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_442
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_443
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_444
timestamp 18001
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_445
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_446
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_447
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_448
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_449
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_450
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_451
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_452
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_453
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_454
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_455
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_456
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_457
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_458
timestamp 18001
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_459
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_460
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_461
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_462
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_463
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_464
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_465
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_466
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_467
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_468
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_469
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_470
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_471
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_472
timestamp 18001
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_473
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_474
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_475
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_476
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_477
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_478
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_479
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_480
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_481
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_482
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_483
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_484
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_485
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_486
timestamp 18001
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_487
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_488
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_489
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_490
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_491
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_492
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_493
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_494
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_495
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_496
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_497
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_498
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_499
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_500
timestamp 18001
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_501
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_502
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_503
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_504
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_505
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_506
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_507
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_508
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_509
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_510
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_511
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_512
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_513
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_514
timestamp 18001
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_515
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_516
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_517
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_518
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_519
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_520
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_521
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_522
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_523
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_524
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_525
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_526
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_527
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_528
timestamp 18001
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_529
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_530
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_531
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_532
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_533
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_534
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_535
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_536
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_537
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_538
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_539
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_540
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_541
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_542
timestamp 18001
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_543
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_544
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_545
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_546
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_547
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_548
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_549
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_550
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_551
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_552
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_553
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_554
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_555
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_556
timestamp 18001
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_557
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_558
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_559
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_560
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_561
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_562
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_563
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_564
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_565
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_566
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_567
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_568
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_569
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_570
timestamp 18001
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_571
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_572
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_573
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_574
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_575
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_576
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_577
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_578
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_579
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_580
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_581
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_582
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_583
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_584
timestamp 18001
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_585
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_586
timestamp 18001
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_587
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_588
timestamp 18001
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_589
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_590
timestamp 18001
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_591
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_592
timestamp 18001
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_593
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_594
timestamp 18001
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_595
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_596
timestamp 18001
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_597
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_598
timestamp 18001
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  team_02_88
timestamp 18001
transform -1 0 28060 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_89
timestamp 18001
transform -1 0 24196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_90
timestamp 18001
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_91
timestamp 18001
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_92
timestamp 18001
transform -1 0 1656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_93
timestamp 18001
transform 1 0 38272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_94
timestamp 18001
transform 1 0 38272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_95
timestamp 18001
transform -1 0 1656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_96
timestamp 18001
transform -1 0 37076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_97
timestamp 18001
transform -1 0 35144 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_98
timestamp 18001
transform -1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_99
timestamp 18001
transform 1 0 37996 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_100
timestamp 18001
transform -1 0 29992 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_101
timestamp 18001
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_102
timestamp 18001
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_103
timestamp 18001
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_104
timestamp 18001
transform 1 0 38272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_105
timestamp 18001
transform 1 0 38272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_106
timestamp 18001
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_107
timestamp 18001
transform -1 0 1656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_108
timestamp 18001
transform -1 0 1932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_109
timestamp 18001
transform -1 0 35788 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_110
timestamp 18001
transform 1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_111
timestamp 18001
transform -1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_112
timestamp 18001
transform -1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_113
timestamp 18001
transform 1 0 38272 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_114
timestamp 18001
transform 1 0 37996 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_115
timestamp 18001
transform -1 0 36432 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_116
timestamp 18001
transform -1 0 34500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_117
timestamp 18001
transform -1 0 1656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_118
timestamp 18001
transform 1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_119
timestamp 18001
transform -1 0 3588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_120
timestamp 18001
transform -1 0 29348 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_121
timestamp 18001
transform 1 0 37720 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_126
timestamp 18001
transform -1 0 38548 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_127
timestamp 18001
transform -1 0 38548 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_128
timestamp 18001
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_129
timestamp 18001
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_130
timestamp 18001
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_131
timestamp 18001
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_132
timestamp 18001
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_133
timestamp 18001
transform -1 0 38548 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_134
timestamp 18001
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_135
timestamp 18001
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_136
timestamp 18001
transform 1 0 31648 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_137
timestamp 18001
transform 1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_138
timestamp 18001
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_139
timestamp 18001
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_140
timestamp 18001
transform -1 0 38548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_141
timestamp 18001
transform 1 0 28428 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_142
timestamp 18001
transform 1 0 30360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_143
timestamp 18001
transform -1 0 38548 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_144
timestamp 18001
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_145
timestamp 18001
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_146
timestamp 18001
transform 1 0 31004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_147
timestamp 18001
transform 1 0 32936 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_148
timestamp 18001
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_149
timestamp 18001
transform -1 0 38548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_150
timestamp 18001
transform 1 0 29072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_151
timestamp 18001
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  team_02_152
timestamp 18001
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire23
timestamp 18001
transform 1 0 2852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire24
timestamp 18001
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire25
timestamp 18001
transform 1 0 36248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire30
timestamp 18001
transform -1 0 13156 0 -1 21760
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 en
port 1 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio_in[0]
port 2 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 gpio_in[10]
port 3 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 gpio_in[11]
port 4 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 gpio_in[12]
port 5 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 gpio_in[13]
port 6 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 gpio_in[14]
port 7 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 gpio_in[15]
port 8 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 gpio_in[16]
port 9 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpio_in[17]
port 10 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 gpio_in[18]
port 11 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpio_in[19]
port 12 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpio_in[1]
port 13 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpio_in[20]
port 14 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpio_in[21]
port 15 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 gpio_in[22]
port 16 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gpio_in[23]
port 17 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 gpio_in[24]
port 18 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 gpio_in[25]
port 19 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 gpio_in[26]
port 20 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 gpio_in[27]
port 21 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpio_in[28]
port 22 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 gpio_in[29]
port 23 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gpio_in[2]
port 24 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpio_in[30]
port 25 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gpio_in[31]
port 26 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 gpio_in[32]
port 27 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 gpio_in[33]
port 28 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpio_in[3]
port 29 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpio_in[4]
port 30 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 gpio_in[5]
port 31 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpio_in[6]
port 32 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpio_in[7]
port 33 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 gpio_in[8]
port 34 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 gpio_in[9]
port 35 nsew signal input
flabel metal3 s 39200 14968 40000 15088 0 FreeSans 480 0 0 0 gpio_oeb[0]
port 36 nsew signal output
flabel metal3 s 39200 31288 40000 31408 0 FreeSans 480 0 0 0 gpio_oeb[10]
port 37 nsew signal output
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpio_oeb[11]
port 38 nsew signal output
flabel metal2 s 36726 39200 36782 40000 0 FreeSans 224 90 0 0 gpio_oeb[12]
port 39 nsew signal output
flabel metal2 s 34794 39200 34850 40000 0 FreeSans 224 90 0 0 gpio_oeb[13]
port 40 nsew signal output
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 gpio_oeb[14]
port 41 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 gpio_oeb[15]
port 42 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 gpio_oeb[16]
port 43 nsew signal output
flabel metal3 s 39200 36048 40000 36168 0 FreeSans 480 0 0 0 gpio_oeb[17]
port 44 nsew signal output
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 gpio_oeb[18]
port 45 nsew signal output
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 gpio_oeb[19]
port 46 nsew signal output
flabel metal3 s 39200 36728 40000 36848 0 FreeSans 480 0 0 0 gpio_oeb[1]
port 47 nsew signal output
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 gpio_oeb[20]
port 48 nsew signal output
flabel metal2 s 5170 39200 5226 40000 0 FreeSans 224 90 0 0 gpio_oeb[21]
port 49 nsew signal output
flabel metal2 s 27066 39200 27122 40000 0 FreeSans 224 90 0 0 gpio_oeb[22]
port 50 nsew signal output
flabel metal2 s 33506 39200 33562 40000 0 FreeSans 224 90 0 0 gpio_oeb[23]
port 51 nsew signal output
flabel metal3 s 39200 2048 40000 2168 0 FreeSans 480 0 0 0 gpio_oeb[24]
port 52 nsew signal output
flabel metal2 s 28354 39200 28410 40000 0 FreeSans 224 90 0 0 gpio_oeb[25]
port 53 nsew signal output
flabel metal2 s 30286 39200 30342 40000 0 FreeSans 224 90 0 0 gpio_oeb[26]
port 54 nsew signal output
flabel metal3 s 39200 34688 40000 34808 0 FreeSans 480 0 0 0 gpio_oeb[27]
port 55 nsew signal output
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 gpio_oeb[28]
port 56 nsew signal output
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 gpio_oeb[29]
port 57 nsew signal output
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 gpio_oeb[2]
port 58 nsew signal output
flabel metal2 s 30930 39200 30986 40000 0 FreeSans 224 90 0 0 gpio_oeb[30]
port 59 nsew signal output
flabel metal2 s 32862 39200 32918 40000 0 FreeSans 224 90 0 0 gpio_oeb[31]
port 60 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 gpio_oeb[32]
port 61 nsew signal output
flabel metal3 s 39200 2728 40000 2848 0 FreeSans 480 0 0 0 gpio_oeb[33]
port 62 nsew signal output
flabel metal2 s 27710 39200 27766 40000 0 FreeSans 224 90 0 0 gpio_oeb[3]
port 63 nsew signal output
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 gpio_oeb[4]
port 64 nsew signal output
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 gpio_oeb[5]
port 65 nsew signal output
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 gpio_oeb[6]
port 66 nsew signal output
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 gpio_oeb[7]
port 67 nsew signal output
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 gpio_oeb[8]
port 68 nsew signal output
flabel metal3 s 39200 39448 40000 39568 0 FreeSans 480 0 0 0 gpio_oeb[9]
port 69 nsew signal output
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 gpio_out[0]
port 70 nsew signal output
flabel metal3 s 39200 27208 40000 27328 0 FreeSans 480 0 0 0 gpio_out[10]
port 71 nsew signal output
flabel metal2 s 23846 39200 23902 40000 0 FreeSans 224 90 0 0 gpio_out[11]
port 72 nsew signal output
flabel metal2 s 25778 39200 25834 40000 0 FreeSans 224 90 0 0 gpio_out[12]
port 73 nsew signal output
flabel metal2 s 26422 39200 26478 40000 0 FreeSans 224 90 0 0 gpio_out[13]
port 74 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 gpio_out[14]
port 75 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 gpio_out[15]
port 76 nsew signal output
flabel metal3 s 39200 35368 40000 35488 0 FreeSans 480 0 0 0 gpio_out[16]
port 77 nsew signal output
flabel metal3 s 39200 34008 40000 34128 0 FreeSans 480 0 0 0 gpio_out[17]
port 78 nsew signal output
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 gpio_out[18]
port 79 nsew signal output
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 gpio_out[19]
port 80 nsew signal output
flabel metal3 s 39200 38088 40000 38208 0 FreeSans 480 0 0 0 gpio_out[1]
port 81 nsew signal output
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 gpio_out[20]
port 82 nsew signal output
flabel metal2 s 35438 39200 35494 40000 0 FreeSans 224 90 0 0 gpio_out[21]
port 83 nsew signal output
flabel metal3 s 39200 33328 40000 33448 0 FreeSans 480 0 0 0 gpio_out[22]
port 84 nsew signal output
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 gpio_out[23]
port 85 nsew signal output
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 gpio_out[24]
port 86 nsew signal output
flabel metal3 s 39200 30608 40000 30728 0 FreeSans 480 0 0 0 gpio_out[25]
port 87 nsew signal output
flabel metal3 s 39200 37408 40000 37528 0 FreeSans 480 0 0 0 gpio_out[26]
port 88 nsew signal output
flabel metal2 s 36082 39200 36138 40000 0 FreeSans 224 90 0 0 gpio_out[27]
port 89 nsew signal output
flabel metal2 s 34150 39200 34206 40000 0 FreeSans 224 90 0 0 gpio_out[28]
port 90 nsew signal output
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 gpio_out[29]
port 91 nsew signal output
flabel metal2 s 29642 39200 29698 40000 0 FreeSans 224 90 0 0 gpio_out[2]
port 92 nsew signal output
flabel metal3 s 39200 3408 40000 3528 0 FreeSans 480 0 0 0 gpio_out[30]
port 93 nsew signal output
flabel metal2 s 3238 39200 3294 40000 0 FreeSans 224 90 0 0 gpio_out[31]
port 94 nsew signal output
flabel metal2 s 28998 39200 29054 40000 0 FreeSans 224 90 0 0 gpio_out[32]
port 95 nsew signal output
flabel metal3 s 39200 38768 40000 38888 0 FreeSans 480 0 0 0 gpio_out[33]
port 96 nsew signal output
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 gpio_out[3]
port 97 nsew signal output
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 gpio_out[4]
port 98 nsew signal output
flabel metal2 s 32218 39200 32274 40000 0 FreeSans 224 90 0 0 gpio_out[5]
port 99 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 gpio_out[6]
port 100 nsew signal output
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 gpio_out[7]
port 101 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 gpio_out[8]
port 102 nsew signal output
flabel metal3 s 39200 7488 40000 7608 0 FreeSans 480 0 0 0 gpio_out[9]
port 103 nsew signal output
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 nrst
port 104 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 105 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 105 nsew power bidirectional
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 vssd1
port 106 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 vssd1
port 106 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 16376 13362 16376 13362 0 _0000_
rlabel metal1 17802 15062 17802 15062 0 _0001_
rlabel metal1 2852 10710 2852 10710 0 _0002_
rlabel metal1 6164 16014 6164 16014 0 _0003_
rlabel metal2 6578 17884 6578 17884 0 _0004_
rlabel metal1 2116 17850 2116 17850 0 _0005_
rlabel metal1 1748 19278 1748 19278 0 _0006_
rlabel metal2 2806 20638 2806 20638 0 _0007_
rlabel metal2 5382 20706 5382 20706 0 _0008_
rlabel metal1 5336 19210 5336 19210 0 _0009_
rlabel metal1 4002 11186 4002 11186 0 _0010_
rlabel metal1 6256 11186 6256 11186 0 _0011_
rlabel metal1 6118 14042 6118 14042 0 _0012_
rlabel metal1 4738 12954 4738 12954 0 _0013_
rlabel metal2 2806 13124 2806 13124 0 _0014_
rlabel metal2 3358 13974 3358 13974 0 _0015_
rlabel metal2 2254 14756 2254 14756 0 _0016_
rlabel metal2 1702 16320 1702 16320 0 _0017_
rlabel metal1 3450 15980 3450 15980 0 _0018_
rlabel metal1 5888 14858 5888 14858 0 _0019_
rlabel metal2 10994 34850 10994 34850 0 _0020_
rlabel metal1 14444 31654 14444 31654 0 _0021_
rlabel metal2 15778 30124 15778 30124 0 _0022_
rlabel metal1 18032 30158 18032 30158 0 _0023_
rlabel metal1 13432 30158 13432 30158 0 _0024_
rlabel metal1 13708 29070 13708 29070 0 _0025_
rlabel metal2 11638 34136 11638 34136 0 _0026_
rlabel metal2 12466 35054 12466 35054 0 _0027_
rlabel metal2 15502 34782 15502 34782 0 _0028_
rlabel metal2 16238 34204 16238 34204 0 _0029_
rlabel metal2 18906 34782 18906 34782 0 _0030_
rlabel metal1 19918 31858 19918 31858 0 _0031_
rlabel metal2 20746 32028 20746 32028 0 _0032_
rlabel metal2 16974 32606 16974 32606 0 _0033_
rlabel metal2 14674 32606 14674 32606 0 _0034_
rlabel metal1 11316 5542 11316 5542 0 _0035_
rlabel metal2 6946 13022 6946 13022 0 _0036_
rlabel metal1 13110 4250 13110 4250 0 _0037_
rlabel metal2 11822 3230 11822 3230 0 _0038_
rlabel metal1 10810 2958 10810 2958 0 _0039_
rlabel metal2 9246 3332 9246 3332 0 _0040_
rlabel metal1 7268 2482 7268 2482 0 _0041_
rlabel metal2 7222 6698 7222 6698 0 _0042_
rlabel metal1 8648 6426 8648 6426 0 _0043_
rlabel metal2 6854 4828 6854 4828 0 _0044_
rlabel metal1 5244 5134 5244 5134 0 _0045_
rlabel metal2 5658 3740 5658 3740 0 _0046_
rlabel metal1 6716 11322 6716 11322 0 _0047_
rlabel metal1 4002 2958 4002 2958 0 _0048_
rlabel metal1 3680 3706 3680 3706 0 _0049_
rlabel metal1 2162 5576 2162 5576 0 _0050_
rlabel metal1 2024 6222 2024 6222 0 _0051_
rlabel metal1 5204 6970 5204 6970 0 _0052_
rlabel metal2 2898 7854 2898 7854 0 _0053_
rlabel metal2 5290 9724 5290 9724 0 _0054_
rlabel metal2 5382 8024 5382 8024 0 _0055_
rlabel metal2 8326 8296 8326 8296 0 _0056_
rlabel metal2 6670 9180 6670 9180 0 _0057_
rlabel metal1 8280 11798 8280 11798 0 _0058_
rlabel metal1 6854 10744 6854 10744 0 _0059_
rlabel metal2 8786 10404 8786 10404 0 _0060_
rlabel metal1 9568 9146 9568 9146 0 _0061_
rlabel metal1 9798 8058 9798 8058 0 _0062_
rlabel metal2 10350 7650 10350 7650 0 _0063_
rlabel metal1 12558 6154 12558 6154 0 _0064_
rlabel metal1 14398 5746 14398 5746 0 _0065_
rlabel metal1 15134 23528 15134 23528 0 _0066_
rlabel via1 6854 15997 6854 15997 0 _0067_
rlabel metal1 9798 26554 9798 26554 0 _0068_
rlabel metal2 8326 26724 8326 26724 0 _0069_
rlabel metal1 7084 25466 7084 25466 0 _0070_
rlabel metal2 5658 26078 5658 26078 0 _0071_
rlabel metal1 5244 24718 5244 24718 0 _0072_
rlabel via1 5927 22202 5927 22202 0 _0073_
rlabel metal2 7038 22814 7038 22814 0 _0074_
rlabel metal1 4554 21658 4554 21658 0 _0075_
rlabel metal2 2346 22814 2346 22814 0 _0076_
rlabel metal1 1932 23290 1932 23290 0 _0077_
rlabel metal1 9062 16626 9062 16626 0 _0078_
rlabel metal2 1794 24956 1794 24956 0 _0079_
rlabel metal2 4094 25500 4094 25500 0 _0080_
rlabel metal2 4002 26724 4002 26724 0 _0081_
rlabel metal1 1840 26894 1840 26894 0 _0082_
rlabel metal1 2162 28152 2162 28152 0 _0083_
rlabel metal1 3450 28730 3450 28730 0 _0084_
rlabel metal2 4738 29376 4738 29376 0 _0085_
rlabel metal1 4186 28730 4186 28730 0 _0086_
rlabel metal1 7682 27982 7682 27982 0 _0087_
rlabel metal1 7268 29206 7268 29206 0 _0088_
rlabel metal2 9154 17714 9154 17714 0 _0089_
rlabel metal2 6946 18972 6946 18972 0 _0090_
rlabel metal2 6670 20060 6670 20060 0 _0091_
rlabel metal2 9430 20808 9430 20808 0 _0092_
rlabel metal1 9338 22066 9338 22066 0 _0093_
rlabel metal1 9154 22746 9154 22746 0 _0094_
rlabel metal2 10534 24412 10534 24412 0 _0095_
rlabel metal1 10488 25806 10488 25806 0 _0096_
rlabel metal1 23092 14586 23092 14586 0 _0097_
rlabel metal2 25530 14756 25530 14756 0 _0098_
rlabel metal2 22126 13668 22126 13668 0 _0099_
rlabel metal1 23782 31790 23782 31790 0 _0100_
rlabel metal1 23874 30294 23874 30294 0 _0101_
rlabel metal1 25760 27914 25760 27914 0 _0102_
rlabel metal1 24012 26554 24012 26554 0 _0103_
rlabel metal2 27922 26622 27922 26622 0 _0104_
rlabel metal1 26404 27506 26404 27506 0 _0105_
rlabel metal1 27232 28186 27232 28186 0 _0106_
rlabel metal1 26496 29818 26496 29818 0 _0107_
rlabel metal1 26358 30804 26358 30804 0 _0108_
rlabel metal2 25622 32674 25622 32674 0 _0109_
rlabel metal1 24978 36346 24978 36346 0 _0110_
rlabel metal2 24610 34782 24610 34782 0 _0111_
rlabel metal1 23092 36346 23092 36346 0 _0112_
rlabel metal2 26266 33218 26266 33218 0 _0113_
rlabel metal1 27416 31926 27416 31926 0 _0114_
rlabel metal1 28980 32334 28980 32334 0 _0115_
rlabel metal1 27646 33626 27646 33626 0 _0116_
rlabel metal1 21344 30362 21344 30362 0 _0117_
rlabel metal2 22494 29274 22494 29274 0 _0118_
rlabel via1 19177 29138 19177 29138 0 _0119_
rlabel metal1 23230 25466 23230 25466 0 _0120_
rlabel metal1 23414 24378 23414 24378 0 _0121_
rlabel metal1 22202 27370 22202 27370 0 _0122_
rlabel via1 22857 28050 22857 28050 0 _0123_
rlabel metal1 20842 29614 20842 29614 0 _0124_
rlabel metal1 22264 31450 22264 31450 0 _0125_
rlabel metal2 18630 16490 18630 16490 0 _0126_
rlabel metal1 21390 15538 21390 15538 0 _0127_
rlabel metal2 19550 16796 19550 16796 0 _0128_
rlabel metal1 21160 14042 21160 14042 0 _0129_
rlabel metal1 19872 12682 19872 12682 0 _0130_
rlabel metal1 19136 11662 19136 11662 0 _0131_
rlabel metal2 20746 10404 20746 10404 0 _0132_
rlabel metal1 20700 9486 20700 9486 0 _0133_
rlabel metal1 21022 8364 21022 8364 0 _0134_
rlabel metal1 20371 6970 20371 6970 0 _0135_
rlabel metal1 20700 5134 20700 5134 0 _0136_
rlabel metal1 21390 3400 21390 3400 0 _0137_
rlabel metal1 22632 3094 22632 3094 0 _0138_
rlabel metal1 24840 3026 24840 3026 0 _0139_
rlabel metal2 9246 29852 9246 29852 0 _0140_
rlabel metal1 10028 28186 10028 28186 0 _0141_
rlabel metal2 11454 29036 11454 29036 0 _0142_
rlabel metal2 10166 30872 10166 30872 0 _0143_
rlabel metal2 12558 32164 12558 32164 0 _0144_
rlabel metal2 10258 32164 10258 32164 0 _0145_
rlabel metal1 10534 34034 10534 34034 0 _0146_
rlabel metal2 9706 33320 9706 33320 0 _0147_
rlabel metal2 6026 33116 6026 33116 0 _0148_
rlabel metal2 9062 30430 9062 30430 0 _0149_
rlabel metal1 7682 31212 7682 31212 0 _0150_
rlabel metal1 5428 32198 5428 32198 0 _0151_
rlabel metal1 3772 30906 3772 30906 0 _0152_
rlabel metal2 2530 31926 2530 31926 0 _0153_
rlabel metal1 3864 32810 3864 32810 0 _0154_
rlabel metal2 2530 33694 2530 33694 0 _0155_
rlabel metal2 2898 34884 2898 34884 0 _0156_
rlabel metal1 4416 34986 4416 34986 0 _0157_
rlabel metal2 5198 36516 5198 36516 0 _0158_
rlabel metal2 7222 36516 7222 36516 0 _0159_
rlabel metal1 7360 35598 7360 35598 0 _0160_
rlabel metal2 8050 35428 8050 35428 0 _0161_
rlabel metal2 13018 28186 13018 28186 0 _0162_
rlabel metal1 13018 27608 13018 27608 0 _0163_
rlabel metal2 15502 28186 15502 28186 0 _0164_
rlabel metal1 16934 27642 16934 27642 0 _0165_
rlabel metal2 17618 28322 17618 28322 0 _0166_
rlabel metal1 15587 22202 15587 22202 0 _0167_
rlabel metal2 23874 20910 23874 20910 0 _0168_
rlabel metal2 28106 20536 28106 20536 0 _0169_
rlabel metal1 29670 19278 29670 19278 0 _0170_
rlabel metal2 28106 16422 28106 16422 0 _0171_
rlabel metal2 30498 16218 30498 16218 0 _0172_
rlabel metal1 32890 16626 32890 16626 0 _0173_
rlabel metal1 34730 17238 34730 17238 0 _0174_
rlabel metal2 35834 17884 35834 17884 0 _0175_
rlabel metal2 25254 15810 25254 15810 0 _0176_
rlabel metal1 21804 17306 21804 17306 0 _0177_
rlabel metal1 22816 16218 22816 16218 0 _0178_
rlabel metal2 27462 35360 27462 35360 0 _0179_
rlabel metal2 16974 17816 16974 17816 0 _0180_
rlabel metal2 19826 18564 19826 18564 0 _0181_
rlabel metal1 19550 18802 19550 18802 0 _0182_
rlabel metal2 14398 8092 14398 8092 0 _0183_
rlabel metal1 14766 7480 14766 7480 0 _0184_
rlabel metal2 16974 7582 16974 7582 0 _0185_
rlabel metal2 17250 8092 17250 8092 0 _0186_
rlabel metal2 17986 9316 17986 9316 0 _0187_
rlabel metal2 18170 10404 18170 10404 0 _0188_
rlabel metal2 17434 11492 17434 11492 0 _0189_
rlabel metal1 17250 12104 17250 12104 0 _0190_
rlabel metal1 15548 12410 15548 12410 0 _0191_
rlabel metal1 13202 11798 13202 11798 0 _0192_
rlabel metal1 12374 11220 12374 11220 0 _0193_
rlabel metal1 11960 9690 11960 9690 0 _0194_
rlabel metal2 13202 9452 13202 9452 0 _0195_
rlabel metal2 12834 8942 12834 8942 0 _0196_
rlabel metal2 14398 10914 14398 10914 0 _0197_
rlabel metal1 15410 13498 15410 13498 0 _0198_
rlabel metal2 14398 15708 14398 15708 0 _0199_
rlabel metal1 11224 15130 11224 15130 0 _0200_
rlabel metal1 9338 16150 9338 16150 0 _0201_
rlabel metal2 9614 14756 9614 14756 0 _0202_
rlabel metal1 8917 13702 8917 13702 0 _0203_
rlabel metal2 9706 13022 9706 13022 0 _0204_
rlabel metal1 11546 13192 11546 13192 0 _0205_
rlabel metal2 13018 14722 13018 14722 0 _0206_
rlabel metal2 13938 20196 13938 20196 0 _0207_
rlabel metal1 12282 19278 12282 19278 0 _0208_
rlabel metal2 9798 19482 9798 19482 0 _0209_
rlabel metal1 9752 18394 9752 18394 0 _0210_
rlabel metal1 9890 17306 9890 17306 0 _0211_
rlabel metal1 11362 17306 11362 17306 0 _0212_
rlabel metal1 14398 17544 14398 17544 0 _0213_
rlabel metal1 15180 18326 15180 18326 0 _0214_
rlabel metal1 15272 19278 15272 19278 0 _0215_
rlabel metal1 16238 19890 16238 19890 0 _0216_
rlabel metal1 18170 21658 18170 21658 0 _0217_
rlabel metal1 14628 21114 14628 21114 0 _0218_
rlabel metal1 12834 21658 12834 21658 0 _0219_
rlabel metal2 11822 21794 11822 21794 0 _0220_
rlabel metal2 10718 21148 10718 21148 0 _0221_
rlabel metal2 19826 20196 19826 20196 0 _0222_
rlabel metal1 18952 20570 18952 20570 0 _0223_
rlabel metal1 18078 18326 18078 18326 0 _0224_
rlabel metal1 17388 12886 17388 12886 0 _0225_
rlabel metal2 27738 6052 27738 6052 0 _0226_
rlabel metal2 26818 6086 26818 6086 0 _0227_
rlabel metal2 27278 6630 27278 6630 0 _0228_
rlabel metal1 28382 6188 28382 6188 0 _0229_
rlabel metal2 29302 6596 29302 6596 0 _0230_
rlabel metal1 29716 6630 29716 6630 0 _0231_
rlabel metal1 30038 6290 30038 6290 0 _0232_
rlabel metal1 31970 6290 31970 6290 0 _0233_
rlabel metal1 32338 6222 32338 6222 0 _0234_
rlabel metal1 32246 6358 32246 6358 0 _0235_
rlabel metal2 32062 5882 32062 5882 0 _0236_
rlabel metal2 32338 6290 32338 6290 0 _0237_
rlabel metal1 29992 6698 29992 6698 0 _0238_
rlabel metal2 30406 7378 30406 7378 0 _0239_
rlabel metal2 27830 7412 27830 7412 0 _0240_
rlabel metal2 27370 7684 27370 7684 0 _0241_
rlabel metal1 26910 7514 26910 7514 0 _0242_
rlabel metal1 27140 8058 27140 8058 0 _0243_
rlabel metal1 28198 7922 28198 7922 0 _0244_
rlabel metal2 28290 8228 28290 8228 0 _0245_
rlabel metal1 28612 8534 28612 8534 0 _0246_
rlabel metal1 29302 7922 29302 7922 0 _0247_
rlabel metal1 30728 7854 30728 7854 0 _0248_
rlabel metal1 31234 6256 31234 6256 0 _0249_
rlabel metal1 31464 7854 31464 7854 0 _0250_
rlabel metal2 31142 8262 31142 8262 0 _0251_
rlabel metal2 30130 8466 30130 8466 0 _0252_
rlabel metal2 28014 8738 28014 8738 0 _0253_
rlabel via2 25254 8483 25254 8483 0 _0254_
rlabel metal1 25530 8602 25530 8602 0 _0255_
rlabel metal1 26220 9146 26220 9146 0 _0256_
rlabel metal1 27600 8942 27600 8942 0 _0257_
rlabel metal2 28198 9350 28198 9350 0 _0258_
rlabel metal1 28796 8466 28796 8466 0 _0259_
rlabel metal2 29762 8772 29762 8772 0 _0260_
rlabel metal1 30590 9044 30590 9044 0 _0261_
rlabel metal1 30774 8908 30774 8908 0 _0262_
rlabel metal2 31050 9316 31050 9316 0 _0263_
rlabel metal2 28382 9350 28382 9350 0 _0264_
rlabel metal2 28474 9826 28474 9826 0 _0265_
rlabel metal2 27186 10438 27186 10438 0 _0266_
rlabel metal2 23184 9554 23184 9554 0 _0267_
rlabel metal1 25898 9554 25898 9554 0 _0268_
rlabel metal1 26128 10710 26128 10710 0 _0269_
rlabel metal1 26956 10574 26956 10574 0 _0270_
rlabel metal2 28290 10234 28290 10234 0 _0271_
rlabel metal1 28888 10166 28888 10166 0 _0272_
rlabel metal1 28934 10234 28934 10234 0 _0273_
rlabel metal2 29210 10914 29210 10914 0 _0274_
rlabel metal1 27876 10166 27876 10166 0 _0275_
rlabel via1 28566 10710 28566 10710 0 _0276_
rlabel metal1 30176 10574 30176 10574 0 _0277_
rlabel metal1 29578 9690 29578 9690 0 _0278_
rlabel metal2 30130 10438 30130 10438 0 _0279_
rlabel metal1 31418 9588 31418 9588 0 _0280_
rlabel metal1 30958 9520 30958 9520 0 _0281_
rlabel metal1 31418 9928 31418 9928 0 _0282_
rlabel metal2 31786 8092 31786 8092 0 _0283_
rlabel metal1 32108 7310 32108 7310 0 _0284_
rlabel metal2 32430 6460 32430 6460 0 _0285_
rlabel metal1 32936 6222 32936 6222 0 _0286_
rlabel metal2 33902 5372 33902 5372 0 _0287_
rlabel metal2 34730 4182 34730 4182 0 _0288_
rlabel metal1 33672 4590 33672 4590 0 _0289_
rlabel metal1 34454 5168 34454 5168 0 _0290_
rlabel metal2 35374 5950 35374 5950 0 _0291_
rlabel metal2 35098 5508 35098 5508 0 _0292_
rlabel metal1 31188 11662 31188 11662 0 _0293_
rlabel metal1 32568 10574 32568 10574 0 _0294_
rlabel metal1 33626 10778 33626 10778 0 _0295_
rlabel metal1 34408 7922 34408 7922 0 _0296_
rlabel metal2 35282 8704 35282 8704 0 _0297_
rlabel metal2 35834 7072 35834 7072 0 _0298_
rlabel metal1 35512 6766 35512 6766 0 _0299_
rlabel metal1 35146 6290 35146 6290 0 _0300_
rlabel metal1 35466 11050 35466 11050 0 _0301_
rlabel metal2 34546 6137 34546 6137 0 _0302_
rlabel metal2 34178 4998 34178 4998 0 _0303_
rlabel metal2 34730 5508 34730 5508 0 _0304_
rlabel metal2 34454 6052 34454 6052 0 _0305_
rlabel metal1 34684 5882 34684 5882 0 _0306_
rlabel metal2 33810 7344 33810 7344 0 _0307_
rlabel metal1 33672 5338 33672 5338 0 _0308_
rlabel metal1 34385 6766 34385 6766 0 _0309_
rlabel metal1 32982 5882 32982 5882 0 _0310_
rlabel metal1 33534 6698 33534 6698 0 _0311_
rlabel metal1 34868 7854 34868 7854 0 _0312_
rlabel metal2 33534 7548 33534 7548 0 _0313_
rlabel metal1 32752 7378 32752 7378 0 _0314_
rlabel metal1 33534 11016 33534 11016 0 _0315_
rlabel metal2 32982 8908 32982 8908 0 _0316_
rlabel metal1 33350 7344 33350 7344 0 _0317_
rlabel metal2 33166 7106 33166 7106 0 _0318_
rlabel metal2 31878 8772 31878 8772 0 _0319_
rlabel metal2 32706 9350 32706 9350 0 _0320_
rlabel metal1 32890 9554 32890 9554 0 _0321_
rlabel metal1 31809 10030 31809 10030 0 _0322_
rlabel metal1 32154 10064 32154 10064 0 _0323_
rlabel metal2 32154 9724 32154 9724 0 _0324_
rlabel metal2 30774 10234 30774 10234 0 _0325_
rlabel metal1 30912 10234 30912 10234 0 _0326_
rlabel metal1 31142 12750 31142 12750 0 _0327_
rlabel metal2 30866 11356 30866 11356 0 _0328_
rlabel metal2 30130 11050 30130 11050 0 _0329_
rlabel metal2 30682 10812 30682 10812 0 _0330_
rlabel metal1 26496 11662 26496 11662 0 _0331_
rlabel metal1 23966 10540 23966 10540 0 _0332_
rlabel metal2 25990 11526 25990 11526 0 _0333_
rlabel metal1 27278 11696 27278 11696 0 _0334_
rlabel metal2 28290 11356 28290 11356 0 _0335_
rlabel metal1 27738 10506 27738 10506 0 _0336_
rlabel metal1 28014 11254 28014 11254 0 _0337_
rlabel metal2 30222 11220 30222 11220 0 _0338_
rlabel metal2 30498 10812 30498 10812 0 _0339_
rlabel metal2 32338 9996 32338 9996 0 _0340_
rlabel metal2 32430 9860 32430 9860 0 _0341_
rlabel metal1 33258 9588 33258 9588 0 _0342_
rlabel metal2 33442 8364 33442 8364 0 _0343_
rlabel metal2 33442 6970 33442 6970 0 _0344_
rlabel metal1 35006 6732 35006 6732 0 _0345_
rlabel via1 34804 6290 34804 6290 0 _0346_
rlabel metal1 35420 6290 35420 6290 0 _0347_
rlabel metal1 35972 6290 35972 6290 0 _0348_
rlabel metal2 35650 6086 35650 6086 0 _0349_
rlabel metal2 36570 7684 36570 7684 0 _0350_
rlabel metal1 36294 6426 36294 6426 0 _0351_
rlabel metal1 35144 10778 35144 10778 0 _0352_
rlabel metal1 35466 11764 35466 11764 0 _0353_
rlabel metal1 34822 14348 34822 14348 0 _0354_
rlabel metal1 34684 14586 34684 14586 0 _0355_
rlabel metal1 35834 11152 35834 11152 0 _0356_
rlabel metal2 36478 9962 36478 9962 0 _0357_
rlabel metal2 27094 14178 27094 14178 0 _0358_
rlabel metal1 26864 13158 26864 13158 0 _0359_
rlabel via1 26826 12138 26826 12138 0 _0360_
rlabel metal1 30774 12614 30774 12614 0 _0361_
rlabel metal1 28244 13158 28244 13158 0 _0362_
rlabel metal2 29854 14484 29854 14484 0 _0363_
rlabel metal1 29854 14042 29854 14042 0 _0364_
rlabel metal2 31050 14416 31050 14416 0 _0365_
rlabel metal2 30682 13362 30682 13362 0 _0366_
rlabel metal1 32024 12070 32024 12070 0 _0367_
rlabel metal2 31602 13260 31602 13260 0 _0368_
rlabel metal1 33212 13974 33212 13974 0 _0369_
rlabel metal1 33166 12886 33166 12886 0 _0370_
rlabel metal1 33580 11526 33580 11526 0 _0371_
rlabel metal1 36264 9622 36264 9622 0 _0372_
rlabel metal1 36340 8466 36340 8466 0 _0373_
rlabel metal1 37582 7888 37582 7888 0 _0374_
rlabel metal1 34408 9690 34408 9690 0 _0375_
rlabel metal1 35466 9690 35466 9690 0 _0376_
rlabel metal1 37168 9622 37168 9622 0 _0377_
rlabel metal1 36708 10778 36708 10778 0 _0378_
rlabel metal1 37674 12614 37674 12614 0 _0379_
rlabel metal1 36340 13974 36340 13974 0 _0380_
rlabel metal1 37122 12852 37122 12852 0 _0381_
rlabel metal1 36754 14042 36754 14042 0 _0382_
rlabel metal1 35604 12954 35604 12954 0 _0383_
rlabel metal1 35688 14042 35688 14042 0 _0384_
rlabel metal1 8142 17748 8142 17748 0 _0385_
rlabel metal2 8510 19142 8510 19142 0 _0386_
rlabel metal1 8602 21012 8602 21012 0 _0387_
rlabel metal2 8694 22814 8694 22814 0 _0388_
rlabel metal2 9614 24242 9614 24242 0 _0389_
rlabel metal1 9936 24718 9936 24718 0 _0390_
rlabel metal1 8694 23562 8694 23562 0 _0391_
rlabel metal1 8786 24378 8786 24378 0 _0392_
rlabel metal1 7176 24786 7176 24786 0 _0393_
rlabel metal2 8142 24378 8142 24378 0 _0394_
rlabel metal1 8840 22746 8840 22746 0 _0395_
rlabel metal1 10902 23664 10902 23664 0 _0396_
rlabel metal1 11040 23766 11040 23766 0 _0397_
rlabel metal1 8402 25942 8402 25942 0 _0398_
rlabel metal2 9798 26044 9798 26044 0 _0399_
rlabel metal1 7636 25806 7636 25806 0 _0400_
rlabel metal1 8648 26010 8648 26010 0 _0401_
rlabel metal1 6900 25262 6900 25262 0 _0402_
rlabel metal2 7130 25466 7130 25466 0 _0403_
rlabel metal2 5842 26316 5842 26316 0 _0404_
rlabel metal1 5888 25262 5888 25262 0 _0405_
rlabel metal2 5658 24820 5658 24820 0 _0406_
rlabel metal1 6118 21658 6118 21658 0 _0407_
rlabel metal1 6210 21386 6210 21386 0 _0408_
rlabel metal2 5198 23562 5198 23562 0 _0409_
rlabel metal1 6578 22678 6578 22678 0 _0410_
rlabel metal1 5060 21454 5060 21454 0 _0411_
rlabel metal1 3174 23120 3174 23120 0 _0412_
rlabel metal1 3220 23698 3220 23698 0 _0413_
rlabel metal1 2553 23086 2553 23086 0 _0414_
rlabel metal2 2070 23902 2070 23902 0 _0415_
rlabel metal2 3266 25126 3266 25126 0 _0416_
rlabel metal1 3404 25874 3404 25874 0 _0417_
rlabel metal1 3818 26384 3818 26384 0 _0418_
rlabel metal2 3174 27404 3174 27404 0 _0419_
rlabel metal1 5014 28016 5014 28016 0 _0420_
rlabel metal1 3542 28526 3542 28526 0 _0421_
rlabel metal2 2990 28730 2990 28730 0 _0422_
rlabel metal1 5106 28084 5106 28084 0 _0423_
rlabel metal1 4600 27846 4600 27846 0 _0424_
rlabel metal2 5474 28118 5474 28118 0 _0425_
rlabel metal1 7268 27982 7268 27982 0 _0426_
rlabel metal1 7314 28118 7314 28118 0 _0427_
rlabel metal1 7452 28730 7452 28730 0 _0428_
rlabel metal1 8556 13430 8556 13430 0 _0429_
rlabel metal1 8280 10234 8280 10234 0 _0430_
rlabel metal1 11178 9418 11178 9418 0 _0431_
rlabel metal2 11362 7072 11362 7072 0 _0432_
rlabel metal2 10810 6664 10810 6664 0 _0433_
rlabel metal1 11776 5746 11776 5746 0 _0434_
rlabel metal1 10902 5610 10902 5610 0 _0435_
rlabel metal1 11500 5814 11500 5814 0 _0436_
rlabel metal2 9706 4964 9706 4964 0 _0437_
rlabel metal1 10074 5338 10074 5338 0 _0438_
rlabel metal2 10166 6664 10166 6664 0 _0439_
rlabel metal2 12926 5508 12926 5508 0 _0440_
rlabel metal1 12696 6290 12696 6290 0 _0441_
rlabel metal2 12374 4556 12374 4556 0 _0442_
rlabel metal2 12650 4556 12650 4556 0 _0443_
rlabel metal1 11270 3468 11270 3468 0 _0444_
rlabel metal1 11546 3536 11546 3536 0 _0445_
rlabel metal1 10350 4046 10350 4046 0 _0446_
rlabel metal1 10534 4080 10534 4080 0 _0447_
rlabel metal2 9982 3808 9982 3808 0 _0448_
rlabel metal2 7590 6834 7590 6834 0 _0449_
rlabel metal2 7866 3910 7866 3910 0 _0450_
rlabel metal2 7774 6732 7774 6732 0 _0451_
rlabel metal1 7406 6324 7406 6324 0 _0452_
rlabel metal2 8234 5984 8234 5984 0 _0453_
rlabel metal1 8510 6256 8510 6256 0 _0454_
rlabel metal2 7130 5372 7130 5372 0 _0455_
rlabel metal1 5934 5678 5934 5678 0 _0456_
rlabel metal1 6026 5338 6026 5338 0 _0457_
rlabel metal2 6026 3638 6026 3638 0 _0458_
rlabel metal1 5796 4114 5796 4114 0 _0459_
rlabel metal2 4002 4114 4002 4114 0 _0460_
rlabel metal1 3818 5644 3818 5644 0 _0461_
rlabel metal1 3404 5202 3404 5202 0 _0462_
rlabel metal1 5382 5882 5382 5882 0 _0463_
rlabel metal2 5290 6766 5290 6766 0 _0464_
rlabel metal2 4094 7378 4094 7378 0 _0465_
rlabel metal2 4738 7990 4738 7990 0 _0466_
rlabel metal1 3956 8466 3956 8466 0 _0467_
rlabel metal1 5198 8398 5198 8398 0 _0468_
rlabel metal1 8142 7718 8142 7718 0 _0469_
rlabel metal2 8602 8126 8602 8126 0 _0470_
rlabel metal2 8510 8704 8510 8704 0 _0471_
rlabel metal1 7176 8058 7176 8058 0 _0472_
rlabel metal2 5842 11764 5842 11764 0 _0473_
rlabel metal2 5842 14246 5842 14246 0 _0474_
rlabel metal1 6686 13974 6686 13974 0 _0475_
rlabel metal1 2116 13362 2116 13362 0 _0476_
rlabel metal1 5106 12818 5106 12818 0 _0477_
rlabel metal1 3956 14382 3956 14382 0 _0478_
rlabel metal1 3818 14450 3818 14450 0 _0479_
rlabel metal1 2484 17170 2484 17170 0 _0480_
rlabel metal2 2438 14858 2438 14858 0 _0481_
rlabel metal2 2438 16524 2438 16524 0 _0482_
rlabel metal1 3082 16082 3082 16082 0 _0483_
rlabel metal1 3450 16150 3450 16150 0 _0484_
rlabel metal1 4692 17850 4692 17850 0 _0485_
rlabel metal1 6210 18190 6210 18190 0 _0486_
rlabel metal1 3174 18122 3174 18122 0 _0487_
rlabel metal1 2622 17680 2622 17680 0 _0488_
rlabel metal1 4002 19754 4002 19754 0 _0489_
rlabel metal1 3726 19278 3726 19278 0 _0490_
rlabel metal2 5750 19856 5750 19856 0 _0491_
rlabel metal1 5014 20026 5014 20026 0 _0492_
rlabel metal1 24334 35734 24334 35734 0 _0493_
rlabel metal2 24242 35292 24242 35292 0 _0494_
rlabel metal1 5244 14586 5244 14586 0 _0495_
rlabel metal1 4416 15674 4416 15674 0 _0496_
rlabel metal1 3956 18870 3956 18870 0 _0497_
rlabel metal1 22356 20230 22356 20230 0 _0498_
rlabel metal1 23230 20400 23230 20400 0 _0499_
rlabel metal1 22816 20910 22816 20910 0 _0500_
rlabel metal2 22218 20264 22218 20264 0 _0501_
rlabel metal2 23966 19550 23966 19550 0 _0502_
rlabel metal1 23016 19822 23016 19822 0 _0503_
rlabel metal1 22126 21046 22126 21046 0 _0504_
rlabel metal1 23368 19346 23368 19346 0 _0505_
rlabel metal2 24242 17204 24242 17204 0 _0506_
rlabel metal1 22678 19822 22678 19822 0 _0507_
rlabel metal1 22586 18700 22586 18700 0 _0508_
rlabel metal1 23874 14416 23874 14416 0 _0509_
rlabel metal1 24334 13906 24334 13906 0 _0510_
rlabel metal1 24012 14382 24012 14382 0 _0511_
rlabel metal1 23828 12818 23828 12818 0 _0512_
rlabel metal1 24288 35258 24288 35258 0 _0513_
rlabel metal2 25254 34748 25254 34748 0 _0514_
rlabel metal1 24610 32198 24610 32198 0 _0515_
rlabel metal1 27416 33490 27416 33490 0 _0516_
rlabel metal1 27922 32742 27922 32742 0 _0517_
rlabel metal1 26818 32402 26818 32402 0 _0518_
rlabel metal1 24840 31110 24840 31110 0 _0519_
rlabel metal1 25438 29648 25438 29648 0 _0520_
rlabel metal1 24104 29818 24104 29818 0 _0521_
rlabel metal2 24426 28764 24426 28764 0 _0522_
rlabel metal1 25162 26316 25162 26316 0 _0523_
rlabel metal1 25760 26010 25760 26010 0 _0524_
rlabel metal1 24932 27438 24932 27438 0 _0525_
rlabel metal2 25254 28560 25254 28560 0 _0526_
rlabel metal2 25254 30124 25254 30124 0 _0527_
rlabel metal1 24978 32368 24978 32368 0 _0528_
rlabel metal1 24196 34714 24196 34714 0 _0529_
rlabel metal1 28428 33626 28428 33626 0 _0530_
rlabel metal1 26910 34714 26910 34714 0 _0531_
rlabel metal2 24978 34884 24978 34884 0 _0532_
rlabel metal1 25300 35802 25300 35802 0 _0533_
rlabel metal1 26266 32538 26266 32538 0 _0534_
rlabel viali 27656 31790 27656 31790 0 _0535_
rlabel metal1 26864 31722 26864 31722 0 _0536_
rlabel metal2 27830 32198 27830 32198 0 _0537_
rlabel metal2 27922 33966 27922 33966 0 _0538_
rlabel metal1 28336 31994 28336 31994 0 _0539_
rlabel metal1 28014 33524 28014 33524 0 _0540_
rlabel metal2 15594 25942 15594 25942 0 _0541_
rlabel metal1 16284 24922 16284 24922 0 _0542_
rlabel metal2 14950 25636 14950 25636 0 _0543_
rlabel metal1 15134 24310 15134 24310 0 _0544_
rlabel metal1 14214 26214 14214 26214 0 _0545_
rlabel metal1 15272 24922 15272 24922 0 _0546_
rlabel metal1 15778 25908 15778 25908 0 _0547_
rlabel metal2 14490 26554 14490 26554 0 _0548_
rlabel metal1 12880 24786 12880 24786 0 _0549_
rlabel metal2 15502 26724 15502 26724 0 _0550_
rlabel metal1 15962 26996 15962 26996 0 _0551_
rlabel metal1 15318 26894 15318 26894 0 _0552_
rlabel metal1 20378 27438 20378 27438 0 _0553_
rlabel metal1 18354 26384 18354 26384 0 _0554_
rlabel metal2 13202 26758 13202 26758 0 _0555_
rlabel via1 13307 25262 13307 25262 0 _0556_
rlabel metal2 15594 24412 15594 24412 0 _0557_
rlabel metal1 15594 25874 15594 25874 0 _0558_
rlabel metal1 14260 25262 14260 25262 0 _0559_
rlabel metal1 13892 25466 13892 25466 0 _0560_
rlabel metal2 14122 26588 14122 26588 0 _0561_
rlabel metal1 13110 25160 13110 25160 0 _0562_
rlabel metal2 13938 24310 13938 24310 0 _0563_
rlabel metal1 13386 24922 13386 24922 0 _0564_
rlabel metal1 13110 27030 13110 27030 0 _0565_
rlabel metal1 13820 25874 13820 25874 0 _0566_
rlabel metal1 15134 24106 15134 24106 0 _0567_
rlabel metal1 14674 24276 14674 24276 0 _0568_
rlabel metal1 14214 24378 14214 24378 0 _0569_
rlabel metal1 19458 22644 19458 22644 0 _0570_
rlabel metal1 18906 24752 18906 24752 0 _0571_
rlabel metal1 19504 22746 19504 22746 0 _0572_
rlabel metal2 20654 26044 20654 26044 0 _0573_
rlabel metal1 16468 24174 16468 24174 0 _0574_
rlabel metal1 16146 24208 16146 24208 0 _0575_
rlabel metal1 17894 24242 17894 24242 0 _0576_
rlabel metal1 19458 23698 19458 23698 0 _0577_
rlabel metal2 14398 24038 14398 24038 0 _0578_
rlabel viali 16701 23698 16701 23698 0 _0579_
rlabel metal1 17342 23732 17342 23732 0 _0580_
rlabel via1 18906 24175 18906 24175 0 _0581_
rlabel metal1 20378 23766 20378 23766 0 _0582_
rlabel metal1 20102 26350 20102 26350 0 _0583_
rlabel metal1 20194 25976 20194 25976 0 _0584_
rlabel metal1 20930 25976 20930 25976 0 _0585_
rlabel metal1 19734 25942 19734 25942 0 _0586_
rlabel metal1 18400 27030 18400 27030 0 _0587_
rlabel metal2 18998 25228 18998 25228 0 _0588_
rlabel metal2 22678 23630 22678 23630 0 _0589_
rlabel metal2 20286 24310 20286 24310 0 _0590_
rlabel metal1 20470 22406 20470 22406 0 _0591_
rlabel metal1 20378 26418 20378 26418 0 _0592_
rlabel metal1 20608 21998 20608 21998 0 _0593_
rlabel via1 21663 25126 21663 25126 0 _0594_
rlabel via1 18630 25738 18630 25738 0 _0595_
rlabel metal1 18354 25262 18354 25262 0 _0596_
rlabel metal2 18814 24990 18814 24990 0 _0597_
rlabel metal1 21390 24820 21390 24820 0 _0598_
rlabel metal2 18906 26180 18906 26180 0 _0599_
rlabel metal1 18354 24922 18354 24922 0 _0600_
rlabel metal2 18722 26044 18722 26044 0 _0601_
rlabel metal2 21390 23868 21390 23868 0 _0602_
rlabel metal1 20654 28050 20654 28050 0 _0603_
rlabel metal1 21160 23698 21160 23698 0 _0604_
rlabel metal1 20654 23018 20654 23018 0 _0605_
rlabel metal1 22080 22542 22080 22542 0 _0606_
rlabel metal1 21850 25194 21850 25194 0 _0607_
rlabel metal2 21850 26214 21850 26214 0 _0608_
rlabel metal1 20378 23120 20378 23120 0 _0609_
rlabel via1 21377 21998 21377 21998 0 _0610_
rlabel metal1 19041 23688 19041 23688 0 _0611_
rlabel metal1 19918 23052 19918 23052 0 _0612_
rlabel metal1 20470 25262 20470 25262 0 _0613_
rlabel metal2 19550 25092 19550 25092 0 _0614_
rlabel metal2 18538 24038 18538 24038 0 _0615_
rlabel metal1 20700 24310 20700 24310 0 _0616_
rlabel metal1 18400 25466 18400 25466 0 _0617_
rlabel metal1 21344 25874 21344 25874 0 _0618_
rlabel metal1 20286 25364 20286 25364 0 _0619_
rlabel metal2 19918 25466 19918 25466 0 _0620_
rlabel metal2 21482 26214 21482 26214 0 _0621_
rlabel metal2 21390 27200 21390 27200 0 _0622_
rlabel metal1 21574 24140 21574 24140 0 _0623_
rlabel metal2 20102 27404 20102 27404 0 _0624_
rlabel metal2 20194 25466 20194 25466 0 _0625_
rlabel metal1 21114 24174 21114 24174 0 _0626_
rlabel metal1 21022 27370 21022 27370 0 _0627_
rlabel metal1 20424 27370 20424 27370 0 _0628_
rlabel metal2 20654 27098 20654 27098 0 _0629_
rlabel metal1 21712 27846 21712 27846 0 _0630_
rlabel metal1 20746 29104 20746 29104 0 _0631_
rlabel metal1 21804 24582 21804 24582 0 _0632_
rlabel metal1 22356 21522 22356 21522 0 _0633_
rlabel metal1 21804 21658 21804 21658 0 _0634_
rlabel metal1 21482 30158 21482 30158 0 _0635_
rlabel metal2 21850 22848 21850 22848 0 _0636_
rlabel metal1 21850 29104 21850 29104 0 _0637_
rlabel metal1 22494 29138 22494 29138 0 _0638_
rlabel metal2 19918 23120 19918 23120 0 _0639_
rlabel metal1 19642 24378 19642 24378 0 _0640_
rlabel metal1 19412 29818 19412 29818 0 _0641_
rlabel metal1 20838 27574 20838 27574 0 _0642_
rlabel metal1 21758 25942 21758 25942 0 _0643_
rlabel via1 22034 24701 22034 24701 0 _0644_
rlabel metal1 22540 24922 22540 24922 0 _0645_
rlabel metal2 22678 25466 22678 25466 0 _0646_
rlabel metal2 21850 24854 21850 24854 0 _0647_
rlabel metal1 22586 24174 22586 24174 0 _0648_
rlabel metal2 22402 27778 22402 27778 0 _0649_
rlabel metal1 20608 28186 20608 28186 0 _0650_
rlabel metal2 20378 29750 20378 29750 0 _0651_
rlabel metal1 21620 28186 21620 28186 0 _0652_
rlabel metal1 19550 14960 19550 14960 0 _0653_
rlabel metal1 17802 14926 17802 14926 0 _0654_
rlabel metal1 20562 15912 20562 15912 0 _0655_
rlabel metal2 20286 15606 20286 15606 0 _0656_
rlabel metal1 20897 16218 20897 16218 0 _0657_
rlabel metal1 20010 16218 20010 16218 0 _0658_
rlabel metal2 20562 14246 20562 14246 0 _0659_
rlabel metal1 19872 13294 19872 13294 0 _0660_
rlabel metal1 20762 13974 20762 13974 0 _0661_
rlabel metal2 19918 12988 19918 12988 0 _0662_
rlabel metal1 20608 12818 20608 12818 0 _0663_
rlabel metal1 25070 13226 25070 13226 0 _0664_
rlabel metal2 25254 14008 25254 14008 0 _0665_
rlabel metal1 24610 13328 24610 13328 0 _0666_
rlabel metal2 24886 13566 24886 13566 0 _0667_
rlabel metal1 24104 13226 24104 13226 0 _0668_
rlabel metal2 22034 11900 22034 11900 0 _0669_
rlabel metal1 23046 11594 23046 11594 0 _0670_
rlabel metal1 23506 11866 23506 11866 0 _0671_
rlabel metal2 22310 11152 22310 11152 0 _0672_
rlabel metal2 24978 10812 24978 10812 0 _0673_
rlabel metal1 24702 8330 24702 8330 0 _0674_
rlabel metal1 23552 12614 23552 12614 0 _0675_
rlabel metal1 24104 11526 24104 11526 0 _0676_
rlabel metal2 25070 9452 25070 9452 0 _0677_
rlabel metal1 25622 6358 25622 6358 0 _0678_
rlabel metal1 26128 6426 26128 6426 0 _0679_
rlabel metal1 25898 6800 25898 6800 0 _0680_
rlabel metal1 25024 6766 25024 6766 0 _0681_
rlabel metal2 24426 6528 24426 6528 0 _0682_
rlabel metal1 25070 10030 25070 10030 0 _0683_
rlabel metal1 24794 10132 24794 10132 0 _0684_
rlabel metal2 23690 8670 23690 8670 0 _0685_
rlabel metal1 24150 9690 24150 9690 0 _0686_
rlabel metal1 23828 10778 23828 10778 0 _0687_
rlabel metal1 24012 10710 24012 10710 0 _0688_
rlabel metal2 23230 11356 23230 11356 0 _0689_
rlabel metal1 24564 10030 24564 10030 0 _0690_
rlabel metal2 24702 10268 24702 10268 0 _0691_
rlabel metal1 24702 7412 24702 7412 0 _0692_
rlabel metal2 25530 6732 25530 6732 0 _0693_
rlabel metal1 26818 4658 26818 4658 0 _0694_
rlabel metal1 26220 5678 26220 5678 0 _0695_
rlabel metal1 25438 5712 25438 5712 0 _0696_
rlabel metal1 25116 5678 25116 5678 0 _0697_
rlabel metal1 25530 4794 25530 4794 0 _0698_
rlabel metal1 25254 5270 25254 5270 0 _0699_
rlabel via1 22034 7803 22034 7803 0 _0700_
rlabel via2 24334 3043 24334 3043 0 _0701_
rlabel metal1 25760 3502 25760 3502 0 _0702_
rlabel metal1 24794 4046 24794 4046 0 _0703_
rlabel metal1 22862 4590 22862 4590 0 _0704_
rlabel metal1 23552 5678 23552 5678 0 _0705_
rlabel metal1 25484 4182 25484 4182 0 _0706_
rlabel metal1 24932 10778 24932 10778 0 _0707_
rlabel metal3 24058 9860 24058 9860 0 _0708_
rlabel metal1 24383 7854 24383 7854 0 _0709_
rlabel metal2 21758 8466 21758 8466 0 _0710_
rlabel metal1 22494 7378 22494 7378 0 _0711_
rlabel metal2 24610 7548 24610 7548 0 _0712_
rlabel metal1 24426 7344 24426 7344 0 _0713_
rlabel metal2 22586 6188 22586 6188 0 _0714_
rlabel metal1 24150 5678 24150 5678 0 _0715_
rlabel metal2 25070 4794 25070 4794 0 _0716_
rlabel metal1 24932 3162 24932 3162 0 _0717_
rlabel metal2 24886 3842 24886 3842 0 _0718_
rlabel metal2 21390 7684 21390 7684 0 _0719_
rlabel metal2 22954 8364 22954 8364 0 _0720_
rlabel metal2 25438 4420 25438 4420 0 _0721_
rlabel metal1 24702 6222 24702 6222 0 _0722_
rlabel via2 23690 10251 23690 10251 0 _0723_
rlabel metal1 21206 10132 21206 10132 0 _0724_
rlabel metal1 22816 10438 22816 10438 0 _0725_
rlabel metal1 22862 9554 22862 9554 0 _0726_
rlabel metal2 22218 9758 22218 9758 0 _0727_
rlabel metal1 23138 6426 23138 6426 0 _0728_
rlabel metal1 22724 7786 22724 7786 0 _0729_
rlabel metal1 21873 7990 21873 7990 0 _0730_
rlabel metal1 24058 7888 24058 7888 0 _0731_
rlabel metal1 23046 7412 23046 7412 0 _0732_
rlabel metal1 20930 7412 20930 7412 0 _0733_
rlabel metal1 22586 5678 22586 5678 0 _0734_
rlabel metal1 21896 5542 21896 5542 0 _0735_
rlabel metal2 22402 5508 22402 5508 0 _0736_
rlabel metal1 22494 5236 22494 5236 0 _0737_
rlabel metal2 23874 4318 23874 4318 0 _0738_
rlabel metal1 24564 3706 24564 3706 0 _0739_
rlabel metal1 9798 29036 9798 29036 0 _0740_
rlabel metal1 11408 29750 11408 29750 0 _0741_
rlabel metal1 11178 30090 11178 30090 0 _0742_
rlabel metal2 12466 31620 12466 31620 0 _0743_
rlabel metal1 10488 31926 10488 31926 0 _0744_
rlabel metal1 10764 33626 10764 33626 0 _0745_
rlabel metal1 9890 32844 9890 32844 0 _0746_
rlabel metal1 6808 33286 6808 33286 0 _0747_
rlabel metal1 7406 32402 7406 32402 0 _0748_
rlabel metal2 7130 33082 7130 33082 0 _0749_
rlabel metal1 7360 30906 7360 30906 0 _0750_
rlabel metal2 7682 31212 7682 31212 0 _0751_
rlabel metal1 4922 32334 4922 32334 0 _0752_
rlabel metal2 6302 32096 6302 32096 0 _0753_
rlabel metal1 4291 32538 4291 32538 0 _0754_
rlabel metal1 3910 30668 3910 30668 0 _0755_
rlabel metal2 3450 33422 3450 33422 0 _0756_
rlabel metal1 3726 32878 3726 32878 0 _0757_
rlabel metal2 3358 35666 3358 35666 0 _0758_
rlabel metal1 3358 34000 3358 34000 0 _0759_
rlabel metal2 5658 36193 5658 36193 0 _0760_
rlabel metal1 5152 36278 5152 36278 0 _0761_
rlabel metal1 7682 36210 7682 36210 0 _0762_
rlabel metal1 5060 36142 5060 36142 0 _0763_
rlabel metal1 7728 36006 7728 36006 0 _0764_
rlabel metal2 8694 36380 8694 36380 0 _0765_
rlabel metal1 24196 17170 24196 17170 0 _0766_
rlabel metal1 24104 17646 24104 17646 0 _0767_
rlabel metal2 24794 17408 24794 17408 0 _0768_
rlabel metal1 24564 17578 24564 17578 0 _0769_
rlabel metal1 21942 19890 21942 19890 0 _0770_
rlabel metal1 22816 19890 22816 19890 0 _0771_
rlabel metal1 23368 19890 23368 19890 0 _0772_
rlabel metal1 23644 17034 23644 17034 0 _0773_
rlabel metal1 24932 17170 24932 17170 0 _0774_
rlabel metal1 27370 17102 27370 17102 0 _0775_
rlabel metal2 25254 16966 25254 16966 0 _0776_
rlabel metal1 25990 17102 25990 17102 0 _0777_
rlabel metal1 24932 18258 24932 18258 0 _0778_
rlabel metal2 25346 18564 25346 18564 0 _0779_
rlabel metal2 25438 18394 25438 18394 0 _0780_
rlabel metal1 24702 19380 24702 19380 0 _0781_
rlabel metal2 24886 18564 24886 18564 0 _0782_
rlabel metal2 26358 19516 26358 19516 0 _0783_
rlabel metal1 25484 18938 25484 18938 0 _0784_
rlabel metal2 26634 17476 26634 17476 0 _0785_
rlabel metal2 33534 18394 33534 18394 0 _0786_
rlabel metal1 26772 17578 26772 17578 0 _0787_
rlabel metal1 26450 17544 26450 17544 0 _0788_
rlabel metal1 28658 20944 28658 20944 0 _0789_
rlabel metal1 28520 18734 28520 18734 0 _0790_
rlabel metal2 28750 17850 28750 17850 0 _0791_
rlabel metal2 28198 17476 28198 17476 0 _0792_
rlabel metal1 29624 18190 29624 18190 0 _0793_
rlabel metal2 32154 19618 32154 19618 0 _0794_
rlabel metal2 29578 19210 29578 19210 0 _0795_
rlabel metal1 29394 17646 29394 17646 0 _0796_
rlabel metal2 26082 20094 26082 20094 0 _0797_
rlabel metal2 26910 19210 26910 19210 0 _0798_
rlabel metal2 28934 18122 28934 18122 0 _0799_
rlabel metal2 29486 17340 29486 17340 0 _0800_
rlabel metal1 29302 17102 29302 17102 0 _0801_
rlabel viali 31234 18258 31234 18258 0 _0802_
rlabel metal1 30452 16762 30452 16762 0 _0803_
rlabel metal1 29854 17204 29854 17204 0 _0804_
rlabel metal2 32798 18938 32798 18938 0 _0805_
rlabel metal1 32706 16762 32706 16762 0 _0806_
rlabel metal1 32706 17306 32706 17306 0 _0807_
rlabel metal1 32706 17204 32706 17204 0 _0808_
rlabel metal1 30774 17102 30774 17102 0 _0809_
rlabel metal1 31947 17238 31947 17238 0 _0810_
rlabel metal2 31418 16388 31418 16388 0 _0811_
rlabel metal2 30682 16524 30682 16524 0 _0812_
rlabel metal2 32246 18224 32246 18224 0 _0813_
rlabel metal1 33396 18734 33396 18734 0 _0814_
rlabel metal2 31602 20026 31602 20026 0 _0815_
rlabel metal1 34730 18836 34730 18836 0 _0816_
rlabel metal2 33626 18020 33626 18020 0 _0817_
rlabel metal2 33258 19516 33258 19516 0 _0818_
rlabel metal1 33626 19142 33626 19142 0 _0819_
rlabel metal1 32062 19414 32062 19414 0 _0820_
rlabel metal2 31418 18734 31418 18734 0 _0821_
rlabel metal2 29946 19550 29946 19550 0 _0822_
rlabel metal1 28474 17612 28474 17612 0 _0823_
rlabel metal1 27830 19380 27830 19380 0 _0824_
rlabel metal1 27186 19278 27186 19278 0 _0825_
rlabel metal2 29026 19108 29026 19108 0 _0826_
rlabel metal1 28658 18394 28658 18394 0 _0827_
rlabel metal1 29624 18258 29624 18258 0 _0828_
rlabel metal1 30866 18258 30866 18258 0 _0829_
rlabel metal1 33580 18870 33580 18870 0 _0830_
rlabel metal1 33074 18394 33074 18394 0 _0831_
rlabel metal2 34638 18428 34638 18428 0 _0832_
rlabel metal2 32154 18020 32154 18020 0 _0833_
rlabel metal2 27186 19499 27186 19499 0 _0834_
rlabel metal1 25760 21114 25760 21114 0 _0835_
rlabel metal1 27600 18938 27600 18938 0 _0836_
rlabel metal1 27692 19278 27692 19278 0 _0837_
rlabel metal1 32154 18870 32154 18870 0 _0838_
rlabel metal1 28934 18938 28934 18938 0 _0839_
rlabel metal1 28702 16082 28702 16082 0 _0840_
rlabel metal2 28290 16864 28290 16864 0 _0841_
rlabel metal1 30726 16558 30726 16558 0 _0842_
rlabel metal2 30590 16966 30590 16966 0 _0843_
rlabel metal1 32890 17544 32890 17544 0 _0844_
rlabel metal2 34270 17612 34270 17612 0 _0845_
rlabel metal1 27340 34986 27340 34986 0 _0846_
rlabel metal1 12742 17850 12742 17850 0 _0847_
rlabel metal2 15226 17952 15226 17952 0 _0848_
rlabel metal2 13294 18428 13294 18428 0 _0849_
rlabel metal2 15042 18938 15042 18938 0 _0850_
rlabel metal1 16008 18666 16008 18666 0 _0851_
rlabel metal1 14858 9078 14858 9078 0 _0852_
rlabel metal1 15272 16082 15272 16082 0 _0853_
rlabel metal2 13846 12444 13846 12444 0 _0854_
rlabel metal1 15456 16082 15456 16082 0 _0855_
rlabel metal1 15640 16150 15640 16150 0 _0856_
rlabel metal1 13294 13940 13294 13940 0 _0857_
rlabel metal2 16054 14416 16054 14416 0 _0858_
rlabel metal2 13846 15674 13846 15674 0 _0859_
rlabel metal2 15318 16388 15318 16388 0 _0860_
rlabel metal1 16744 16762 16744 16762 0 _0861_
rlabel metal2 18630 20162 18630 20162 0 _0862_
rlabel metal1 17480 18734 17480 18734 0 _0863_
rlabel metal1 13892 20910 13892 20910 0 _0864_
rlabel metal2 13478 21318 13478 21318 0 _0865_
rlabel metal1 17434 16082 17434 16082 0 _0866_
rlabel metal2 18722 18496 18722 18496 0 _0867_
rlabel viali 16790 10027 16790 10027 0 _0868_
rlabel metal1 16790 15606 16790 15606 0 _0869_
rlabel metal1 16882 15402 16882 15402 0 _0870_
rlabel via2 17342 16235 17342 16235 0 _0871_
rlabel metal2 17158 9860 17158 9860 0 _0872_
rlabel metal1 16514 9350 16514 9350 0 _0873_
rlabel metal2 15318 9146 15318 9146 0 _0874_
rlabel metal2 14582 9588 14582 9588 0 _0875_
rlabel metal1 13984 10234 13984 10234 0 _0876_
rlabel metal1 13524 10778 13524 10778 0 _0877_
rlabel metal1 13156 12410 13156 12410 0 _0878_
rlabel metal1 12788 12954 12788 12954 0 _0879_
rlabel metal1 11914 13872 11914 13872 0 _0880_
rlabel metal2 12926 14756 12926 14756 0 _0881_
rlabel metal2 13294 16116 13294 16116 0 _0882_
rlabel metal1 12788 16762 12788 16762 0 _0883_
rlabel metal1 13432 17306 13432 17306 0 _0884_
rlabel metal1 12650 18768 12650 18768 0 _0885_
rlabel metal1 13156 18938 13156 18938 0 _0886_
rlabel metal1 12880 19414 12880 19414 0 _0887_
rlabel metal1 15778 20944 15778 20944 0 _0888_
rlabel metal1 16468 21046 16468 21046 0 _0889_
rlabel metal1 18998 19822 18998 19822 0 _0890_
rlabel metal1 15778 9588 15778 9588 0 _0891_
rlabel metal2 15410 9894 15410 9894 0 _0892_
rlabel metal1 14122 13226 14122 13226 0 _0893_
rlabel metal2 13386 13634 13386 13634 0 _0894_
rlabel metal2 13754 14756 13754 14756 0 _0895_
rlabel metal1 13202 15402 13202 15402 0 _0896_
rlabel metal1 13248 18122 13248 18122 0 _0897_
rlabel metal1 13800 18394 13800 18394 0 _0898_
rlabel metal1 17986 20876 17986 20876 0 _0899_
rlabel metal2 18538 20604 18538 20604 0 _0900_
rlabel metal1 16284 15674 16284 15674 0 _0901_
rlabel metal2 15594 16388 15594 16388 0 _0902_
rlabel metal1 15088 16762 15088 16762 0 _0903_
rlabel metal1 14858 17306 14858 17306 0 _0904_
rlabel metal1 14674 18122 14674 18122 0 _0905_
rlabel metal1 14720 24718 14720 24718 0 _0906_
rlabel metal2 14398 25534 14398 25534 0 _0907_
rlabel metal2 30682 33456 30682 33456 0 _0908_
rlabel metal1 17020 13702 17020 13702 0 _0909_
rlabel metal1 10626 24752 10626 24752 0 _0910_
rlabel metal1 12880 6358 12880 6358 0 _0911_
rlabel metal2 31418 32198 31418 32198 0 _0912_
rlabel metal1 28198 23018 28198 23018 0 _0913_
rlabel metal1 25438 22746 25438 22746 0 _0914_
rlabel metal1 29532 21114 29532 21114 0 _0915_
rlabel metal1 33718 20978 33718 20978 0 _0916_
rlabel metal1 32384 21998 32384 21998 0 _0917_
rlabel metal1 35788 14314 35788 14314 0 _0918_
rlabel metal1 30176 3434 30176 3434 0 _0919_
rlabel metal1 29440 5134 29440 5134 0 _0920_
rlabel metal1 29118 6732 29118 6732 0 _0921_
rlabel metal1 22494 10506 22494 10506 0 _0922_
rlabel metal2 22586 20774 22586 20774 0 _0923_
rlabel metal1 23874 18054 23874 18054 0 _0924_
rlabel metal1 24242 13498 24242 13498 0 _0925_
rlabel metal1 17066 20502 17066 20502 0 _0926_
rlabel metal2 17894 10234 17894 10234 0 _0927_
rlabel metal1 16560 9486 16560 9486 0 _0928_
rlabel metal1 14996 8806 14996 8806 0 _0929_
rlabel metal1 21850 7820 21850 7820 0 _0930_
rlabel metal1 29118 19754 29118 19754 0 _0931_
rlabel metal1 13616 34170 13616 34170 0 _0932_
rlabel metal1 17840 34918 17840 34918 0 _0933_
rlabel metal2 17526 32538 17526 32538 0 _0934_
rlabel metal1 17710 31858 17710 31858 0 _0935_
rlabel metal2 17342 30192 17342 30192 0 _0936_
rlabel metal1 17388 30702 17388 30702 0 _0937_
rlabel metal2 18814 30124 18814 30124 0 _0938_
rlabel via1 20746 15062 20746 15062 0 _0939_
rlabel metal2 19734 14518 19734 14518 0 _0940_
rlabel metal1 19412 15062 19412 15062 0 _0941_
rlabel metal1 18032 15674 18032 15674 0 _0942_
rlabel metal1 17618 15402 17618 15402 0 _0943_
rlabel metal1 19320 13838 19320 13838 0 _0944_
rlabel metal1 8142 18292 8142 18292 0 _0945_
rlabel metal2 7498 18768 7498 18768 0 _0946_
rlabel metal1 7406 20944 7406 20944 0 _0947_
rlabel metal2 8234 24514 8234 24514 0 _0948_
rlabel metal2 8510 24956 8510 24956 0 _0949_
rlabel metal1 9108 24310 9108 24310 0 _0950_
rlabel metal2 7682 24225 7682 24225 0 _0951_
rlabel via1 7314 24259 7314 24259 0 _0952_
rlabel metal1 7084 24582 7084 24582 0 _0953_
rlabel metal2 7314 26146 7314 26146 0 _0954_
rlabel metal2 7866 24548 7866 24548 0 _0955_
rlabel metal1 8786 12138 8786 12138 0 _0956_
rlabel metal1 10488 8806 10488 8806 0 _0957_
rlabel metal1 9936 8942 9936 8942 0 _0958_
rlabel metal2 10994 5916 10994 5916 0 _0959_
rlabel metal2 11178 5236 11178 5236 0 _0960_
rlabel metal1 10994 5814 10994 5814 0 _0961_
rlabel metal1 9476 5202 9476 5202 0 _0962_
rlabel metal1 9568 5746 9568 5746 0 _0963_
rlabel metal2 9660 5746 9660 5746 0 _0964_
rlabel metal1 8832 5134 8832 5134 0 _0965_
rlabel metal1 10350 5610 10350 5610 0 _0966_
rlabel metal2 4554 18564 4554 18564 0 _0967_
rlabel metal2 4968 14994 4968 14994 0 _0968_
rlabel metal1 5336 13906 5336 13906 0 _0969_
rlabel metal1 4462 14518 4462 14518 0 _0970_
rlabel metal1 4738 14926 4738 14926 0 _0971_
rlabel metal1 4968 14586 4968 14586 0 _0972_
rlabel metal1 5474 14994 5474 14994 0 _0973_
rlabel metal1 24886 35632 24886 35632 0 _0974_
rlabel metal2 23782 35972 23782 35972 0 _0975_
rlabel metal2 29026 35768 29026 35768 0 _0976_
rlabel metal1 27232 33490 27232 33490 0 _0977_
rlabel metal2 32062 34850 32062 34850 0 _0978_
rlabel metal1 29256 36346 29256 36346 0 _0979_
rlabel metal1 29394 35802 29394 35802 0 _0980_
rlabel metal1 30314 34714 30314 34714 0 _0981_
rlabel metal1 28290 35088 28290 35088 0 _0982_
rlabel metal2 32154 34850 32154 34850 0 _0983_
rlabel metal1 25852 34578 25852 34578 0 _0984_
rlabel metal1 32016 34646 32016 34646 0 _0985_
rlabel metal1 30590 35462 30590 35462 0 _0986_
rlabel metal2 30222 35292 30222 35292 0 _0987_
rlabel metal2 30360 34578 30360 34578 0 _0988_
rlabel metal2 30498 34204 30498 34204 0 _0989_
rlabel metal1 22356 36142 22356 36142 0 _0990_
rlabel metal1 20976 33014 20976 33014 0 _0991_
rlabel metal1 20332 34646 20332 34646 0 _0992_
rlabel metal1 22034 33048 22034 33048 0 _0993_
rlabel via1 22042 32742 22042 32742 0 _0994_
rlabel metal2 21850 35224 21850 35224 0 _0995_
rlabel metal1 21528 35530 21528 35530 0 _0996_
rlabel metal2 19642 36822 19642 36822 0 _0997_
rlabel metal1 20148 35666 20148 35666 0 _0998_
rlabel metal1 20102 35598 20102 35598 0 _0999_
rlabel metal1 19918 35462 19918 35462 0 _1000_
rlabel metal2 12650 30362 12650 30362 0 _1001_
rlabel metal2 11822 31076 11822 31076 0 _1002_
rlabel metal1 10334 33558 10334 33558 0 _1003_
rlabel metal1 10396 32878 10396 32878 0 _1004_
rlabel metal2 8602 33082 8602 33082 0 _1005_
rlabel metal1 10626 32810 10626 32810 0 _1006_
rlabel metal1 6440 31994 6440 31994 0 _1007_
rlabel metal2 6946 33252 6946 33252 0 _1008_
rlabel metal1 7130 34170 7130 34170 0 _1009_
rlabel metal1 6762 34000 6762 34000 0 _1010_
rlabel metal1 8418 32810 8418 32810 0 _1011_
rlabel metal1 15134 35122 15134 35122 0 _1012_
rlabel metal1 11454 34578 11454 34578 0 _1013_
rlabel metal2 13110 35462 13110 35462 0 _1014_
rlabel metal1 15824 34714 15824 34714 0 _1015_
rlabel metal1 16606 34578 16606 34578 0 _1016_
rlabel metal2 18354 34612 18354 34612 0 _1017_
rlabel metal1 17848 31994 17848 31994 0 _1018_
rlabel metal1 15226 31212 15226 31212 0 _1019_
rlabel metal2 18630 31552 18630 31552 0 _1020_
rlabel metal2 18262 32334 18262 32334 0 _1021_
rlabel metal1 18722 32232 18722 32232 0 _1022_
rlabel metal1 18952 31994 18952 31994 0 _1023_
rlabel metal1 17204 32810 17204 32810 0 _1024_
rlabel metal1 17342 33014 17342 33014 0 _1025_
rlabel metal1 15134 31994 15134 31994 0 _1026_
rlabel metal2 14214 32708 14214 32708 0 _1027_
rlabel metal1 16330 31348 16330 31348 0 _1028_
rlabel metal1 14674 31824 14674 31824 0 _1029_
rlabel metal2 15778 30906 15778 30906 0 _1030_
rlabel metal1 16790 30294 16790 30294 0 _1031_
rlabel metal2 16698 30634 16698 30634 0 _1032_
rlabel metal2 14582 30498 14582 30498 0 _1033_
rlabel metal1 14260 30226 14260 30226 0 _1034_
rlabel metal1 14398 30736 14398 30736 0 _1035_
rlabel metal2 30774 25058 30774 25058 0 _1036_
rlabel metal1 31786 27506 31786 27506 0 _1037_
rlabel metal2 32706 27404 32706 27404 0 _1038_
rlabel metal2 35650 26724 35650 26724 0 _1039_
rlabel metal1 36708 29206 36708 29206 0 _1040_
rlabel metal2 36846 28764 36846 28764 0 _1041_
rlabel metal2 37674 28526 37674 28526 0 _1042_
rlabel metal1 37674 22032 37674 22032 0 _1043_
rlabel metal1 36064 19482 36064 19482 0 _1044_
rlabel metal2 37582 21522 37582 21522 0 _1045_
rlabel metal1 36570 19414 36570 19414 0 _1046_
rlabel metal1 37628 22610 37628 22610 0 _1047_
rlabel metal1 34086 19822 34086 19822 0 _1048_
rlabel metal2 37950 22916 37950 22916 0 _1049_
rlabel metal2 37490 23460 37490 23460 0 _1050_
rlabel metal1 38134 25160 38134 25160 0 _1051_
rlabel metal2 37306 23494 37306 23494 0 _1052_
rlabel metal1 37260 23494 37260 23494 0 _1053_
rlabel metal1 36524 22202 36524 22202 0 _1054_
rlabel metal1 36478 22542 36478 22542 0 _1055_
rlabel metal2 36202 19006 36202 19006 0 _1056_
rlabel metal1 36754 19482 36754 19482 0 _1057_
rlabel metal1 36754 23154 36754 23154 0 _1058_
rlabel metal1 37720 24106 37720 24106 0 _1059_
rlabel metal1 36846 22746 36846 22746 0 _1060_
rlabel metal1 36340 23290 36340 23290 0 _1061_
rlabel metal1 36325 24174 36325 24174 0 _1062_
rlabel metal1 35558 19380 35558 19380 0 _1063_
rlabel metal1 36294 20434 36294 20434 0 _1064_
rlabel metal2 37858 20740 37858 20740 0 _1065_
rlabel metal1 37306 19890 37306 19890 0 _1066_
rlabel metal1 36386 20842 36386 20842 0 _1067_
rlabel metal2 36754 20128 36754 20128 0 _1068_
rlabel metal2 36018 20060 36018 20060 0 _1069_
rlabel metal2 36064 20910 36064 20910 0 _1070_
rlabel metal1 35926 24276 35926 24276 0 _1071_
rlabel metal2 36846 24548 36846 24548 0 _1072_
rlabel metal1 35696 24718 35696 24718 0 _1073_
rlabel metal1 35512 20570 35512 20570 0 _1074_
rlabel metal1 35972 21114 35972 21114 0 _1075_
rlabel metal1 36662 20944 36662 20944 0 _1076_
rlabel metal1 36064 21522 36064 21522 0 _1077_
rlabel viali 33840 19819 33840 19819 0 _1078_
rlabel metal2 33626 20162 33626 20162 0 _1079_
rlabel metal2 33902 20638 33902 20638 0 _1080_
rlabel metal1 34960 21590 34960 21590 0 _1081_
rlabel metal1 35190 21658 35190 21658 0 _1082_
rlabel metal1 34408 21998 34408 21998 0 _1083_
rlabel metal2 35374 21828 35374 21828 0 _1084_
rlabel metal1 34822 21998 34822 21998 0 _1085_
rlabel metal2 34454 22406 34454 22406 0 _1086_
rlabel metal1 35282 23698 35282 23698 0 _1087_
rlabel metal2 34822 23222 34822 23222 0 _1088_
rlabel metal1 34868 24786 34868 24786 0 _1089_
rlabel metal1 34684 22202 34684 22202 0 _1090_
rlabel metal2 34638 23222 34638 23222 0 _1091_
rlabel metal2 33902 21318 33902 21318 0 _1092_
rlabel metal1 33718 22542 33718 22542 0 _1093_
rlabel metal1 32568 20910 32568 20910 0 _1094_
rlabel metal1 31878 20434 31878 20434 0 _1095_
rlabel metal2 31786 21284 31786 21284 0 _1096_
rlabel metal2 32706 21726 32706 21726 0 _1097_
rlabel metal1 33074 22508 33074 22508 0 _1098_
rlabel metal2 33074 21522 33074 21522 0 _1099_
rlabel metal1 32844 22406 32844 22406 0 _1100_
rlabel metal1 33718 22678 33718 22678 0 _1101_
rlabel metal2 34362 23222 34362 23222 0 _1102_
rlabel metal1 34546 24582 34546 24582 0 _1103_
rlabel metal2 34546 24004 34546 24004 0 _1104_
rlabel metal1 33994 24752 33994 24752 0 _1105_
rlabel metal1 33212 22202 33212 22202 0 _1106_
rlabel metal1 33166 23732 33166 23732 0 _1107_
rlabel metal1 30682 22576 30682 22576 0 _1108_
rlabel metal2 30406 21114 30406 21114 0 _1109_
rlabel metal2 30314 22950 30314 22950 0 _1110_
rlabel metal2 31786 22780 31786 22780 0 _1111_
rlabel metal1 32476 22202 32476 22202 0 _1112_
rlabel metal2 32154 22916 32154 22916 0 _1113_
rlabel metal1 32752 23698 32752 23698 0 _1114_
rlabel metal1 33304 24786 33304 24786 0 _1115_
rlabel metal2 32890 24004 32890 24004 0 _1116_
rlabel metal2 32706 24582 32706 24582 0 _1117_
rlabel metal1 31556 23290 31556 23290 0 _1118_
rlabel metal1 31694 24140 31694 24140 0 _1119_
rlabel metal1 30360 23630 30360 23630 0 _1120_
rlabel metal1 29026 21658 29026 21658 0 _1121_
rlabel metal1 28474 22066 28474 22066 0 _1122_
rlabel metal1 29118 22644 29118 22644 0 _1123_
rlabel metal2 30222 23222 30222 23222 0 _1124_
rlabel metal2 30406 23970 30406 23970 0 _1125_
rlabel metal1 32292 24786 32292 24786 0 _1126_
rlabel metal1 31786 24208 31786 24208 0 _1127_
rlabel metal2 31602 24616 31602 24616 0 _1128_
rlabel metal1 30406 23834 30406 23834 0 _1129_
rlabel metal1 28934 24242 28934 24242 0 _1130_
rlabel metal2 28842 23494 28842 23494 0 _1131_
rlabel metal1 29762 24208 29762 24208 0 _1132_
rlabel metal2 29210 20468 29210 20468 0 _1133_
rlabel metal2 27278 20876 27278 20876 0 _1134_
rlabel metal2 29578 24548 29578 24548 0 _1135_
rlabel metal1 29624 24786 29624 24786 0 _1136_
rlabel metal1 31970 24786 31970 24786 0 _1137_
rlabel metal1 32798 25228 32798 25228 0 _1138_
rlabel metal2 33626 25058 33626 25058 0 _1139_
rlabel metal2 34914 24922 34914 24922 0 _1140_
rlabel metal1 35926 25806 35926 25806 0 _1141_
rlabel metal2 36662 23936 36662 23936 0 _1142_
rlabel metal2 37030 24582 37030 24582 0 _1143_
rlabel metal1 37398 25228 37398 25228 0 _1144_
rlabel metal1 37582 26418 37582 26418 0 _1145_
rlabel metal1 37306 27574 37306 27574 0 _1146_
rlabel metal2 37858 25670 37858 25670 0 _1147_
rlabel viali 37565 27438 37565 27438 0 _1148_
rlabel metal1 35512 28594 35512 28594 0 _1149_
rlabel metal1 37214 27302 37214 27302 0 _1150_
rlabel metal1 37720 27438 37720 27438 0 _1151_
rlabel metal2 37030 28730 37030 28730 0 _1152_
rlabel metal2 37582 28288 37582 28288 0 _1153_
rlabel metal2 38042 27676 38042 27676 0 _1154_
rlabel metal1 36478 26996 36478 26996 0 _1155_
rlabel metal1 36800 25262 36800 25262 0 _1156_
rlabel metal1 36524 26350 36524 26350 0 _1157_
rlabel metal1 36478 26894 36478 26894 0 _1158_
rlabel metal2 35466 25398 35466 25398 0 _1159_
rlabel metal1 35328 26554 35328 26554 0 _1160_
rlabel metal1 35558 25908 35558 25908 0 _1161_
rlabel metal1 36202 26010 36202 26010 0 _1162_
rlabel metal1 34638 24922 34638 24922 0 _1163_
rlabel metal2 34362 25670 34362 25670 0 _1164_
rlabel metal2 32154 28594 32154 28594 0 _1165_
rlabel metal2 33626 26316 33626 26316 0 _1166_
rlabel metal1 34730 25806 34730 25806 0 _1167_
rlabel metal1 32798 25908 32798 25908 0 _1168_
rlabel metal2 31510 27642 31510 27642 0 _1169_
rlabel metal2 32430 26656 32430 26656 0 _1170_
rlabel metal2 33442 25092 33442 25092 0 _1171_
rlabel metal2 33166 25636 33166 25636 0 _1172_
rlabel metal2 32706 25092 32706 25092 0 _1173_
rlabel metal1 32430 25466 32430 25466 0 _1174_
rlabel metal2 31142 26690 31142 26690 0 _1175_
rlabel metal2 32246 24956 32246 24956 0 _1176_
rlabel metal2 31142 24990 31142 24990 0 _1177_
rlabel metal2 30958 25738 30958 25738 0 _1178_
rlabel metal1 31280 24922 31280 24922 0 _1179_
rlabel metal2 29026 24242 29026 24242 0 _1180_
rlabel metal2 29118 24956 29118 24956 0 _1181_
rlabel via1 27646 20842 27646 20842 0 _1182_
rlabel metal1 30912 20434 30912 20434 0 _1183_
rlabel metal1 28152 20910 28152 20910 0 _1184_
rlabel metal1 28152 18258 28152 18258 0 _1185_
rlabel metal1 28244 18394 28244 18394 0 _1186_
rlabel metal2 27830 23290 27830 23290 0 _1187_
rlabel metal1 26818 21998 26818 21998 0 _1188_
rlabel metal1 27508 22066 27508 22066 0 _1189_
rlabel metal2 26818 22916 26818 22916 0 _1190_
rlabel metal1 27554 23120 27554 23120 0 _1191_
rlabel metal1 28198 22202 28198 22202 0 _1192_
rlabel metal1 27692 22746 27692 22746 0 _1193_
rlabel metal1 27416 23086 27416 23086 0 _1194_
rlabel metal1 28152 23290 28152 23290 0 _1195_
rlabel metal2 28290 23800 28290 23800 0 _1196_
rlabel metal1 27876 24378 27876 24378 0 _1197_
rlabel metal1 31418 25330 31418 25330 0 _1198_
rlabel metal1 31510 25398 31510 25398 0 _1199_
rlabel metal1 32476 25126 32476 25126 0 _1200_
rlabel metal1 33074 25772 33074 25772 0 _1201_
rlabel metal1 34776 25874 34776 25874 0 _1202_
rlabel metal1 35880 26010 35880 26010 0 _1203_
rlabel metal2 36570 26758 36570 26758 0 _1204_
rlabel metal1 37490 27098 37490 27098 0 _1205_
rlabel metal1 38180 27642 38180 27642 0 _1206_
rlabel metal2 37306 28900 37306 28900 0 _1207_
rlabel metal1 37858 28186 37858 28186 0 _1208_
rlabel metal1 32890 29818 32890 29818 0 _1209_
rlabel metal1 32660 30226 32660 30226 0 _1210_
rlabel metal2 37490 29274 37490 29274 0 _1211_
rlabel metal1 32798 30668 32798 30668 0 _1212_
rlabel metal1 32982 29274 32982 29274 0 _1213_
rlabel metal1 32430 30736 32430 30736 0 _1214_
rlabel metal1 32016 30906 32016 30906 0 _1215_
rlabel metal2 23966 23290 23966 23290 0 _1216_
rlabel metal1 25346 25466 25346 25466 0 _1217_
rlabel metal1 25116 24378 25116 24378 0 _1218_
rlabel metal1 25530 25228 25530 25228 0 _1219_
rlabel metal2 27002 25092 27002 25092 0 _1220_
rlabel metal1 29440 26350 29440 26350 0 _1221_
rlabel metal1 28428 25670 28428 25670 0 _1222_
rlabel metal1 28152 26554 28152 26554 0 _1223_
rlabel metal1 30452 28526 30452 28526 0 _1224_
rlabel metal1 30774 28390 30774 28390 0 _1225_
rlabel metal1 29118 28560 29118 28560 0 _1226_
rlabel metal1 28566 29512 28566 29512 0 _1227_
rlabel metal1 30452 28730 30452 28730 0 _1228_
rlabel metal1 34408 29138 34408 29138 0 _1229_
rlabel metal1 33212 28526 33212 28526 0 _1230_
rlabel metal1 34546 28084 34546 28084 0 _1231_
rlabel metal2 33074 27914 33074 27914 0 _1232_
rlabel metal1 34454 29274 34454 29274 0 _1233_
rlabel metal1 33948 29614 33948 29614 0 _1234_
rlabel metal2 34546 30430 34546 30430 0 _1235_
rlabel metal1 35282 30362 35282 30362 0 _1236_
rlabel via1 33902 32402 33902 32402 0 _1237_
rlabel metal1 34270 32946 34270 32946 0 _1238_
rlabel metal2 34638 32708 34638 32708 0 _1239_
rlabel metal1 33810 32810 33810 32810 0 _1240_
rlabel metal1 32614 32198 32614 32198 0 _1241_
rlabel metal1 32928 32538 32928 32538 0 _1242_
rlabel metal1 31786 3468 31786 3468 0 _1243_
rlabel metal2 31326 3366 31326 3366 0 _1244_
rlabel metal1 30820 3502 30820 3502 0 _1245_
rlabel metal1 26174 4080 26174 4080 0 _1246_
rlabel metal2 27738 3332 27738 3332 0 _1247_
rlabel metal1 27140 3570 27140 3570 0 _1248_
rlabel metal1 26220 4250 26220 4250 0 _1249_
rlabel metal1 28014 4012 28014 4012 0 _1250_
rlabel metal2 27922 4182 27922 4182 0 _1251_
rlabel metal1 27646 3604 27646 3604 0 _1252_
rlabel metal1 32859 4114 32859 4114 0 _1253_
rlabel metal2 31142 3808 31142 3808 0 _1254_
rlabel metal2 32338 3332 32338 3332 0 _1255_
rlabel metal1 32430 4046 32430 4046 0 _1256_
rlabel metal1 34040 4658 34040 4658 0 _1257_
rlabel metal2 33166 4658 33166 4658 0 _1258_
rlabel metal1 32154 5236 32154 5236 0 _1259_
rlabel metal2 27830 4454 27830 4454 0 _1260_
rlabel metal1 28382 4590 28382 4590 0 _1261_
rlabel metal2 28566 3230 28566 3230 0 _1262_
rlabel metal2 29578 3876 29578 3876 0 _1263_
rlabel metal2 28658 4454 28658 4454 0 _1264_
rlabel metal1 29946 5168 29946 5168 0 _1265_
rlabel metal2 29394 4998 29394 4998 0 _1266_
rlabel via1 29854 5338 29854 5338 0 _1267_
rlabel metal1 30406 5134 30406 5134 0 _1268_
rlabel metal1 31142 3162 31142 3162 0 _1269_
rlabel metal1 32062 5168 32062 5168 0 _1270_
rlabel metal1 32660 5202 32660 5202 0 _1271_
rlabel metal1 32522 5236 32522 5236 0 _1272_
rlabel metal2 32798 5508 32798 5508 0 _1273_
rlabel metal1 29670 5338 29670 5338 0 _1274_
rlabel metal2 30682 6086 30682 6086 0 _1275_
rlabel metal1 29532 3706 29532 3706 0 _1276_
rlabel metal1 28980 6290 28980 6290 0 _1277_
rlabel metal3 575 33796 575 33796 0 clk
rlabel via2 14214 14331 14214 14331 0 clknet_0_clk
rlabel metal1 15088 14382 15088 14382 0 clknet_2_0__leaf_clk
rlabel metal2 18722 33116 18722 33116 0 clknet_2_1__leaf_clk
rlabel metal1 34270 16082 34270 16082 0 clknet_2_2__leaf_clk
rlabel metal1 32890 34510 32890 34510 0 clknet_2_3__leaf_clk
rlabel metal2 2530 11696 2530 11696 0 clknet_leaf_0_clk
rlabel metal2 19366 32708 19366 32708 0 clknet_leaf_10_clk
rlabel metal1 12880 29070 12880 29070 0 clknet_leaf_11_clk
rlabel metal2 19274 21522 19274 21522 0 clknet_leaf_12_clk
rlabel metal1 21574 29614 21574 29614 0 clknet_leaf_13_clk
rlabel metal1 21114 31790 21114 31790 0 clknet_leaf_14_clk
rlabel metal1 27002 35700 27002 35700 0 clknet_leaf_15_clk
rlabel metal1 32890 34034 32890 34034 0 clknet_leaf_16_clk
rlabel metal2 35466 28016 35466 28016 0 clknet_leaf_17_clk
rlabel metal1 27646 23630 27646 23630 0 clknet_leaf_18_clk
rlabel metal2 24978 18156 24978 18156 0 clknet_leaf_19_clk
rlabel metal1 1472 18190 1472 18190 0 clknet_leaf_1_clk
rlabel metal2 36754 13872 36754 13872 0 clknet_leaf_20_clk
rlabel metal1 35374 13362 35374 13362 0 clknet_leaf_21_clk
rlabel metal1 23460 3434 23460 3434 0 clknet_leaf_23_clk
rlabel metal1 21850 13940 21850 13940 0 clknet_leaf_24_clk
rlabel metal1 19044 15470 19044 15470 0 clknet_leaf_25_clk
rlabel metal2 15778 13600 15778 13600 0 clknet_leaf_26_clk
rlabel metal2 15870 5168 15870 5168 0 clknet_leaf_27_clk
rlabel metal2 14490 7990 14490 7990 0 clknet_leaf_28_clk
rlabel metal2 2668 6868 2668 6868 0 clknet_leaf_29_clk
rlabel metal2 12742 15266 12742 15266 0 clknet_leaf_2_clk
rlabel metal2 12558 20978 12558 20978 0 clknet_leaf_3_clk
rlabel metal1 10074 20910 10074 20910 0 clknet_leaf_4_clk
rlabel metal1 1748 22542 1748 22542 0 clknet_leaf_5_clk
rlabel metal2 2714 25806 2714 25806 0 clknet_leaf_6_clk
rlabel metal2 8970 29104 8970 29104 0 clknet_leaf_7_clk
rlabel metal1 2070 31994 2070 31994 0 clknet_leaf_8_clk
rlabel metal1 15870 34034 15870 34034 0 clknet_leaf_9_clk
rlabel metal2 21482 10234 21482 10234 0 dut.actual_duty_x\[0\]
rlabel metal1 21620 9622 21620 9622 0 dut.actual_duty_x\[1\]
rlabel metal2 21850 8670 21850 8670 0 dut.actual_duty_x\[2\]
rlabel metal2 21482 7140 21482 7140 0 dut.actual_duty_x\[3\]
rlabel metal1 21735 5202 21735 5202 0 dut.actual_duty_x\[4\]
rlabel metal2 27186 4811 27186 4811 0 dut.actual_duty_x\[5\]
rlabel metal1 29072 3026 29072 3026 0 dut.actual_duty_x\[6\]
rlabel metal2 27002 3196 27002 3196 0 dut.actual_duty_x\[7\]
rlabel metal2 25898 21046 25898 21046 0 dut.actual_duty_y\[0\]
rlabel metal1 28750 21998 28750 21998 0 dut.actual_duty_y\[1\]
rlabel via2 33074 20485 33074 20485 0 dut.actual_duty_y\[2\]
rlabel via2 33074 20859 33074 20859 0 dut.actual_duty_y\[3\]
rlabel metal1 32108 17170 32108 17170 0 dut.actual_duty_y\[4\]
rlabel metal1 33718 17578 33718 17578 0 dut.actual_duty_y\[5\]
rlabel metal1 37076 18734 37076 18734 0 dut.actual_duty_y\[6\]
rlabel metal2 37122 18258 37122 18258 0 dut.actual_duty_y\[7\]
rlabel metal1 20194 20230 20194 20230 0 dut.ball_pos_x\[0\]
rlabel metal1 18998 20298 18998 20298 0 dut.ball_pos_x\[1\]
rlabel metal2 17618 18530 17618 18530 0 dut.ball_pos_x\[2\]
rlabel metal1 18492 18734 18492 18734 0 dut.ball_pos_y\[0\]
rlabel metal1 21436 18734 21436 18734 0 dut.ball_pos_y\[1\]
rlabel metal2 21482 19176 21482 19176 0 dut.ball_pos_y\[2\]
rlabel metal1 14996 14518 14996 14518 0 dut.clk_en
rlabel metal1 5014 12410 5014 12410 0 dut.clkdiv_inst.counter\[0\]
rlabel metal1 5290 16694 5290 16694 0 dut.clkdiv_inst.counter\[10\]
rlabel metal2 5106 17918 5106 17918 0 dut.clkdiv_inst.counter\[11\]
rlabel metal2 4462 17442 4462 17442 0 dut.clkdiv_inst.counter\[12\]
rlabel metal1 3496 18938 3496 18938 0 dut.clkdiv_inst.counter\[13\]
rlabel metal1 4048 18734 4048 18734 0 dut.clkdiv_inst.counter\[14\]
rlabel metal1 4508 19822 4508 19822 0 dut.clkdiv_inst.counter\[15\]
rlabel metal1 4738 18700 4738 18700 0 dut.clkdiv_inst.counter\[16\]
rlabel metal1 5014 12104 5014 12104 0 dut.clkdiv_inst.counter\[1\]
rlabel viali 4822 12138 4822 12138 0 dut.clkdiv_inst.counter\[2\]
rlabel metal1 7498 13906 7498 13906 0 dut.clkdiv_inst.counter\[3\]
rlabel metal1 5106 14450 5106 14450 0 dut.clkdiv_inst.counter\[4\]
rlabel metal2 2714 13889 2714 13889 0 dut.clkdiv_inst.counter\[5\]
rlabel metal1 5704 14450 5704 14450 0 dut.clkdiv_inst.counter\[6\]
rlabel metal1 4002 14926 4002 14926 0 dut.clkdiv_inst.counter\[7\]
rlabel metal1 2254 17136 2254 17136 0 dut.clkdiv_inst.counter\[8\]
rlabel metal1 4784 15334 4784 15334 0 dut.clkdiv_inst.counter\[9\]
rlabel metal1 2162 10574 2162 10574 0 dut.clkdiv_inst.reset_n
rlabel metal1 3956 18938 3956 18938 0 dut.clkdiv_inst.sck
rlabel metal2 24426 36550 24426 36550 0 dut.cs_n_lcd
rlabel metal1 23230 30838 23230 30838 0 dut.data_in\[0\]
rlabel metal2 23138 29342 23138 29342 0 dut.data_in\[1\]
rlabel metal2 20286 29410 20286 29410 0 dut.data_in\[2\]
rlabel metal1 24150 26010 24150 26010 0 dut.data_in\[3\]
rlabel metal1 24840 24582 24840 24582 0 dut.data_in\[4\]
rlabel metal1 24058 27302 24058 27302 0 dut.data_in\[5\]
rlabel metal1 23782 28594 23782 28594 0 dut.data_in\[6\]
rlabel metal1 20746 29206 20746 29206 0 dut.data_in\[7\]
rlabel metal1 23506 31858 23506 31858 0 dut.data_in\[9\]
rlabel metal1 18906 16762 18906 16762 0 dut.ir_sensor_array.bit_count\[0\]
rlabel metal1 20010 15334 20010 15334 0 dut.ir_sensor_array.bit_count\[1\]
rlabel metal1 21068 16422 21068 16422 0 dut.ir_sensor_array.bit_count\[2\]
rlabel metal1 20240 14586 20240 14586 0 dut.ir_sensor_array.bit_count\[3\]
rlabel metal2 20286 13668 20286 13668 0 dut.ir_sensor_array.bit_count\[4\]
rlabel metal1 20608 12750 20608 12750 0 dut.ir_sensor_array.bit_count\[5\]
rlabel metal1 13708 13430 13708 13430 0 dut.ir_sensor_array.final_sensor_data\[10\]
rlabel metal1 13478 13294 13478 13294 0 dut.ir_sensor_array.final_sensor_data\[11\]
rlabel metal2 13110 9758 13110 9758 0 dut.ir_sensor_array.final_sensor_data\[12\]
rlabel metal1 13754 8942 13754 8942 0 dut.ir_sensor_array.final_sensor_data\[13\]
rlabel metal1 15042 9588 15042 9588 0 dut.ir_sensor_array.final_sensor_data\[14\]
rlabel metal2 14858 12789 14858 12789 0 dut.ir_sensor_array.final_sensor_data\[15\]
rlabel metal2 14030 13498 14030 13498 0 dut.ir_sensor_array.final_sensor_data\[16\]
rlabel metal2 14858 15776 14858 15776 0 dut.ir_sensor_array.final_sensor_data\[17\]
rlabel metal2 13662 15810 13662 15810 0 dut.ir_sensor_array.final_sensor_data\[18\]
rlabel metal2 13570 15674 13570 15674 0 dut.ir_sensor_array.final_sensor_data\[19\]
rlabel metal1 16008 8942 16008 8942 0 dut.ir_sensor_array.final_sensor_data\[1\]
rlabel metal1 11776 13906 11776 13906 0 dut.ir_sensor_array.final_sensor_data\[20\]
rlabel metal2 12650 13634 12650 13634 0 dut.ir_sensor_array.final_sensor_data\[21\]
rlabel metal1 13110 13872 13110 13872 0 dut.ir_sensor_array.final_sensor_data\[22\]
rlabel metal1 13156 13294 13156 13294 0 dut.ir_sensor_array.final_sensor_data\[23\]
rlabel metal1 14168 15130 14168 15130 0 dut.ir_sensor_array.final_sensor_data\[24\]
rlabel metal1 14306 19414 14306 19414 0 dut.ir_sensor_array.final_sensor_data\[25\]
rlabel metal2 13478 18700 13478 18700 0 dut.ir_sensor_array.final_sensor_data\[26\]
rlabel metal2 13386 18938 13386 18938 0 dut.ir_sensor_array.final_sensor_data\[27\]
rlabel metal1 12834 17578 12834 17578 0 dut.ir_sensor_array.final_sensor_data\[28\]
rlabel metal1 13018 17612 13018 17612 0 dut.ir_sensor_array.final_sensor_data\[29\]
rlabel metal2 16422 9486 16422 9486 0 dut.ir_sensor_array.final_sensor_data\[2\]
rlabel metal1 13524 17646 13524 17646 0 dut.ir_sensor_array.final_sensor_data\[30\]
rlabel metal1 15824 17850 15824 17850 0 dut.ir_sensor_array.final_sensor_data\[31\]
rlabel metal1 17204 18802 17204 18802 0 dut.ir_sensor_array.final_sensor_data\[32\]
rlabel metal1 16560 20434 16560 20434 0 dut.ir_sensor_array.final_sensor_data\[33\]
rlabel metal2 17986 21284 17986 21284 0 dut.ir_sensor_array.final_sensor_data\[34\]
rlabel metal1 18078 20842 18078 20842 0 dut.ir_sensor_array.final_sensor_data\[35\]
rlabel metal2 15594 21114 15594 21114 0 dut.ir_sensor_array.final_sensor_data\[36\]
rlabel metal1 13846 22066 13846 22066 0 dut.ir_sensor_array.final_sensor_data\[37\]
rlabel metal1 14076 20978 14076 20978 0 dut.ir_sensor_array.final_sensor_data\[38\]
rlabel metal1 14168 20842 14168 20842 0 dut.ir_sensor_array.final_sensor_data\[39\]
rlabel metal2 17802 7956 17802 7956 0 dut.ir_sensor_array.final_sensor_data\[3\]
rlabel metal1 18584 8806 18584 8806 0 dut.ir_sensor_array.final_sensor_data\[4\]
rlabel metal1 17434 9996 17434 9996 0 dut.ir_sensor_array.final_sensor_data\[5\]
rlabel metal2 18538 10234 18538 10234 0 dut.ir_sensor_array.final_sensor_data\[6\]
rlabel metal2 18446 11968 18446 11968 0 dut.ir_sensor_array.final_sensor_data\[7\]
rlabel metal1 13432 12818 13432 12818 0 dut.ir_sensor_array.final_sensor_data\[8\]
rlabel metal1 14168 12750 14168 12750 0 dut.ir_sensor_array.final_sensor_data\[9\]
rlabel metal1 20424 11730 20424 11730 0 dut.ir_sensor_array.latch
rlabel metal1 17986 13906 17986 13906 0 dut.ir_sensor_array.state\[0\]
rlabel metal1 19044 14994 19044 14994 0 dut.ir_sensor_array.state\[1\]
rlabel metal1 18998 12954 18998 12954 0 dut.ir_sensor_array.state\[2\]
rlabel metal1 10074 29478 10074 29478 0 dut.lcd1602.cnt_200ms\[0\]
rlabel metal1 6314 31858 6314 31858 0 dut.lcd1602.cnt_200ms\[10\]
rlabel metal2 6762 31552 6762 31552 0 dut.lcd1602.cnt_200ms\[11\]
rlabel metal2 5842 31484 5842 31484 0 dut.lcd1602.cnt_200ms\[12\]
rlabel metal1 4002 31892 4002 31892 0 dut.lcd1602.cnt_200ms\[13\]
rlabel metal2 5658 32538 5658 32538 0 dut.lcd1602.cnt_200ms\[14\]
rlabel metal1 4278 33422 4278 33422 0 dut.lcd1602.cnt_200ms\[15\]
rlabel metal2 5106 34204 5106 34204 0 dut.lcd1602.cnt_200ms\[16\]
rlabel metal2 6118 35428 6118 35428 0 dut.lcd1602.cnt_200ms\[17\]
rlabel metal1 6624 36142 6624 36142 0 dut.lcd1602.cnt_200ms\[18\]
rlabel metal1 7268 36074 7268 36074 0 dut.lcd1602.cnt_200ms\[19\]
rlabel metal1 11845 29070 11845 29070 0 dut.lcd1602.cnt_200ms\[1\]
rlabel metal1 8234 35802 8234 35802 0 dut.lcd1602.cnt_200ms\[20\]
rlabel metal1 8694 35156 8694 35156 0 dut.lcd1602.cnt_200ms\[21\]
rlabel metal2 12926 28934 12926 28934 0 dut.lcd1602.cnt_200ms\[2\]
rlabel metal1 11960 30770 11960 30770 0 dut.lcd1602.cnt_200ms\[3\]
rlabel metal2 11822 32810 11822 32810 0 dut.lcd1602.cnt_200ms\[4\]
rlabel metal2 11362 32028 11362 32028 0 dut.lcd1602.cnt_200ms\[5\]
rlabel metal1 10074 33388 10074 33388 0 dut.lcd1602.cnt_200ms\[6\]
rlabel metal1 8924 32946 8924 32946 0 dut.lcd1602.cnt_200ms\[7\]
rlabel metal2 7498 32606 7498 32606 0 dut.lcd1602.cnt_200ms\[8\]
rlabel metal1 6992 31858 6992 31858 0 dut.lcd1602.cnt_200ms\[9\]
rlabel metal2 13478 34612 13478 34612 0 dut.lcd1602.cnt_500hz\[0\]
rlabel metal1 15410 31790 15410 31790 0 dut.lcd1602.cnt_500hz\[10\]
rlabel metal1 16192 30362 16192 30362 0 dut.lcd1602.cnt_500hz\[11\]
rlabel metal1 17388 30362 17388 30362 0 dut.lcd1602.cnt_500hz\[12\]
rlabel metal2 15042 29886 15042 29886 0 dut.lcd1602.cnt_500hz\[13\]
rlabel metal1 15134 30158 15134 30158 0 dut.lcd1602.cnt_500hz\[14\]
rlabel metal2 13110 34544 13110 34544 0 dut.lcd1602.cnt_500hz\[1\]
rlabel metal2 13938 34884 13938 34884 0 dut.lcd1602.cnt_500hz\[2\]
rlabel metal2 15042 34476 15042 34476 0 dut.lcd1602.cnt_500hz\[3\]
rlabel metal1 18216 33830 18216 33830 0 dut.lcd1602.cnt_500hz\[4\]
rlabel metal2 17434 34850 17434 34850 0 dut.lcd1602.cnt_500hz\[5\]
rlabel metal1 17434 31926 17434 31926 0 dut.lcd1602.cnt_500hz\[6\]
rlabel metal1 17618 32810 17618 32810 0 dut.lcd1602.cnt_500hz\[7\]
rlabel metal1 18308 32198 18308 32198 0 dut.lcd1602.cnt_500hz\[8\]
rlabel metal2 16330 33150 16330 33150 0 dut.lcd1602.cnt_500hz\[9\]
rlabel metal1 13432 24786 13432 24786 0 dut.lcd1602.currentState\[0\]
rlabel metal1 12926 24174 12926 24174 0 dut.lcd1602.currentState\[1\]
rlabel metal1 13938 27982 13938 27982 0 dut.lcd1602.currentState\[2\]
rlabel metal1 15318 27438 15318 27438 0 dut.lcd1602.currentState\[3\]
rlabel metal1 18538 28186 18538 28186 0 dut.lcd1602.currentState\[4\]
rlabel metal1 16652 22066 16652 22066 0 dut.lcd1602.currentState\[5\]
rlabel metal1 19320 29750 19320 29750 0 dut.lcd1602.lcd_ctrl
rlabel metal1 24610 32436 24610 32436 0 dut.lcd1602.out_valid
rlabel metal1 21758 10098 21758 10098 0 dut.microstep_x.clk_en
rlabel metal1 8602 12682 8602 12682 0 dut.microstep_x.ctr\[0\]
rlabel metal1 11178 4590 11178 4590 0 dut.microstep_x.ctr\[10\]
rlabel metal1 13156 3502 13156 3502 0 dut.microstep_x.ctr\[11\]
rlabel metal1 10258 3604 10258 3604 0 dut.microstep_x.ctr\[12\]
rlabel metal1 9154 4556 9154 4556 0 dut.microstep_x.ctr\[13\]
rlabel metal1 9108 2482 9108 2482 0 dut.microstep_x.ctr\[14\]
rlabel metal2 8602 7038 8602 7038 0 dut.microstep_x.ctr\[15\]
rlabel viali 10153 6222 10153 6222 0 dut.microstep_x.ctr\[16\]
rlabel metal1 6762 5236 6762 5236 0 dut.microstep_x.ctr\[17\]
rlabel metal2 6578 4454 6578 4454 0 dut.microstep_x.ctr\[18\]
rlabel metal2 7130 3910 7130 3910 0 dut.microstep_x.ctr\[19\]
rlabel metal1 9154 12274 9154 12274 0 dut.microstep_x.ctr\[1\]
rlabel metal1 4462 3706 4462 3706 0 dut.microstep_x.ctr\[20\]
rlabel metal2 5014 3672 5014 3672 0 dut.microstep_x.ctr\[21\]
rlabel metal1 4140 5746 4140 5746 0 dut.microstep_x.ctr\[22\]
rlabel metal1 5244 6290 5244 6290 0 dut.microstep_x.ctr\[23\]
rlabel metal1 3726 6970 3726 6970 0 dut.microstep_x.ctr\[24\]
rlabel metal1 4600 7174 4600 7174 0 dut.microstep_x.ctr\[25\]
rlabel metal2 6026 8364 6026 8364 0 dut.microstep_x.ctr\[26\]
rlabel metal1 7130 8500 7130 8500 0 dut.microstep_x.ctr\[27\]
rlabel metal2 9154 8058 9154 8058 0 dut.microstep_x.ctr\[28\]
rlabel metal2 8142 9316 8142 9316 0 dut.microstep_x.ctr\[29\]
rlabel metal2 9798 12036 9798 12036 0 dut.microstep_x.ctr\[2\]
rlabel metal1 8464 10438 8464 10438 0 dut.microstep_x.ctr\[3\]
rlabel metal1 11454 10574 11454 10574 0 dut.microstep_x.ctr\[4\]
rlabel metal2 10902 9112 10902 9112 0 dut.microstep_x.ctr\[5\]
rlabel via1 11730 8398 11730 8398 0 dut.microstep_x.ctr\[6\]
rlabel metal2 11546 7242 11546 7242 0 dut.microstep_x.ctr\[7\]
rlabel metal1 14306 6766 14306 6766 0 dut.microstep_x.ctr\[8\]
rlabel metal1 13616 5678 13616 5678 0 dut.microstep_x.ctr\[9\]
rlabel metal1 34316 17034 34316 17034 0 dut.microstep_y.clk_en
rlabel metal2 7590 16660 7590 16660 0 dut.microstep_y.ctr\[0\]
rlabel metal1 11638 26894 11638 26894 0 dut.microstep_y.ctr\[10\]
rlabel metal1 9614 26350 9614 26350 0 dut.microstep_y.ctr\[11\]
rlabel metal1 8234 25466 8234 25466 0 dut.microstep_y.ctr\[12\]
rlabel metal1 6486 24786 6486 24786 0 dut.microstep_y.ctr\[13\]
rlabel metal1 6164 24922 6164 24922 0 dut.microstep_y.ctr\[14\]
rlabel metal1 7728 24106 7728 24106 0 dut.microstep_y.ctr\[15\]
rlabel metal2 6854 22916 6854 22916 0 dut.microstep_y.ctr\[16\]
rlabel metal1 5198 21522 5198 21522 0 dut.microstep_y.ctr\[17\]
rlabel metal2 4002 23936 4002 23936 0 dut.microstep_y.ctr\[18\]
rlabel metal1 3404 23630 3404 23630 0 dut.microstep_y.ctr\[19\]
rlabel metal1 7406 17510 7406 17510 0 dut.microstep_y.ctr\[1\]
rlabel metal1 3312 24106 3312 24106 0 dut.microstep_y.ctr\[20\]
rlabel metal2 4738 24684 4738 24684 0 dut.microstep_y.ctr\[21\]
rlabel metal2 4002 27846 4002 27846 0 dut.microstep_y.ctr\[22\]
rlabel metal1 4370 27438 4370 27438 0 dut.microstep_y.ctr\[23\]
rlabel metal1 3864 27982 3864 27982 0 dut.microstep_y.ctr\[24\]
rlabel metal2 3358 28016 3358 28016 0 dut.microstep_y.ctr\[25\]
rlabel metal1 5658 27880 5658 27880 0 dut.microstep_y.ctr\[26\]
rlabel metal1 6900 28594 6900 28594 0 dut.microstep_y.ctr\[27\]
rlabel metal2 8234 28220 8234 28220 0 dut.microstep_y.ctr\[28\]
rlabel metal1 7452 28526 7452 28526 0 dut.microstep_y.ctr\[29\]
rlabel metal2 7958 18020 7958 18020 0 dut.microstep_y.ctr\[2\]
rlabel metal2 8326 18428 8326 18428 0 dut.microstep_y.ctr\[3\]
rlabel metal2 7774 20604 7774 20604 0 dut.microstep_y.ctr\[4\]
rlabel metal1 8280 20570 8280 20570 0 dut.microstep_y.ctr\[5\]
rlabel metal1 9108 23698 9108 23698 0 dut.microstep_y.ctr\[6\]
rlabel metal2 9246 23494 9246 23494 0 dut.microstep_y.ctr\[7\]
rlabel metal2 12098 25024 12098 25024 0 dut.microstep_y.ctr\[8\]
rlabel metal1 12052 25874 12052 25874 0 dut.microstep_y.ctr\[9\]
rlabel metal1 24472 15130 24472 15130 0 dut.pid_x.x_pid.last_error\[1\]
rlabel metal1 23598 13260 23598 13260 0 dut.pid_x.x_pid.last_error\[2\]
rlabel metal2 24702 14552 24702 14552 0 dut.pid_x.x_pid.last_error\[3\]
rlabel metal1 25944 16218 25944 16218 0 dut.pid_y.y_pid.last_error\[1\]
rlabel metal2 24058 16320 24058 16320 0 dut.pid_y.y_pid.last_error\[2\]
rlabel metal1 23644 17714 23644 17714 0 dut.pid_y.y_pid.last_error\[3\]
rlabel metal1 27508 14926 27508 14926 0 dut.pwm_a_inst_x.count_d\[0\]
rlabel metal1 37069 6970 37069 6970 0 dut.pwm_a_inst_x.count_d\[10\]
rlabel metal1 35006 9928 35006 9928 0 dut.pwm_a_inst_x.count_d\[11\]
rlabel metal1 37122 10098 37122 10098 0 dut.pwm_a_inst_x.count_d\[12\]
rlabel metal2 36938 11356 36938 11356 0 dut.pwm_a_inst_x.count_d\[13\]
rlabel metal2 37030 13090 37030 13090 0 dut.pwm_a_inst_x.count_d\[14\]
rlabel metal1 36938 14450 36938 14450 0 dut.pwm_a_inst_x.count_d\[15\]
rlabel metal1 34868 13226 34868 13226 0 dut.pwm_a_inst_x.count_d\[16\]
rlabel metal1 35374 14586 35374 14586 0 dut.pwm_a_inst_x.count_d\[17\]
rlabel metal2 27002 15028 27002 15028 0 dut.pwm_a_inst_x.count_d\[1\]
rlabel metal1 27140 12410 27140 12410 0 dut.pwm_a_inst_x.count_d\[2\]
rlabel metal1 29440 12750 29440 12750 0 dut.pwm_a_inst_x.count_d\[3\]
rlabel metal1 29578 14314 29578 14314 0 dut.pwm_a_inst_x.count_d\[4\]
rlabel metal2 31234 14178 31234 14178 0 dut.pwm_a_inst_x.count_d\[5\]
rlabel metal2 31142 13090 31142 13090 0 dut.pwm_a_inst_x.count_d\[6\]
rlabel metal1 32844 13226 32844 13226 0 dut.pwm_a_inst_x.count_d\[7\]
rlabel metal1 33212 12614 33212 12614 0 dut.pwm_a_inst_x.count_d\[8\]
rlabel metal1 36846 8602 36846 8602 0 dut.pwm_a_inst_x.count_d\[9\]
rlabel metal2 28198 15266 28198 15266 0 dut.pwm_a_inst_x.count_q\[0\]
rlabel metal1 34592 10778 34592 10778 0 dut.pwm_a_inst_x.count_q\[10\]
rlabel metal1 34960 9554 34960 9554 0 dut.pwm_a_inst_x.count_q\[11\]
rlabel metal1 35512 7854 35512 7854 0 dut.pwm_a_inst_x.count_q\[12\]
rlabel metal1 36156 7718 36156 7718 0 dut.pwm_a_inst_x.count_q\[13\]
rlabel metal1 38226 12818 38226 12818 0 dut.pwm_a_inst_x.count_q\[14\]
rlabel metal1 38548 13906 38548 13906 0 dut.pwm_a_inst_x.count_q\[15\]
rlabel metal1 36248 13498 36248 13498 0 dut.pwm_a_inst_x.count_q\[16\]
rlabel metal2 37306 15130 37306 15130 0 dut.pwm_a_inst_x.count_q\[17\]
rlabel metal2 34730 14892 34730 14892 0 dut.pwm_a_inst_x.count_q\[18\]
rlabel metal1 34776 14518 34776 14518 0 dut.pwm_a_inst_x.count_q\[19\]
rlabel metal1 28520 13906 28520 13906 0 dut.pwm_a_inst_x.count_q\[1\]
rlabel metal1 28566 13260 28566 13260 0 dut.pwm_a_inst_x.count_q\[2\]
rlabel metal1 28750 12954 28750 12954 0 dut.pwm_a_inst_x.count_q\[3\]
rlabel metal2 32982 10914 32982 10914 0 dut.pwm_a_inst_x.count_q\[4\]
rlabel metal2 30774 13600 30774 13600 0 dut.pwm_a_inst_x.count_q\[5\]
rlabel metal2 33258 10778 33258 10778 0 dut.pwm_a_inst_x.count_q\[6\]
rlabel metal1 33902 13906 33902 13906 0 dut.pwm_a_inst_x.count_q\[7\]
rlabel metal2 32798 11900 32798 11900 0 dut.pwm_a_inst_x.count_q\[8\]
rlabel metal2 36754 9316 36754 9316 0 dut.pwm_a_inst_x.count_q\[9\]
rlabel metal1 37398 7514 37398 7514 0 dut.pwm_a_inst_x.pwm_out
rlabel metal1 24840 23018 24840 23018 0 dut.pwm_a_inst_y.count_d\[0\]
rlabel metal1 33626 27642 33626 27642 0 dut.pwm_a_inst_y.count_d\[10\]
rlabel metal1 35006 29512 35006 29512 0 dut.pwm_a_inst_y.count_d\[11\]
rlabel metal1 34592 30090 34592 30090 0 dut.pwm_a_inst_y.count_d\[12\]
rlabel metal1 35466 30634 35466 30634 0 dut.pwm_a_inst_y.count_d\[13\]
rlabel metal1 34776 33014 34776 33014 0 dut.pwm_a_inst_y.count_d\[14\]
rlabel metal2 33534 33252 33534 33252 0 dut.pwm_a_inst_y.count_d\[15\]
rlabel metal2 32154 32674 32154 32674 0 dut.pwm_a_inst_y.count_d\[16\]
rlabel metal2 30682 32028 30682 32028 0 dut.pwm_a_inst_y.count_d\[17\]
rlabel metal1 23598 23222 23598 23222 0 dut.pwm_a_inst_y.count_d\[1\]
rlabel metal2 24794 24990 24794 24990 0 dut.pwm_a_inst_y.count_d\[2\]
rlabel metal1 26450 25160 26450 25160 0 dut.pwm_a_inst_y.count_d\[3\]
rlabel metal1 28382 25976 28382 25976 0 dut.pwm_a_inst_y.count_d\[4\]
rlabel metal1 28474 27030 28474 27030 0 dut.pwm_a_inst_y.count_d\[5\]
rlabel metal2 28290 28254 28290 28254 0 dut.pwm_a_inst_y.count_d\[6\]
rlabel metal2 28566 29478 28566 29478 0 dut.pwm_a_inst_y.count_d\[7\]
rlabel metal1 30452 29206 30452 29206 0 dut.pwm_a_inst_y.count_d\[8\]
rlabel metal1 34868 26894 34868 26894 0 dut.pwm_a_inst_y.count_d\[9\]
rlabel via2 26450 23069 26450 23069 0 dut.pwm_a_inst_y.count_q\[0\]
rlabel metal1 35190 28424 35190 28424 0 dut.pwm_a_inst_y.count_q\[10\]
rlabel metal2 36478 29036 36478 29036 0 dut.pwm_a_inst_y.count_q\[11\]
rlabel metal1 36432 31790 36432 31790 0 dut.pwm_a_inst_y.count_q\[12\]
rlabel metal1 37076 29478 37076 29478 0 dut.pwm_a_inst_y.count_q\[13\]
rlabel metal1 36708 32742 36708 32742 0 dut.pwm_a_inst_y.count_q\[14\]
rlabel metal1 35328 33422 35328 33422 0 dut.pwm_a_inst_y.count_q\[15\]
rlabel metal1 33442 32402 33442 32402 0 dut.pwm_a_inst_y.count_q\[16\]
rlabel metal1 32614 31790 32614 31790 0 dut.pwm_a_inst_y.count_q\[17\]
rlabel metal2 32154 30430 32154 30430 0 dut.pwm_a_inst_y.count_q\[18\]
rlabel metal1 32476 30090 32476 30090 0 dut.pwm_a_inst_y.count_q\[19\]
rlabel metal1 26542 22576 26542 22576 0 dut.pwm_a_inst_y.count_q\[1\]
rlabel metal1 27094 24106 27094 24106 0 dut.pwm_a_inst_y.count_q\[2\]
rlabel metal2 27462 24956 27462 24956 0 dut.pwm_a_inst_y.count_q\[3\]
rlabel metal1 31993 26962 31993 26962 0 dut.pwm_a_inst_y.count_q\[4\]
rlabel metal2 31786 27268 31786 27268 0 dut.pwm_a_inst_y.count_q\[5\]
rlabel metal1 29992 28594 29992 28594 0 dut.pwm_a_inst_y.count_q\[6\]
rlabel metal1 29670 29614 29670 29614 0 dut.pwm_a_inst_y.count_q\[7\]
rlabel metal2 31878 27846 31878 27846 0 dut.pwm_a_inst_y.count_q\[8\]
rlabel viali 34998 28458 34998 28458 0 dut.pwm_a_inst_y.count_q\[9\]
rlabel metal2 38042 28220 38042 28220 0 dut.pwm_a_inst_y.pwm_out
rlabel metal1 27554 36346 27554 36346 0 dut.sclk_lcd
rlabel metal1 25484 34034 25484 34034 0 dut.sdo_lcd
rlabel metal1 27554 32878 27554 32878 0 dut.spi.bit_counter_q\[0\]
rlabel metal1 27968 32810 27968 32810 0 dut.spi.bit_counter_q\[1\]
rlabel metal2 28750 33184 28750 33184 0 dut.spi.bit_counter_q\[2\]
rlabel metal1 29118 34612 29118 34612 0 dut.spi.bit_counter_q\[3\]
rlabel metal2 28382 36516 28382 36516 0 dut.spi.clk_counter_d\[0\]
rlabel metal2 29394 36516 29394 36516 0 dut.spi.clk_counter_d\[1\]
rlabel metal1 31878 34476 31878 34476 0 dut.spi.clk_counter_d\[2\]
rlabel metal1 30682 35802 30682 35802 0 dut.spi.clk_counter_d\[3\]
rlabel metal2 31786 34340 31786 34340 0 dut.spi.clk_counter_d\[4\]
rlabel metal1 29854 34068 29854 34068 0 dut.spi.clk_counter_d\[5\]
rlabel metal1 28750 36176 28750 36176 0 dut.spi.clk_counter_q\[0\]
rlabel metal1 29210 36142 29210 36142 0 dut.spi.clk_counter_q\[1\]
rlabel metal2 32430 34918 32430 34918 0 dut.spi.clk_counter_q\[2\]
rlabel metal2 32246 35802 32246 35802 0 dut.spi.clk_counter_q\[3\]
rlabel metal1 30590 34578 30590 34578 0 dut.spi.clk_counter_q\[4\]
rlabel metal1 29486 34578 29486 34578 0 dut.spi.clk_counter_q\[5\]
rlabel metal1 19734 33082 19734 33082 0 dut.spi.cs_low_counter_d\[0\]
rlabel metal2 21758 34374 21758 34374 0 dut.spi.cs_low_counter_d\[1\]
rlabel metal1 22264 33082 22264 33082 0 dut.spi.cs_low_counter_d\[2\]
rlabel metal1 20644 35258 20644 35258 0 dut.spi.cs_low_counter_d\[3\]
rlabel metal1 20194 36856 20194 36856 0 dut.spi.cs_low_counter_d\[4\]
rlabel metal1 19504 35802 19504 35802 0 dut.spi.cs_low_counter_d\[5\]
rlabel metal1 20700 33830 20700 33830 0 dut.spi.cs_low_counter_q\[0\]
rlabel metal1 20378 34578 20378 34578 0 dut.spi.cs_low_counter_q\[1\]
rlabel metal1 21942 34476 21942 34476 0 dut.spi.cs_low_counter_q\[2\]
rlabel metal2 22218 35700 22218 35700 0 dut.spi.cs_low_counter_q\[3\]
rlabel metal1 21252 36890 21252 36890 0 dut.spi.cs_low_counter_q\[4\]
rlabel metal2 21022 35802 21022 35802 0 dut.spi.cs_low_counter_q\[5\]
rlabel metal1 24656 31450 24656 31450 0 dut.spi.shift_reg_q\[0\]
rlabel via1 25438 30022 25438 30022 0 dut.spi.shift_reg_q\[1\]
rlabel metal1 24012 29002 24012 29002 0 dut.spi.shift_reg_q\[2\]
rlabel metal1 27094 26962 27094 26962 0 dut.spi.shift_reg_q\[3\]
rlabel metal1 26036 26554 26036 26554 0 dut.spi.shift_reg_q\[4\]
rlabel metal1 26082 27574 26082 27574 0 dut.spi.shift_reg_q\[5\]
rlabel metal1 25944 28730 25944 28730 0 dut.spi.shift_reg_q\[6\]
rlabel metal2 26082 30192 26082 30192 0 dut.spi.shift_reg_q\[7\]
rlabel metal1 25208 31790 25208 31790 0 dut.spi.shift_reg_q\[8\]
rlabel metal2 27646 35564 27646 35564 0 dut.spi.spi_clk_q
rlabel metal1 26312 36210 26312 36210 0 dut.spi.state_q\[0\]
rlabel metal2 23874 35088 23874 35088 0 dut.spi.state_q\[1\]
rlabel metal1 24012 36142 24012 36142 0 dut.spi.state_q\[2\]
rlabel metal1 1518 10234 1518 10234 0 en
rlabel metal2 14858 1520 14858 1520 0 gpio_in[6]
rlabel metal2 38410 27183 38410 27183 0 gpio_out[10]
rlabel metal1 23966 37094 23966 37094 0 gpio_out[11]
rlabel metal1 25944 37094 25944 37094 0 gpio_out[12]
rlabel metal1 26542 37094 26542 37094 0 gpio_out[13]
rlabel metal1 1426 24650 1426 24650 0 gpio_out[7]
rlabel metal2 21298 1520 21298 1520 0 gpio_out[8]
rlabel metal2 38410 7633 38410 7633 0 gpio_out[9]
rlabel metal1 1886 10676 1886 10676 0 net1
rlabel metal1 38180 7854 38180 7854 0 net10
rlabel metal1 29716 37434 29716 37434 0 net100
rlabel metal1 7176 2822 7176 2822 0 net101
rlabel metal3 751 5508 751 5508 0 net102
rlabel metal2 5198 1027 5198 1027 0 net103
rlabel via2 38502 35445 38502 35445 0 net104
rlabel metal2 38502 34221 38502 34221 0 net105
rlabel metal3 751 3468 751 3468 0 net106
rlabel metal3 751 29988 751 29988 0 net107
rlabel metal1 1518 37434 1518 37434 0 net108
rlabel metal1 35512 37434 35512 37434 0 net109
rlabel metal1 25300 11730 25300 11730 0 net11
rlabel via2 38502 33371 38502 33371 0 net110
rlabel metal3 751 29308 751 29308 0 net111
rlabel metal2 30314 1588 30314 1588 0 net112
rlabel via2 38502 30685 38502 30685 0 net113
rlabel via2 38226 37451 38226 37451 0 net114
rlabel metal1 36156 37434 36156 37434 0 net115
rlabel metal1 34224 37434 34224 37434 0 net116
rlabel metal3 751 36788 751 36788 0 net117
rlabel via2 38502 3485 38502 3485 0 net118
rlabel metal1 3312 37434 3312 37434 0 net119
rlabel metal1 19550 28118 19550 28118 0 net12
rlabel metal1 29072 37434 29072 37434 0 net120
rlabel metal2 37950 38131 37950 38131 0 net121
rlabel metal2 33166 15504 33166 15504 0 net122
rlabel metal1 32936 15402 32936 15402 0 net123
rlabel metal1 30452 30294 30452 30294 0 net124
rlabel metal2 29946 30872 29946 30872 0 net125
rlabel metal2 38502 15181 38502 15181 0 net126
rlabel metal2 38502 36941 38502 36941 0 net127
rlabel metal2 27738 1520 27738 1520 0 net128
rlabel metal2 27094 1520 27094 1520 0 net129
rlabel metal1 12650 31858 12650 31858 0 net13
rlabel metal3 751 2788 751 2788 0 net130
rlabel metal3 751 6868 751 6868 0 net131
rlabel metal3 751 6188 751 6188 0 net132
rlabel via2 38502 36091 38502 36091 0 net133
rlabel metal3 751 35428 751 35428 0 net134
rlabel metal3 751 4148 751 4148 0 net135
rlabel metal1 31648 37230 31648 37230 0 net136
rlabel metal1 5244 37230 5244 37230 0 net137
rlabel metal1 27140 37230 27140 37230 0 net138
rlabel metal1 33580 37230 33580 37230 0 net139
rlabel metal2 16330 34255 16330 34255 0 net14
rlabel metal2 38502 2193 38502 2193 0 net140
rlabel metal1 28428 37230 28428 37230 0 net141
rlabel metal1 30360 37230 30360 37230 0 net142
rlabel metal2 38502 34833 38502 34833 0 net143
rlabel metal3 751 4828 751 4828 0 net144
rlabel metal3 751 28628 751 28628 0 net145
rlabel metal1 31004 37230 31004 37230 0 net146
rlabel metal1 32936 37230 32936 37230 0 net147
rlabel metal3 820 9588 820 9588 0 net148
rlabel metal2 38502 2873 38502 2873 0 net149
rlabel metal1 13018 5168 13018 5168 0 net15
rlabel metal2 29026 1520 29026 1520 0 net150
rlabel metal2 24518 1520 24518 1520 0 net151
rlabel metal1 32292 37230 32292 37230 0 net152
rlabel metal1 7912 35054 7912 35054 0 net153
rlabel metal1 17250 13940 17250 13940 0 net154
rlabel metal2 2990 11458 2990 11458 0 net155
rlabel metal1 7682 13362 7682 13362 0 net156
rlabel metal1 8372 16966 8372 16966 0 net157
rlabel metal1 23690 25262 23690 25262 0 net158
rlabel metal1 23092 28526 23092 28526 0 net159
rlabel metal1 10580 3502 10580 3502 0 net16
rlabel metal1 23828 24174 23828 24174 0 net160
rlabel metal1 24334 30770 24334 30770 0 net161
rlabel metal1 23138 31654 23138 31654 0 net162
rlabel metal2 11270 9758 11270 9758 0 net163
rlabel metal2 9706 9418 9706 9418 0 net164
rlabel metal1 24288 14586 24288 14586 0 net165
rlabel metal1 7084 20434 7084 20434 0 net166
rlabel metal1 9384 10030 9384 10030 0 net167
rlabel metal2 22218 31484 22218 31484 0 net168
rlabel metal1 5796 12138 5796 12138 0 net169
rlabel metal1 6532 21522 6532 21522 0 net17
rlabel metal1 6440 11118 6440 11118 0 net170
rlabel metal1 7360 17578 7360 17578 0 net171
rlabel metal2 8786 18054 8786 18054 0 net172
rlabel metal1 26266 15470 26266 15470 0 net173
rlabel metal2 7958 21114 7958 21114 0 net174
rlabel metal1 7590 20876 7590 20876 0 net175
rlabel metal1 4508 19346 4508 19346 0 net176
rlabel metal1 25668 31994 25668 31994 0 net177
rlabel metal2 27002 31042 27002 31042 0 net178
rlabel metal1 8510 13226 8510 13226 0 net179
rlabel metal1 16606 23154 16606 23154 0 net18
rlabel metal1 8648 12614 8648 12614 0 net180
rlabel metal1 8924 18394 8924 18394 0 net181
rlabel metal1 2530 11084 2530 11084 0 net182
rlabel metal1 9614 30260 9614 30260 0 net183
rlabel metal1 28566 36108 28566 36108 0 net184
rlabel metal1 7958 29478 7958 29478 0 net185
rlabel metal1 7728 9622 7728 9622 0 net186
rlabel metal2 21850 27268 21850 27268 0 net187
rlabel metal1 7498 11118 7498 11118 0 net188
rlabel metal2 11730 34782 11730 34782 0 net189
rlabel metal1 21666 27370 21666 27370 0 net19
rlabel metal1 7958 9996 7958 9996 0 net190
rlabel metal2 11362 16796 11362 16796 0 net191
rlabel via1 25070 32402 25070 32402 0 net192
rlabel metal1 20010 12750 20010 12750 0 net193
rlabel metal1 2162 24752 2162 24752 0 net194
rlabel metal1 2852 6290 2852 6290 0 net195
rlabel metal1 2576 26962 2576 26962 0 net196
rlabel metal2 31694 34816 31694 34816 0 net197
rlabel metal2 6854 36618 6854 36618 0 net198
rlabel metal1 18538 16082 18538 16082 0 net199
rlabel metal1 15042 2618 15042 2618 0 net2
rlabel metal1 26818 31892 26818 31892 0 net20
rlabel metal1 14996 31790 14996 31790 0 net200
rlabel metal2 3266 35258 3266 35258 0 net201
rlabel metal1 14536 29818 14536 29818 0 net202
rlabel metal1 7452 31314 7452 31314 0 net203
rlabel metal1 5060 33490 5060 33490 0 net204
rlabel metal1 4876 31790 4876 31790 0 net205
rlabel metal1 3450 3094 3450 3094 0 net206
rlabel metal2 4646 30940 4646 30940 0 net207
rlabel metal2 5566 35938 5566 35938 0 net208
rlabel metal1 4278 35088 4278 35088 0 net209
rlabel metal1 30820 32334 30820 32334 0 net21
rlabel metal1 20424 17102 20424 17102 0 net210
rlabel metal1 3818 33966 3818 33966 0 net211
rlabel metal1 5152 29614 5152 29614 0 net212
rlabel metal2 8970 36550 8970 36550 0 net213
rlabel metal1 8004 36142 8004 36142 0 net214
rlabel metal1 5888 9554 5888 9554 0 net215
rlabel metal1 26358 26860 26358 26860 0 net216
rlabel metal1 27186 26282 27186 26282 0 net217
rlabel metal1 14582 30770 14582 30770 0 net218
rlabel metal1 25760 28050 25760 28050 0 net219
rlabel metal1 33672 32946 33672 32946 0 net22
rlabel metal1 27471 27642 27471 27642 0 net220
rlabel metal1 37674 10710 37674 10710 0 net221
rlabel metal2 24886 26554 24886 26554 0 net222
rlabel metal1 24334 26894 24334 26894 0 net223
rlabel metal1 5382 28152 5382 28152 0 net224
rlabel metal1 35144 31790 35144 31790 0 net225
rlabel metal1 9890 32946 9890 32946 0 net226
rlabel metal1 10672 31722 10672 31722 0 net227
rlabel metal1 25760 29682 25760 29682 0 net228
rlabel metal2 27554 29852 27554 29852 0 net229
rlabel metal1 2760 24786 2760 24786 0 net23
rlabel viali 4646 36143 4646 36143 0 net230
rlabel metal1 20010 34544 20010 34544 0 net231
rlabel metal1 20194 33592 20194 33592 0 net232
rlabel metal1 6394 8466 6394 8466 0 net233
rlabel metal1 16008 18938 16008 18938 0 net234
rlabel metal1 2898 17612 2898 17612 0 net235
rlabel metal1 34178 32742 34178 32742 0 net236
rlabel metal1 29164 29546 29164 29546 0 net237
rlabel metal2 4738 28288 4738 28288 0 net238
rlabel metal1 4968 6358 4968 6358 0 net239
rlabel metal2 3818 21012 3818 21012 0 net24
rlabel metal1 27646 14042 27646 14042 0 net240
rlabel metal1 27416 14450 27416 14450 0 net241
rlabel metal1 25530 28084 25530 28084 0 net242
rlabel metal1 27738 28594 27738 28594 0 net243
rlabel metal1 2438 19346 2438 19346 0 net244
rlabel metal1 10350 25874 10350 25874 0 net245
rlabel metal1 24794 28050 24794 28050 0 net246
rlabel metal1 25530 29206 25530 29206 0 net247
rlabel metal2 16882 20672 16882 20672 0 net248
rlabel metal1 5842 24106 5842 24106 0 net249
rlabel metal2 36202 8092 36202 8092 0 net25
rlabel metal1 15548 32878 15548 32878 0 net250
rlabel metal2 11546 29410 11546 29410 0 net251
rlabel metal1 24334 30158 24334 30158 0 net252
rlabel metal1 11500 30226 11500 30226 0 net253
rlabel metal1 4738 4590 4738 4590 0 net254
rlabel metal1 6118 3060 6118 3060 0 net255
rlabel metal1 13064 5678 13064 5678 0 net256
rlabel metal1 4784 23018 4784 23018 0 net257
rlabel metal1 9706 3366 9706 3366 0 net258
rlabel metal1 9522 29104 9522 29104 0 net259
rlabel metal1 35098 13974 35098 13974 0 net26
rlabel metal1 10580 28050 10580 28050 0 net260
rlabel metal1 9798 25976 9798 25976 0 net261
rlabel metal1 8786 2618 8786 2618 0 net262
rlabel metal1 6072 4590 6072 4590 0 net263
rlabel metal2 3266 14620 3266 14620 0 net264
rlabel metal1 5980 13906 5980 13906 0 net265
rlabel metal1 3266 24208 3266 24208 0 net266
rlabel metal1 5244 18258 5244 18258 0 net267
rlabel metal1 3680 24174 3680 24174 0 net268
rlabel metal1 7406 25806 7406 25806 0 net269
rlabel metal2 31786 13294 31786 13294 0 net27
rlabel metal1 13156 5202 13156 5202 0 net270
rlabel metal1 6210 25942 6210 25942 0 net271
rlabel metal1 10074 7888 10074 7888 0 net272
rlabel metal1 8648 21998 8648 21998 0 net273
rlabel metal1 16974 21522 16974 21522 0 net274
rlabel metal1 4048 5678 4048 5678 0 net275
rlabel metal2 5566 16524 5566 16524 0 net276
rlabel metal1 22632 17306 22632 17306 0 net277
rlabel metal1 11224 3706 11224 3706 0 net278
rlabel metal2 4278 29308 4278 29308 0 net279
rlabel metal1 17549 18326 17549 18326 0 net28
rlabel metal2 2806 26741 2806 26741 0 net280
rlabel metal1 2714 13294 2714 13294 0 net281
rlabel metal1 28060 32402 28060 32402 0 net282
rlabel metal1 37490 14042 37490 14042 0 net283
rlabel metal1 21620 7378 21620 7378 0 net284
rlabel metal2 4830 7548 4830 7548 0 net285
rlabel metal2 11638 21046 11638 21046 0 net286
rlabel metal1 3910 19414 3910 19414 0 net287
rlabel metal1 18492 33898 18492 33898 0 net288
rlabel metal2 30774 33082 30774 33082 0 net289
rlabel via1 17074 18666 17074 18666 0 net29
rlabel metal1 30590 33558 30590 33558 0 net290
rlabel metal1 13938 34986 13938 34986 0 net291
rlabel metal2 2898 16592 2898 16592 0 net292
rlabel metal1 33028 31790 33028 31790 0 net293
rlabel metal1 27830 33456 27830 33456 0 net294
rlabel metal1 2576 14314 2576 14314 0 net295
rlabel metal2 11730 31484 11730 31484 0 net296
rlabel metal2 21574 13124 21574 13124 0 net297
rlabel metal1 18538 14246 18538 14246 0 net298
rlabel metal2 18814 14620 18814 14620 0 net299
rlabel metal1 1656 10642 1656 10642 0 net3
rlabel metal1 14306 18190 14306 18190 0 net30
rlabel metal1 11362 33456 11362 33456 0 net300
rlabel metal1 17020 20842 17020 20842 0 net301
rlabel metal2 16054 34748 16054 34748 0 net302
rlabel metal1 33350 14042 33350 14042 0 net303
rlabel metal1 8970 26350 8970 26350 0 net304
rlabel metal1 11316 24786 11316 24786 0 net305
rlabel metal1 13754 6290 13754 6290 0 net306
rlabel metal1 15410 8602 15410 8602 0 net307
rlabel metal1 13616 9690 13616 9690 0 net308
rlabel metal1 7866 6222 7866 6222 0 net309
rlabel metal2 14766 13804 14766 13804 0 net31
rlabel metal1 14674 15130 14674 15130 0 net310
rlabel metal1 14214 12342 14214 12342 0 net311
rlabel metal1 16376 30702 16376 30702 0 net312
rlabel metal2 36662 15164 36662 15164 0 net313
rlabel metal1 12098 3570 12098 3570 0 net314
rlabel metal1 12834 19278 12834 19278 0 net315
rlabel metal1 17664 18258 17664 18258 0 net316
rlabel metal1 12926 13328 12926 13328 0 net317
rlabel metal1 24334 22950 24334 22950 0 net318
rlabel metal1 12972 22406 12972 22406 0 net319
rlabel metal1 18860 13906 18860 13906 0 net32
rlabel metal2 12006 17680 12006 17680 0 net320
rlabel metal1 10304 13906 10304 13906 0 net321
rlabel metal1 4830 32538 4830 32538 0 net322
rlabel metal2 13478 20060 13478 20060 0 net323
rlabel metal1 13616 17714 13616 17714 0 net33
rlabel metal1 18446 16966 18446 16966 0 net34
rlabel metal2 20010 14926 20010 14926 0 net35
rlabel metal1 37950 20842 37950 20842 0 net36
rlabel metal1 36478 19346 36478 19346 0 net37
rlabel metal1 37582 19278 37582 19278 0 net38
rlabel metal1 32062 16592 32062 16592 0 net39
rlabel metal2 38226 27404 38226 27404 0 net4
rlabel metal1 34776 19142 34776 19142 0 net40
rlabel metal1 36386 19924 36386 19924 0 net41
rlabel metal1 26680 21522 26680 21522 0 net42
rlabel metal1 15916 28186 15916 28186 0 net43
rlabel metal1 33212 18190 33212 18190 0 net44
rlabel metal1 34960 4590 34960 4590 0 net45
rlabel metal1 30866 4046 30866 4046 0 net46
rlabel metal2 28198 3434 28198 3434 0 net47
rlabel metal2 22034 5814 22034 5814 0 net48
rlabel metal2 27462 4046 27462 4046 0 net49
rlabel metal2 24242 37060 24242 37060 0 net5
rlabel metal2 3910 11356 3910 11356 0 net50
rlabel metal1 8839 3094 8839 3094 0 net51
rlabel metal1 5789 7786 5789 7786 0 net52
rlabel metal2 2714 16524 2714 16524 0 net53
rlabel metal1 7459 14314 7459 14314 0 net54
rlabel metal2 10442 18156 10442 18156 0 net55
rlabel metal1 5159 16082 5159 16082 0 net56
rlabel metal2 12558 3842 12558 3842 0 net57
rlabel metal1 19097 7446 19097 7446 0 net58
rlabel metal2 15502 16558 15502 16558 0 net59
rlabel metal1 25806 37230 25806 37230 0 net6
rlabel metal2 16146 18802 16146 18802 0 net60
rlabel metal2 20010 16439 20010 16439 0 net61
rlabel metal2 5014 19992 5014 19992 0 net62
rlabel metal1 9913 27030 9913 27030 0 net63
rlabel metal2 5750 35938 5750 35938 0 net64
rlabel via1 8142 33507 8142 33507 0 net65
rlabel metal2 7038 32623 7038 32623 0 net66
rlabel metal1 9023 20502 9023 20502 0 net67
rlabel metal1 16199 21590 16199 21590 0 net68
rlabel metal2 20010 34986 20010 34986 0 net69
rlabel metal2 27002 37060 27002 37060 0 net7
rlabel metal2 14950 33558 14950 33558 0 net70
rlabel metal1 19366 20774 19366 20774 0 net71
rlabel metal1 3956 21522 3956 21522 0 net72
rlabel metal2 20838 19074 20838 19074 0 net73
rlabel metal2 28014 16252 28014 16252 0 net74
rlabel metal2 21666 13090 21666 13090 0 net75
rlabel metal2 37490 12138 37490 12138 0 net76
rlabel metal1 35243 16490 35243 16490 0 net77
rlabel metal2 37490 7735 37490 7735 0 net78
rlabel metal2 20378 20910 20378 20910 0 net79
rlabel metal1 1702 24718 1702 24718 0 net8
rlabel metal2 25530 20672 25530 20672 0 net80
rlabel metal2 21390 35836 21390 35836 0 net81
rlabel metal1 27370 36822 27370 36822 0 net82
rlabel metal2 21114 29750 21114 29750 0 net83
rlabel metal1 31786 31831 31786 31831 0 net84
rlabel metal1 35151 33558 35151 33558 0 net85
rlabel metal2 32982 27574 32982 27574 0 net86
rlabel metal2 22034 20417 22034 20417 0 net87
rlabel metal1 27784 37434 27784 37434 0 net88
rlabel metal2 23874 1588 23874 1588 0 net89
rlabel metal2 21390 2587 21390 2587 0 net9
rlabel metal2 36110 1588 36110 1588 0 net90
rlabel metal2 35466 1588 35466 1588 0 net91
rlabel metal3 751 36108 751 36108 0 net92
rlabel metal1 38548 36754 38548 36754 0 net93
rlabel metal3 38878 31348 38878 31348 0 net94
rlabel metal3 751 34748 751 34748 0 net95
rlabel metal1 36800 37434 36800 37434 0 net96
rlabel metal1 34868 37434 34868 37434 0 net97
rlabel metal2 29670 1588 29670 1588 0 net98
rlabel metal1 38272 36754 38272 36754 0 net99
rlabel metal1 1380 11118 1380 11118 0 nrst
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
