* NGSPICE file created from team_07.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_40_12 abstract view
.subckt sky130_ef_sc_hd__decap_40_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_4 abstract view
.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_8 abstract view
.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_07 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
X_05903_ top0.CPU.register.registers\[770\] top0.CPU.register.registers\[802\] top0.CPU.register.registers\[834\]
+ top0.CPU.register.registers\[866\] net831 net796 vssd1 vssd1 vccd1 vccd1 _02560_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08731__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06883_ net860 _03531_ _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__a21oi_4
X_09671_ net768 _05186_ net651 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06968__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05834_ _02489_ _02490_ net729 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
X_08622_ net714 net214 net310 net330 net2495 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__a32o_1
XFILLER_55_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05765_ _02384_ net632 net626 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nand3_2
XFILLER_70_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08553_ net153 net678 net397 net362 net2272 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__a32o_1
XANTENNA__07332__B _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _02769_ net527 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ net160 net614 net386 net369 net2659 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a32o_1
XANTENNA__05848__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05696_ top0.MMIO.WBData_i\[18\] vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__inv_2
XANTENNA__07837__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07435_ net469 _03403_ _03820_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a21bo_1
X_11299__951 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__inv_2
XANTENNA_fanout427_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05943__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07366_ _03918_ _03922_ net456 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__mux2_1
XANTENNA__08798__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06317_ top0.CPU.register.registers\[412\] top0.CPU.register.registers\[444\] top0.CPU.register.registers\[476\]
+ top0.CPU.register.registers\[508\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02974_
+ sky130_fd_sc_hd__mux4_1
X_09105_ top0.CPU.register.registers\[88\] net568 vssd1 vssd1 vccd1 vccd1 _04827_
+ sky130_fd_sc_hd__or2_1
X_07297_ net489 _03953_ _03755_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_98_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09036_ net217 net613 _04805_ net351 net3216 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__a32o_1
X_06248_ _02901_ _02904_ net780 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
XANTENNA__08163__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout796_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold362 top0.CPU.register.registers\[872\] vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold351 top0.CPU.register.registers\[117\] vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ top0.CPU.register.registers\[533\] top0.CPU.register.registers\[565\] top0.CPU.register.registers\[597\]
+ top0.CPU.register.registers\[629\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02836_
+ sky130_fd_sc_hd__mux4_1
Xhold340 top0.CPU.register.registers\[962\] vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 top0.CPU.register.registers\[932\] vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 top0.CPU.register.registers\[374\] vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 top0.CPU.register.registers\[635\] vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout820 net822 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_4
X_09938_ top0.CPU.internalMem.pcOut\[23\] _05421_ _05410_ vssd1 vssd1 vccd1 vccd1
+ _05432_ sky130_fd_sc_hd__a21o_1
Xfanout842 net844 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_4
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 net834 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_4
X_10556__208 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__inv_2
Xfanout864 net868 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_4
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_2
XFILLER_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 top0.CPU.register.registers\[77\] vssd1 vssd1 vccd1 vccd1 net3273 sky130_fd_sc_hd__dlygate4sd3_1
X_09869_ top0.CPU.internalMem.pcOut\[18\] _05359_ vssd1 vssd1 vccd1 vccd1 _05369_
+ sky130_fd_sc_hd__nand2_1
Xfanout897 net904 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_51_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 top0.CPU.register.registers\[90\] vssd1 vssd1 vccd1 vccd1 net3262 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout886 net887 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06959__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11900_ net1592 _01539_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[393\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1084 top0.CPU.register.registers\[197\] vssd1 vssd1 vccd1 vccd1 net3306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1073 top0.CPU.register.registers\[264\] vssd1 vssd1 vccd1 vccd1 net3295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 top0.CPU.register.registers\[107\] vssd1 vssd1 vccd1 vccd1 net3284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11831_ net1523 _01470_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[324\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1095 top0.CPU.register.registers\[130\] vssd1 vssd1 vccd1 vccd1 net3317 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07242__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ net1454 _01401_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[255\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11693_ net1385 _01332_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08354__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12314_ net2006 _01953_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[807\]
+ sky130_fd_sc_hd__dfrtp_1
X_11092__744 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__inv_2
XANTENNA__10108__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ net1937 _01884_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[738\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06435__A1_N net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ net1868 _01815_ net1081 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[669\]
+ sky130_fd_sc_hd__dfrtp_1
X_11133__785 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__inv_2
XANTENNA__08961__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10124__A _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08713__A0 _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05870__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10009_ top0.CPU.internalMem.pcOut\[29\] _05496_ vssd1 vssd1 vccd1 vccd1 _05498_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_82_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06178__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08492__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ net455 _03726_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__or2_1
X_10997__649 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__inv_2
X_07151_ net532 _03403_ net472 vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__mux2_1
XFILLER_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06102_ top0.CPU.register.registers\[140\] top0.CPU.register.registers\[172\] top0.CPU.register.registers\[204\]
+ top0.CPU.register.registers\[236\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02759_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08244__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09633__B1_N _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10018__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741__393 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__inv_2
X_07082_ _03713_ _03737_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__or2_1
XANTENNA__08795__A3 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06033_ top0.CPU.register.registers\[521\] top0.CPU.register.registers\[553\] top0.CPU.register.registers\[585\]
+ top0.CPU.register.registers\[617\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02690_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08547__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06102__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout138 net140 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
Xfanout127 net128 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08952__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout116 _05643_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_93_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07984_ top0.CPU.internalMem.pcOut\[5\] net640 _04613_ _04614_ net635 vssd1 vssd1
+ vccd1 vccd1 _04615_ sky130_fd_sc_hd__o221a_4
Xfanout149 _05012_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_2
X_09723_ top0.CPU.internalMem.pcOut\[7\] _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__nand2_1
X_06935_ net863 _03587_ net858 vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__o21ai_1
X_09654_ net3379 top0.MISOtoMMIO\[5\] _05173_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux2_1
X_06866_ _02618_ _02685_ _02716_ net542 vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a31o_1
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout377_A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08180__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05817_ _02380_ _02447_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__nand2_2
X_08605_ net2952 net330 net315 _04540_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a22o_1
X_06797_ _03452_ _03453_ net873 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux2_1
X_09585_ top0.display.counter\[2\] _05122_ _05124_ top0.display.counter\[3\] vssd1
+ vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05748_ net545 _02404_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__nor2_1
X_08536_ _04718_ net388 net361 net2702 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ _04684_ net407 net372 net2767 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05679_ net769 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08483__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07418_ net450 _03755_ _03927_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_21_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08398_ _04663_ net396 net378 net2827 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07349_ _03740_ _04003_ _04004_ net443 _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1163 vssd1 vssd1 vccd1 vccd1 team_07_1163/HI gpio_out[29] sky130_fd_sc_hd__conb_1
X_11076__728 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__inv_2
X_10436__88 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__inv_2
Xteam_07_1141 vssd1 vssd1 vccd1 vccd1 team_07_1141/HI gpio_out[7] sky130_fd_sc_hd__conb_1
Xteam_07_1152 vssd1 vssd1 vccd1 vccd1 team_07_1152/HI gpio_out[18] sky130_fd_sc_hd__conb_1
XFILLER_12_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xteam_07_1185 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] team_07_1185/LO sky130_fd_sc_hd__conb_1
Xteam_07_1174 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] team_07_1174/LO sky130_fd_sc_hd__conb_1
Xteam_07_1196 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] team_07_1196/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ _04938_ _05594_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__or2_1
XANTENNA__07780__A1_N _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ net205 net2992 net350 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
XANTENNA__07994__A1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117__769 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__inv_2
Xhold170 top0.CPU.register.registers\[175\] vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
X_12030_ net1722 _01669_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[523\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08113__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 top0.CPU.register.registers\[818\] vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 top0.CPU.register.registers\[747\] vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05852__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_4
Xfanout672 net673 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_4
Xfanout661 _04954_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_2
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08171__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08068__B net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ net1506 _01453_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08474__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10684__336 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__inv_2
X_11745_ net1437 _01384_ net1059 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05907__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06485__A1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08084__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11676_ net1368 _01315_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[169\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06580__S1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10725__377 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__B _02729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12228_ net1920 _01867_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[721\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08934__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10578__230 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ net1851 _01798_ net1101 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619__271 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__inv_2
XFILLER_77_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12596__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ _03373_ _03374_ _03375_ _03376_ net757 net862 vssd1 vssd1 vccd1 vccd1 _03377_
+ sky130_fd_sc_hd__mux4_1
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06651_ _03304_ _03305_ _03306_ _03307_ net756 net749 vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__mux4_1
XFILLER_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06582_ net871 _03236_ net752 vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a21o_1
X_09370_ net2822 _04568_ net606 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08321_ net545 _02403_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor2_1
XANTENNA__09111__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06020__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ net2756 net417 _04711_ net491 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a22o_1
X_07203_ net457 _03859_ _03831_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08217__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_08183_ net504 net174 net620 net427 net2346 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_95_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07134_ net447 net536 net475 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__mux2_1
XANTENNA__06941__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11407__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ _03403_ _03262_ net468 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__mux2_1
XANTENNA__09029__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06016_ net784 _02672_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout494_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06087__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07967_ _04069_ net232 net227 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ top0.CPU.control.funct7\[1\] net631 _02453_ vssd1 vssd1 vccd1 vccd1 _05218_
+ sky130_fd_sc_hd__and3_1
X_06918_ _03177_ _03198_ _03572_ _03574_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout759_A _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ top0.CPU.internalMem.pcOut\[20\] net638 net633 _04543_ vssd1 vssd1 vccd1
+ vccd1 _04544_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06164__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ net142 _05164_ net660 vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a21oi_1
X_06849_ _02619_ _02686_ _02718_ net540 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout926_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09568_ _04292_ net233 net228 net632 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_104_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ net154 net682 net397 net366 net2667 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a32o_1
XANTENNA__08456__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ top0.MMIO.WBData_i\[28\] net137 vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__or2_1
XANTENNA__06011__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ net1222 _01169_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ clknet_leaf_70_clk _01109_ net1117 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09405__A1 top0.MMIO.WBData_i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11392_ clknet_leaf_59_clk _01040_ net1091 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08759__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ net2238 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06314__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net144 _05160_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nand2_1
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06078__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__A3 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net1705 _01652_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05745__A3 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout491 net496 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06298__S net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11245__897 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__inv_2
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12777_ top0.display.sclk vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
X_11098__750 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__inv_2
XANTENNA__08998__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11728_ net1420 _01367_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ net1351 _01298_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[152\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07407__A0 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold917 top0.CPU.register.registers\[659\] vssd1 vssd1 vccd1 vccd1 net3139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold906 top0.CPU.intMemAddr\[0\] vssd1 vssd1 vccd1 vccd1 net3128 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold928 top0.CPU.register.registers\[121\] vssd1 vssd1 vccd1 vccd1 net3150 sky130_fd_sc_hd__dlygate4sd3_1
X_11139__791 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__inv_2
Xhold939 top0.CPU.register.registers\[270\] vssd1 vssd1 vccd1 vccd1 net3161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06069__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_90_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__09175__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ net3010 net284 net275 _04493_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__a22o_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07821_ _04475_ net561 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__nor2_1
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07752_ _02635_ _03836_ _04053_ _03848_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_121_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08686__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ net450 _04267_ _03849_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a21o_1
X_06703_ _03357_ _03358_ _03339_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09422_ _04933_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__and2b_1
X_06634_ net869 _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__or2_1
XANTENNA__06792__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _02366_ _02367_ _04986_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.state_n\[3\]
+ sky130_fd_sc_hd__o21bai_1
X_08304_ net3148 _04571_ net415 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__mux2_1
X_06565_ net858 _03216_ _03220_ _03208_ _03212_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__o32ai_4
XFILLER_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10245__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09284_ _04942_ _04943_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__nand2_1
X_06496_ _03134_ _03150_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__xor2_1
XFILLER_21_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ net495 net166 net681 net421 net2586 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ net2986 net427 _04683_ net508 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
X_10406__58 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__inv_2
X_07117_ net454 _03719_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_132_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ net511 net181 net694 net434 net2338 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_132_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07048_ _03702_ _03703_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__or2_1
Xclkload90 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09166__A3 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__A3 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08999_ net214 net691 net271 net259 net2650 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__a32o_1
XANTENNA__07515__B _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__A1 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08677__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12700_ clknet_leaf_75_clk _02335_ net1124 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.storeCt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12631_ clknet_leaf_73_clk _02266_ net1127 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05896__C1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06783__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ clknet_leaf_55_clk _02201_ net1038 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_11513_ net1205 _01152_ net980 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12493_ net2185 _02132_ net958 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[986\]
+ sky130_fd_sc_hd__dfrtp_1
X_11444_ clknet_leaf_78_clk _01092_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.Op\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11375_ clknet_leaf_76_clk top0.CPU.internalMem.load2Ct_n\[1\] net1123 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.load2Ct\[1\] sky130_fd_sc_hd__dfrtp_1
X_10796__448 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__inv_2
XANTENNA__08601__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10326_ net2234 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__clkbuf_1
X_10540__192 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__inv_2
X_10420__72 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__inv_2
X_10257_ net3096 net118 net112 _05651_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a22o_1
XFILLER_78_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10837__489 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__inv_2
XANTENNA__09193__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05925__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ net609 _04930_ net149 vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08301__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07425__B _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08117__A1 _04528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08668__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06774__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05887__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06350_ net540 _03006_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__nand2_1
XANTENNA__07628__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06281_ top0.CPU.register.registers\[410\] top0.CPU.register.registers\[442\] top0.CPU.register.registers\[474\]
+ top0.CPU.register.registers\[506\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02938_
+ sky130_fd_sc_hd__mux4_1
XFILLER_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08020_ net210 net705 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__and2_1
XANTENNA__06491__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold703 top0.CPU.register.registers\[664\] vssd1 vssd1 vccd1 vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold714 top0.CPU.register.registers\[444\] vssd1 vssd1 vccd1 vccd1 net2936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 top0.CPU.register.registers\[782\] vssd1 vssd1 vccd1 vccd1 net2947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 top0.CPU.register.registers\[730\] vssd1 vssd1 vccd1 vccd1 net2958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold758 top0.CPU.intMem_out\[5\] vssd1 vssd1 vccd1 vccd1 net2980 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _05439_ _05449_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__nand2_1
Xhold769 top0.CPU.register.registers\[468\] vssd1 vssd1 vccd1 vccd1 net2991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 top0.CPU.register.registers\[512\] vssd1 vssd1 vccd1 vccd1 net2969 sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ _04641_ net552 _04774_ net263 net3343 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__a32o_1
XANTENNA__09553__A0 top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05835__S net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ net183 net3210 net356 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__mux2_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08784_ net191 net688 net327 net292 net2478 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a32o_1
XANTENNA__06462__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05996_ top0.CPU.register.registers\[519\] top0.CPU.register.registers\[551\] top0.CPU.register.registers\[583\]
+ top0.CPU.register.registers\[615\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02653_
+ sky130_fd_sc_hd__mux4_1
X_07804_ net537 net536 _03129_ net447 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__and4_1
XANTENNA__07903__X _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07735_ _03871_ _03879_ net345 vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__mux2_1
XFILLER_93_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout457_A _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__B1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ top0.MMIO.WBData_i\[1\] net147 net143 top0.MISOtoMMIO\[1\] _05014_ vssd1
+ vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__o221a_1
XFILLER_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07331__A2 _03504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ _03834_ _03838_ net517 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout624_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06617_ top0.CPU.register.registers\[261\] top0.CPU.register.registers\[293\] top0.CPU.register.registers\[325\]
+ top0.CPU.register.registers\[357\] net934 net900 vssd1 vssd1 vccd1 vccd1 _03274_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_101_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09608__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ net530 net531 net470 vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__mux2_1
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09336_ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__inv_2
XANTENNA__09084__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06548_ top0.CPU.register.registers\[657\] top0.CPU.register.registers\[689\] top0.CPU.register.registers\[721\]
+ top0.CPU.register.registers\[753\] net913 net879 vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__mux4_1
XFILLER_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _02366_ _04850_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10483__135 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__inv_2
X_08218_ net508 net203 net684 net423 net2368 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a32o_1
X_06479_ top0.CPU.register.registers\[789\] top0.CPU.register.registers\[821\] top0.CPU.register.registers\[853\]
+ top0.CPU.register.registers\[885\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03136_
+ sky130_fd_sc_hd__mux4_1
X_09198_ net603 _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__nor2_1
XFILLER_20_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__10217__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ net211 net616 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10524__176 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__inv_2
XFILLER_121_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ top0.display.delayctr\[17\] _05574_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__nand2_1
XANTENNA__09139__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ top0.CPU.internalMem.pcOut\[31\] _05517_ net652 vssd1 vssd1 vccd1 vccd1 _05529_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__08347__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08121__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold30 top0.CPU.register.registers\[3\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 top0.CPU.register.registers\[98\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 top0.CPU.register.registers\[681\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 top0.CPU.register.registers\[843\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold74 top0.CPU.register.registers\[994\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 top0.CPU.register.registers\[617\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold85 top0.CPU.register.registers\[546\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11993_ net1685 _01632_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06756__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08076__B net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12614_ clknet_leaf_80_clk _02249_ net1113 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10209__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12545_ clknet_leaf_69_clk _02184_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08283__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08822__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ net2168 _02115_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[969\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09619__C net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06605__A _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ clknet_leaf_68_clk _01075_ net1101 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_5 en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10397__49 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08050__A3 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net3279 net119 net113 _05673_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22o_1
XANTENNA__08338__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09535__A0 top0.CPU.control.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06692__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06340__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05850_ top0.CPU.register.registers\[15\] top0.CPU.register.registers\[47\] top0.CPU.register.registers\[79\]
+ top0.CPU.register.registers\[111\] net849 net814 vssd1 vssd1 vccd1 vccd1 _02507_
+ sky130_fd_sc_hd__mux4_1
Xfanout1050 net1055 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1083 net1087 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06444__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1061 net1063 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout1072 net1074 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_2
Xfanout1094 net1106 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_2
XANTENNA__06995__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ _03906_ _04168_ _04169_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__and4_1
X_05781_ top0.CPU.register.registers\[535\] top0.CPU.register.registers\[567\] top0.CPU.register.registers\[599\]
+ top0.CPU.register.registers\[631\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02438_
+ sky130_fd_sc_hd__mux4_1
X_11260__912 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__inv_2
XANTENNA__06058__Y _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07451_ _03282_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06402_ _02983_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__xor2_1
XFILLER_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301__953 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__inv_2
X_07382_ _03919_ _03950_ net459 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__mux2_1
X_10467__119 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__inv_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06333_ net786 _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__and2_1
X_09121_ _04703_ net555 _04832_ net252 net3244 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a32o_1
XANTENNA__08274__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_123_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_135_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06824__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ _04674_ net556 _04810_ net256 net3232 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__a32o_1
X_06264_ top0.CPU.register.registers\[281\] top0.CPU.register.registers\[313\] top0.CPU.register.registers\[345\]
+ top0.CPU.register.registers\[377\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02921_
+ sky130_fd_sc_hd__mux4_1
XFILLER_135_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08003_ top0.CPU.internalMem.pcOut\[1\] net640 net635 _04629_ vssd1 vssd1 vccd1 vccd1
+ _04630_ sky130_fd_sc_hd__o211a_4
XANTENNA__05767__A_N net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06195_ _02850_ _02851_ net580 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_2
Xhold511 top0.CPU.register.registers\[355\] vssd1 vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 top0.CPU.register.registers\[341\] vssd1 vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 top0.CPU.register.registers\[734\] vssd1 vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 top0.CPU.register.registers\[491\] vssd1 vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 top0.CPU.register.registers\[316\] vssd1 vssd1 vccd1 vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08041__A3 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 top0.CPU.register.registers\[642\] vssd1 vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 top0.CPU.register.registers\[600\] vssd1 vssd1 vccd1 vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 top0.CPU.register.registers\[186\] vssd1 vssd1 vccd1 vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 top0.CPU.register.registers\[919\] vssd1 vssd1 vccd1 vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09526__A0 top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1114_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold599 top0.CPU.register.registers\[914\] vssd1 vssd1 vccd1 vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net585 _02910_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__nor2_1
Xhold1200 top0.MMIO.WBData_i\[23\] vssd1 vssd1 vccd1 vccd1 net3422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09885_ _05379_ _05380_ _05383_ _05110_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout574_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05792__C top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ net714 net176 net276 net283 net2717 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__a32o_1
Xhold1211 top0.CPU.intMem_out\[29\] vssd1 vssd1 vccd1 vccd1 net3433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1222 top0.wishbone0.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net3444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07001__B2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08836_ net210 net3157 net353 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__mux2_1
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout741_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05979_ net583 _02634_ _02620_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08767_ _04691_ net317 net290 net2640 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07718_ _03720_ _03972_ _04370_ _03849_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__o221a_1
X_08698_ net224 net3080 net358 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__mux2_1
X_07649_ _04301_ _04303_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ top0.display.delayctr\[20\] top0.display.delayctr\[21\] top0.display.delayctr\[22\]
+ top0.display.delayctr\[23\] vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__or4_1
XFILLER_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11044__696 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_114_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08804__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08280__A3 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ net2022 _01969_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06425__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ net1953 _01900_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_135_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08568__A1 _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ net1884 _01831_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XANTENNA__06674__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
X_10025_ _05487_ _05498_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__nand2_1
XFILLER_49_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06426__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08099__A3 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ net1668 _01615_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_118_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_105_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12528_ net2220 _02167_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1021\]
+ sky130_fd_sc_hd__dfrtp_1
X_12459_ net2151 _02098_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[952\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09756__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08559__A1 _04492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
X_10852__504 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__inv_2
XFILLER_113_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06951_ top0.CPU.register.registers\[536\] top0.CPU.register.registers\[568\] top0.CPU.register.registers\[600\]
+ top0.CPU.register.registers\[632\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03608_
+ sky130_fd_sc_hd__mux4_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ net768 net237 _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__a2bb2o_1
X_05902_ top0.CPU.register.registers\[898\] top0.CPU.register.registers\[930\] top0.CPU.register.registers\[962\]
+ top0.CPU.register.registers\[994\] net831 net796 vssd1 vssd1 vccd1 vccd1 _02559_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08696__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ net720 net167 net322 net331 net2315 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__a32o_1
X_06882_ net864 _03534_ _03537_ _03538_ net747 vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_87_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07534__A2 _03504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06968__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05833_ top0.CPU.register.registers\[18\] top0.CPU.register.registers\[50\] top0.CPU.register.registers\[82\]
+ top0.CPU.register.registers\[114\] net846 net811 vssd1 vssd1 vccd1 vccd1 _02490_
+ sky130_fd_sc_hd__mux4_1
XFILLER_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05764_ _02384_ net632 net626 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__and3_1
X_08552_ net159 net668 net385 net361 net2323 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__a32o_1
X_07503_ _04155_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__nand2_1
XANTENNA__08495__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ net166 net614 net389 net369 net2359 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a32o_1
XANTENNA__07298__A1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05695_ top0.MMIO.WBData_i\[21\] vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout155_A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07434_ _03995_ _03998_ net345 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__mux2_1
XANTENNA__06516__Y _03173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07365_ net339 _04019_ _04021_ net441 _04020_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1064_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_X clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06316_ _02971_ _02972_ net726 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_1
X_09104_ _04695_ net268 net251 net2737 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a22o_1
X_07296_ _03920_ _03952_ net478 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_98_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09035_ top0.CPU.register.registers\[136\] net573 vssd1 vssd1 vccd1 vccd1 _04805_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07470__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06247_ _02902_ _02903_ net731 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__mux2_1
XFILLER_132_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 top0.CPU.register.registers\[375\] vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 top0.CPU.register.registers\[928\] vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ top0.CPU.register.registers\[661\] top0.CPU.register.registers\[693\] top0.CPU.register.registers\[725\]
+ top0.CPU.register.registers\[757\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02835_
+ sky130_fd_sc_hd__mux4_1
Xhold352 net51 vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 top0.CPU.register.registers\[970\] vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 top0.CPU.register.registers\[168\] vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 top0.CPU.intMemAddr\[4\] vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 top0.CPU.register.registers\[376\] vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06656__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout821 net822 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_2
Xfanout810 net819 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_4
X_09937_ _05429_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__nor2_1
Xfanout832 net834 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
X_10595__247 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__inv_2
Xfanout865 net868 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout854 top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09562__Y _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout876 net885 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_2
Xfanout898 net900 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_4
X_09868_ _05355_ _05365_ _05363_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__o21bai_1
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 top0.CPU.register.registers\[120\] vssd1 vssd1 vccd1 vccd1 net3263 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 top0.CPU.register.registers\[183\] vssd1 vssd1 vccd1 vccd1 net3252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06959__S1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout887 net891 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
Xhold1085 top0.CPU.register.registers\[202\] vssd1 vssd1 vccd1 vccd1 net3307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 top0.CPU.register.registers\[147\] vssd1 vssd1 vccd1 vccd1 net3296 sky130_fd_sc_hd__dlygate4sd3_1
X_10636__288 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__inv_2
X_09799_ top0.CPU.internalMem.pcOut\[12\] _05304_ net648 vssd1 vssd1 vccd1 vccd1 _02189_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ net187 net673 net318 net287 net2257 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a32o_1
XFILLER_85_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07804__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1063 top0.CPU.register.registers\[404\] vssd1 vssd1 vccd1 vccd1 net3285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1052 top0.CPU.register.registers\[409\] vssd1 vssd1 vccd1 vccd1 net3274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1096 top0.CPU.register.registers\[365\] vssd1 vssd1 vccd1 vccd1 net3318 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net1522 _01469_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[323\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07015__S net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net1453 _01400_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[254\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__C net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08486__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489__141 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__inv_2
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10293__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ net1384 _01331_ net968 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[185\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08238__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ net2005 _01952_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06895__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05994__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367__19 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__inv_2
X_12244_ net1936 _01883_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[737\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08410__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ net1867 _01814_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[668\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06647__S0 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05870__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ top0.CPU.internalMem.pcOut\[29\] _05496_ vssd1 vssd1 vccd1 vccd1 _05497_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08477__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11959_ net1651 _01598_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_43_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08229__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ net531 net530 net472 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__mux2_1
X_06101_ top0.CPU.control.rs2\[3\] _02753_ _02757_ net774 vssd1 vssd1 vccd1 vccd1
+ _02758_ sky130_fd_sc_hd__o211a_1
X_07081_ _03713_ _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_113_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06886__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06032_ top0.CPU.register.registers\[649\] top0.CPU.register.registers\[681\] top0.CPU.register.registers\[713\]
+ top0.CPU.register.registers\[745\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02689_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09095__B net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06638__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout128 _05101_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout117 net124 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_2
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_2
X_07983_ top0.CPU.intMem_out\[5\] net629 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and2_1
X_09722_ net590 _04604_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a21o_1
XANTENNA__05766__A1 _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05843__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381__33 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__inv_2
X_06934_ net750 _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__nor2_1
X_09653_ net3387 net3379 _05173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
X_06865_ _02618_ _02685_ net542 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout272_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05816_ _02449_ _02452_ _02341_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a21o_1
X_09584_ net666 _05126_ _05127_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__and3_1
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08604_ net2929 net330 _04739_ net717 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06796_ top0.CPU.register.registers\[908\] top0.CPU.register.registers\[940\] top0.CPU.register.registers\[972\]
+ top0.CPU.register.registers\[1004\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03453_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ net3367 net363 _04730_ _02399_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__a22o_1
XANTENNA__07911__X _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05747_ _02393_ _02402_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__and2_2
XANTENNA__08468__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980__632 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__inv_2
XANTENNA_fanout537_A _03092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05678_ top0.MMIO.WBData_i\[31\] vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__inv_2
X_08466_ _04683_ net400 net371 net2637 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout704_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _04662_ net395 net378 net2698 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07348_ _02730_ _03518_ _03738_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__and3_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08174__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_07_1142 vssd1 vssd1 vccd1 vccd1 team_07_1142/HI gpio_out[8] sky130_fd_sc_hd__conb_1
Xteam_07_1153 vssd1 vssd1 vccd1 vccd1 team_07_1153/HI gpio_out[19] sky130_fd_sc_hd__conb_1
XANTENNA__08235__A3 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1197 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] team_07_1197/LO sky130_fd_sc_hd__conb_1
XANTENNA__08640__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1186 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] team_07_1186/LO sky130_fd_sc_hd__conb_1
Xteam_07_1175 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] team_07_1175/LO sky130_fd_sc_hd__conb_1
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ net244 _03934_ _03935_ net448 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__a22o_1
Xteam_07_1164 vssd1 vssd1 vccd1 vccd1 team_07_1164/HI gpio_out[30] sky130_fd_sc_hd__conb_1
XANTENNA__08190__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ net3113 net119 net112 _05590_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a22o_1
XANTENNA__07358__X _04015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ net152 net613 _04802_ net349 net3176 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__a32o_1
XANTENNA__07994__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold171 top0.CPU.register.registers\[813\] vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 top0.CPU.intMemAddr\[21\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06629__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 top0.CPU.register.registers\[165\] vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07746__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 top0.CPU.register.registers\[833\] vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 _02369_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_2
Xfanout640 net641 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06954__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05852__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09292__Y _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout673 net677 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
Xfanout684 net687 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_4
Xfanout662 _04954_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout695 net698 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_4
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08171__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ net1505 _01452_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[306\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08459__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11744_ net1436 _01383_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08474__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ net1367 _01314_ net1009 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07682__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08084__B _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__A3 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100__752 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__inv_2
XANTENNA__06868__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08631__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08304__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06172__X _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ net1919 _01866_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[720\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10135__A _02887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ net1850 _01797_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[651\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12089_ net1781 _01728_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[582\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08698__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__A_N net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07163__B _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08162__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ top0.CPU.register.registers\[514\] top0.CPU.register.registers\[546\] top0.CPU.register.registers\[578\]
+ top0.CPU.register.registers\[610\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__mux4_1
X_10964__616 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__inv_2
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06581_ net762 _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__and2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08320_ net948 _02391_ net545 vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__or3_1
XANTENNA__05899__A top0.CPU.decoder.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__A0 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06476__A2 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ net209 net668 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__and2_1
X_05706__1 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__inv_2
XANTENNA__08870__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ net539 _03053_ net474 vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__mux2_1
X_08182_ net504 net177 net619 net427 net2302 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a32o_1
XANTENNA__06859__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08622__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07133_ net535 _03129_ net473 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout118_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ net530 net532 net472 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__mux2_1
X_10858__510 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06015_ top0.CPU.register.registers\[902\] top0.CPU.register.registers\[934\] top0.CPU.register.registers\[966\]
+ top0.CPU.register.registers\[998\] net844 net809 vssd1 vssd1 vccd1 vccd1 _02672_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07728__A2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06087__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10193__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ net720 net511 net181 net547 net2313 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a32o_1
X_09705_ top0.CPU.internalMem.pcOut\[5\] _05217_ net650 vssd1 vssd1 vccd1 vccd1 _02182_
+ sky130_fd_sc_hd__mux2_1
X_06917_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__inv_2
XANTENNA__08689__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ _04476_ _04541_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a21o_1
X_09636_ _02748_ _05150_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_94_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06164__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ _03490_ net526 vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07361__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07900__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout821_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ net589 _04632_ _05111_ _02351_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06779_ top0.CPU.register.registers\[14\] top0.CPU.register.registers\[46\] top0.CPU.register.registers\[78\]
+ top0.CPU.register.registers\[110\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03436_
+ sky130_fd_sc_hd__mux4_1
X_09498_ top0.MMIO.WBData_i\[6\] net139 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout919_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net158 net679 net386 net365 net2687 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__a32o_1
XANTENNA__06011__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08449_ net2864 net215 net373 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06417__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ clknet_leaf_66_clk _01108_ net1104 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09405__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08613__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ clknet_leaf_59_clk _01039_ net1091 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10342_ net2253 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08124__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05978__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10273_ net2978 net121 net113 _05658_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a22o_1
X_12012_ net1704 _01651_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[505\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06078__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10651__303 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__inv_2
XFILLER_93_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout481 _02575_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_2
XFILLER_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_2
Xfanout492 net496 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xclkbuf_leaf_85_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ net767 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07104__A0 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09644__A2 _05169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ net1419 _01366_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ net1350 _01297_ net965 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[151\]
+ sky130_fd_sc_hd__dfrtp_1
X_11589_ net1281 _01228_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07407__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold907 top0.CPU.register.registers\[275\] vssd1 vssd1 vccd1 vccd1 net3129 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold918 top0.CPU.register.registers\[881\] vssd1 vssd1 vccd1 vccd1 net3140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 top0.CPU.register.registers\[506\] vssd1 vssd1 vccd1 vccd1 net3151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06069__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07820_ _02339_ _02385_ _02387_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__or3_1
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08383__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _03720_ _04057_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__nor2_1
XANTENNA__07174__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ _03340_ _03357_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__and3_1
XANTENNA__08686__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ net442 _04152_ _04266_ _03760_ _04335_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_121_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09421_ top0.CPU.Op\[5\] _02409_ net626 _05000_ _05005_ vssd1 vssd1 vccd1 vccd1 _05025_
+ sky130_fd_sc_hd__o41ai_1
XFILLER_65_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06633_ top0.CPU.register.registers\[515\] top0.CPU.register.registers\[547\] top0.CPU.register.registers\[579\]
+ top0.CPU.register.registers\[611\] net913 net879 vssd1 vssd1 vccd1 vccd1 _03290_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09096__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ _04995_ _04997_ _04998_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.state_n\[2\]
+ sky130_fd_sc_hd__or3_1
XANTENNA__06077__X _02734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06564_ net858 _03216_ _03220_ _03208_ _03212_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__o32a_4
X_08303_ net2854 _04566_ net415 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__mux2_1
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08843__A0 _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07646__A1 _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ top0.wishbone0.curr_state\[1\] top0.wishbone0.curr_state\[2\] net1 vssd1
+ vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout235_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06495_ _03134_ net447 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__or2_1
XANTENNA__07646__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ net497 net215 net680 net421 net2364 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a32o_1
XANTENNA__06952__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout402_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08165_ net223 net620 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07116_ net477 _03754_ _03771_ _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_132_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08096_ net509 net184 net696 net434 net2377 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a32o_1
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08071__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload80 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07047_ net519 _03701_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__xor2_2
XANTENNA__07068__B _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09020__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout869_A top0.CPU.decoder.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net168 net696 net277 net260 net2415 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__a32o_1
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07084__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ net637 _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_67_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07885__A1 top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09619_ _02715_ _04952_ net660 _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__nor4_1
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ clknet_leaf_80_clk _02265_ net1113 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07023__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05991__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08119__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09087__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ clknet_leaf_54_clk _02200_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08834__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ net1204 _01151_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09298__X _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12492_ net2184 _02131_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[985\]
+ sky130_fd_sc_hd__dfrtp_1
X_11443_ clknet_leaf_78_clk _01091_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.Op\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11374_ clknet_leaf_74_clk top0.CPU.internalMem.load2Ct_n\[0\] net1123 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.load2Ct\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06163__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06073__B1 _02729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171__823 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__inv_2
XANTENNA__05820__A0 _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ net2225 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10256_ _04938_ _05134_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__or2_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11212__864 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ net129 _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__nor2_1
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_74_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09078__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06280_ top0.CPU.register.registers\[282\] top0.CPU.register.registers\[314\] top0.CPU.register.registers\[346\]
+ top0.CPU.register.registers\[378\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02937_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07169__A _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold737 top0.CPU.register.registers\[775\] vssd1 vssd1 vccd1 vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 top0.CPU.register.registers\[519\] vssd1 vssd1 vccd1 vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 top0.CPU.register.registers\[262\] vssd1 vssd1 vccd1 vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
X_10820__472 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__inv_2
XANTENNA__11721__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold726 top0.CPU.register.registers\[497\] vssd1 vssd1 vccd1 vccd1 net2948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 top0.CPU.register.registers\[415\] vssd1 vssd1 vccd1 vccd1 net2981 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ top0.CPU.internalMem.pcOut\[26\] _05459_ vssd1 vssd1 vccd1 vccd1 _05462_
+ sky130_fd_sc_hd__xnor2_1
Xhold748 top0.CPU.register.registers\[669\] vssd1 vssd1 vccd1 vccd1 net2970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08699__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__X _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ top0.CPU.register.registers\[219\] net567 vssd1 vssd1 vccd1 vccd1 _04774_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09002__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ net187 net3280 net355 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__mux2_1
XANTENNA__06520__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _03482_ net526 _03519_ net524 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout185_A _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
X_08783_ net195 net687 net319 net291 net2367 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a32o_1
XANTENNA__06462__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05995_ top0.CPU.register.registers\[647\] top0.CPU.register.registers\[679\] top0.CPU.register.registers\[711\]
+ top0.CPU.register.registers\[743\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02652_
+ sky130_fd_sc_hd__mux4_1
X_07734_ net451 _04028_ _04033_ _03846_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__a22o_1
X_07665_ _03445_ _04320_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07632__A _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06616_ net864 _03268_ _03271_ _03272_ net860 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout352_A _04798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ net2860 _04949_ _05015_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1094_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_36_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A2 _05006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07596_ net245 _03957_ _04169_ net441 _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__o221a_1
XANTENNA__05973__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ _04975_ _04983_ _02517_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a21o_1
XFILLER_80_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06547_ net540 _03200_ _02812_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _04918_ _04926_ _04927_ _04898_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a211o_1
XANTENNA__09084__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__A1 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ top0.CPU.register.registers\[917\] top0.CPU.register.registers\[949\] top0.CPU.register.registers\[981\]
+ top0.CPU.register.registers\[1013\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03135_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_134_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155__807 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__inv_2
X_08217_ net2962 net424 _04701_ net516 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ top0.display.state\[2\] _04857_ _02359_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__o21ai_1
X_08148_ net2887 net426 _04674_ net503 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a22o_1
XANTENNA__08044__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08595__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08079_ net3118 net436 _04662_ net500 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a22o_1
X_10110_ top0.display.delayctr\[17\] _05574_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__or2_1
XANTENNA__07807__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10041_ top0.CPU.internalMem.pcOut\[31\] _05517_ vssd1 vssd1 vccd1 vccd1 _05528_
+ sky130_fd_sc_hd__or2_1
XFILLER_88_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold31 top0.CPU.register.registers\[8\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xhold20 top0.CPU.register.registers\[0\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 top0.CPU.register.registers\[434\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top0.CPU.register.registers\[626\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 top0.CPU.register.registers\[427\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
X_11049__701 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__inv_2
Xhold86 top0.CPU.register.registers\[51\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ net1684 _01631_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[485\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold97 top0.CPU.register.registers\[882\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 top0.CPU.register.registers\[739\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05869__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05964__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ clknet_leaf_80_clk _02248_ net1112 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
X_10763__415 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__inv_2
XANTENNA__08807__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ clknet_leaf_78_clk _02183_ net1115 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08283__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08822__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ net2167 _02114_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[968\]
+ sky130_fd_sc_hd__dfrtp_1
X_10804__456 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__inv_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ clknet_leaf_60_clk _01074_ net1094 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08035__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10308_ _03700_ net551 net144 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06141__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06692__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ net11 net656 net595 top0.MMIO.WBData_i\[18\] vssd1 vssd1 vccd1 vccd1 _02285_
+ sky130_fd_sc_hd__a22o_1
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
XFILLER_79_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1051 net1054 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1062 net1063 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1095 net1097 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout1084 net1087 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05780_ top0.CPU.register.registers\[663\] top0.CPU.register.registers\[695\] top0.CPU.register.registers\[727\]
+ top0.CPU.register.registers\[759\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02437_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08510__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08267__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07171__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07450_ _03364_ _03381_ _03380_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a21o_1
XFILLER_50_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11340__992 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__inv_2
X_06401_ _02927_ _02944_ _02962_ net544 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a31o_1
X_07381_ _03951_ _03980_ net458 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__mux2_1
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06332_ top0.CPU.register.registers\[925\] top0.CPU.register.registers\[957\] top0.CPU.register.registers\[989\]
+ top0.CPU.register.registers\[1021\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__mux4_1
X_09120_ top0.CPU.register.registers\[78\] net569 vssd1 vssd1 vccd1 vccd1 _04832_
+ sky130_fd_sc_hd__or2_1
X_09051_ top0.CPU.register.registers\[125\] net569 vssd1 vssd1 vccd1 vccd1 _04810_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_116_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10547__199 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__inv_2
X_08002_ top0.CPU.intMem_out\[1\] net630 _04588_ _04628_ vssd1 vssd1 vccd1 vccd1 _04629_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06263_ top0.CPU.register.registers\[409\] top0.CPU.register.registers\[441\] top0.CPU.register.registers\[473\]
+ top0.CPU.register.registers\[505\] net825 net790 vssd1 vssd1 vccd1 vccd1 _02920_
+ sky130_fd_sc_hd__mux4_1
X_06194_ net822 net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a21oi_2
Xhold501 top0.CPU.register.registers\[795\] vssd1 vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 top0.CPU.register.registers\[627\] vssd1 vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 net41 vssd1 vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_1
Xhold534 top0.CPU.register.registers\[826\] vssd1 vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 top0.CPU.register.registers\[174\] vssd1 vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05846__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold578 net43 vssd1 vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 top0.CPU.register.registers\[911\] vssd1 vssd1 vccd1 vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 top0.CPU.register.registers\[733\] vssd1 vssd1 vccd1 vccd1 net2789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 top0.CPU.register.registers\[975\] vssd1 vssd1 vccd1 vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ top0.CPU.internalMem.pcOut\[24\] net645 _05443_ _05446_ vssd1 vssd1 vccd1
+ vccd1 _02201_ sky130_fd_sc_hd__o22a_1
XANTENNA__08329__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1107_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _05381_ _05382_ net647 vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__o21a_1
X_08904_ net718 net218 net277 net283 net2438 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__a32o_1
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07346__B _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1223 top0.MMIO.WBData_i\[11\] vssd1 vssd1 vccd1 vccd1 net3445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 top0.CPU.intMem_out\[3\] vssd1 vssd1 vccd1 vccd1 net3434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_4_0_clk_X clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 top0.display.delayctr\[17\] vssd1 vssd1 vccd1 vccd1 net3423 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07001__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08835_ _04498_ net3154 net354 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__mux2_1
X_08766_ _04690_ net324 net292 net2605 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a22o_1
XANTENNA__08729__Y _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout567_A _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05978_ net583 _02634_ _02620_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a21boi_4
X_07717_ net485 _03945_ _04373_ net244 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout734_A _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ net212 net3041 net359 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
XANTENNA__06199__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450__102 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__inv_2
XANTENNA__06249__Y _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08501__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07648_ net245 _03911_ _04304_ net449 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05946__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout901_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ net449 _03379_ net444 _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__o31a_1
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09289__A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ top0.display.delayctr\[24\] top0.display.delayctr\[25\] top0.display.delayctr\[26\]
+ top0.display.delayctr\[27\] vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__or4_2
XFILLER_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08265__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06371__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ net769 top0.CPU.intMemAddr\[7\] net610 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__o21a_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12260_ net1952 _01899_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[753\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08017__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ net1883 _01830_ net1101 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[684\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__08132__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06674__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__X _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__nand2_1
XANTENNA__06426__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11283__935 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__inv_2
X_11975_ net1667 _01614_ net1000 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08087__B net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324__976 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__inv_2
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08307__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07563__A1_N _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06362__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__C net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12527_ net2219 _02166_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1020\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08831__A top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net2150 _02097_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[951\]
+ sky130_fd_sc_hd__dfrtp_1
X_11409_ clknet_leaf_87_clk _01057_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11218__870 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__inv_2
XANTENNA__06622__Y _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12389_ net2081 _02028_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06351__A top0.CPU.control.funct7\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891__543 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__inv_2
XFILLER_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07519__B1 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ top0.CPU.register.registers\[664\] top0.CPU.register.registers\[696\] top0.CPU.register.registers\[728\]
+ top0.CPU.register.registers\[760\] net923 net889 vssd1 vssd1 vccd1 vccd1 _03607_
+ sky130_fd_sc_hd__mux4_1
X_06881_ net871 _03535_ net751 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21o_1
X_05901_ _02556_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08731__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05832_ top0.CPU.register.registers\[146\] top0.CPU.register.registers\[178\] top0.CPU.register.registers\[210\]
+ top0.CPU.register.registers\[242\] net846 net811 vssd1 vssd1 vccd1 vccd1 _02489_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10932__584 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__inv_2
X_08620_ net715 net171 net312 net330 net2502 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__a32o_1
X_05763_ top0.CPU.Op\[4\] _02371_ _02373_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__or3_1
X_08551_ net161 net668 net391 net361 net2307 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__a32o_1
X_05694_ top0.MMIO.WBData_i\[30\] vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__inv_2
X_07502_ _04156_ _04157_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__or2_1
X_08482_ net214 net616 net390 net369 net2551 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a32o_1
X_07433_ _04070_ _04071_ net344 vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_46_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout148_A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07364_ _02698_ _03540_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__xor2_1
X_09103_ _04694_ net552 _04826_ net251 net3262 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__a32o_1
XANTENNA__06353__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06315_ top0.CPU.register.registers\[28\] top0.CPU.register.registers\[60\] top0.CPU.register.registers\[92\]
+ top0.CPU.register.registers\[124\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02972_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ _03950_ _03951_ net459 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__mux2_1
X_09034_ net180 net613 _04804_ net351 net3325 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_98_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06246_ top0.CPU.register.registers\[280\] top0.CPU.register.registers\[312\] top0.CPU.register.registers\[344\]
+ top0.CPU.register.registers\[376\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02903_
+ sky130_fd_sc_hd__mux4_1
Xhold320 top0.CPU.register.registers\[717\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09747__B2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06105__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold331 top0.CPU.register.registers\[702\] vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 top0.CPU.intMemAddr\[27\] vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ net246 _02771_ _02791_ _02832_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand4_2
Xhold353 top0.CPU.register.registers\[451\] vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold375 top0.CPU.register.registers\[322\] vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
Xhold386 top0.CPU.register.registers\[695\] vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 top0.CPU.register.registers\[835\] vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06656__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold397 top0.CPU.register.registers\[559\] vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout822 top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__buf_2
XFILLER_104_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout811 net819 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_2
X_09936_ _05387_ _05402_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_2
X_11267__919 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__inv_2
Xfanout855 net857 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_129_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout844 net854 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
Xfanout866 net868 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
XANTENNA_fanout851_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout899 net900 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout949_A top0.CPU.decoder.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _05365_ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__or2_1
Xhold1042 top0.CPU.register.registers\[240\] vssd1 vssd1 vccd1 vccd1 net3264 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 top0.CPU.register.registers\[263\] vssd1 vssd1 vccd1 vccd1 net3242 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 net879 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
Xfanout888 net891 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_4
Xhold1031 top0.CPU.register.registers\[281\] vssd1 vssd1 vccd1 vccd1 net3253 sky130_fd_sc_hd__dlygate4sd3_1
X_11011__663 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__inv_2
X_08818_ net191 net677 net327 net288 net2317 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__a32o_1
X_09798_ net240 _05300_ _05301_ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__o31ai_1
Xhold1075 top0.CPU.register.registers\[72\] vssd1 vssd1 vccd1 vccd1 net3297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07804__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1064 top0.CPU.register.registers\[407\] vssd1 vssd1 vccd1 vccd1 net3286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 top0.CPU.register.registers\[64\] vssd1 vssd1 vccd1 vccd1 net3275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1097 top0.CPU.register.registers\[403\] vssd1 vssd1 vccd1 vccd1 net3319 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ top0.CPU.register.registers\[365\] net572 _04736_ vssd1 vssd1 vccd1 vccd1
+ _04748_ sky130_fd_sc_hd__o21a_1
XANTENNA__06200__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1086 top0.CPU.register.registers\[148\] vssd1 vssd1 vccd1 vccd1 net3308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11760_ net1452 _01399_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ net1383 _01330_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[184\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08127__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08238__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08789__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net2004 _01951_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06870__S net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__X _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06895__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09738__A1 top0.CPU.control.funct7\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ net1935 _01882_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[736\]
+ sky130_fd_sc_hd__dfrtp_1
X_10875__527 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08410__A1 _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06647__S1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ net1866 _01813_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08961__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10916__568 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__inv_2
X_10007_ _03003_ _04489_ net589 vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__mux2_1
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07714__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769__421 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11958_ net1650 _01597_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[451\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11889_ net1581 _01528_ net1050 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08229__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07437__C1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06100_ net740 _02756_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__or2_1
XANTENNA__07988__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07080_ _02428_ _02430_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__nand2_1
XANTENNA__06780__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06031_ top0.CPU.register.registers\[777\] top0.CPU.register.registers\[809\] top0.CPU.register.registers\[841\]
+ top0.CPU.register.registers\[873\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02688_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06886__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06638__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08952__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout129 _05638_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
X_07982_ net562 _04612_ _04588_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_93_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout118 net124 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09392__A _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ top0.CPU.control.funct7\[2\] net631 _02453_ vssd1 vssd1 vccd1 vccd1 _05232_
+ sky130_fd_sc_hd__and3_1
X_06933_ _03588_ _03589_ net869 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__mux2_1
X_09652_ top0.MISOtoMMIO\[2\] net3387 _05173_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
X_06864_ _03507_ _03518_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__xnor2_2
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08180__A3 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06795_ top0.CPU.register.registers\[780\] top0.CPU.register.registers\[812\] top0.CPU.register.registers\[844\]
+ top0.CPU.register.registers\[876\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03452_
+ sky130_fd_sc_hd__mux4_1
XFILLER_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09583_ _05121_ _05125_ top0.display.counter\[2\] vssd1 vssd1 vccd1 vccd1 _05127_
+ sky130_fd_sc_hd__or3b_1
X_05815_ _02449_ _02452_ _02341_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__a21oi_4
X_08603_ net205 net314 vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05746_ _02393_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__nand2_1
X_08534_ _02404_ net202 net673 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__and3_1
XFILLER_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08465_ _04682_ net396 net370 net3078 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
X_07416_ _03263_ _03385_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nor2_1
XANTENNA__07691__A2 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ _04661_ net385 net377 net2608 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07347_ _04002_ _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__and2_1
Xteam_07_1154 vssd1 vssd1 vccd1 vccd1 team_07_1154/HI gpio_out[20] sky130_fd_sc_hd__conb_1
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10562__214 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__inv_2
Xteam_07_1143 vssd1 vssd1 vccd1 vccd1 team_07_1143/HI gpio_out[9] sky130_fd_sc_hd__conb_1
XANTENNA_fanout899_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1165 vssd1 vssd1 vccd1 vccd1 team_07_1165/HI gpio_out[31] sky130_fd_sc_hd__conb_1
Xteam_07_1187 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] team_07_1187/LO sky130_fd_sc_hd__conb_1
X_07278_ _03735_ _03768_ net488 vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__mux2_1
Xteam_07_1176 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] team_07_1176/LO sky130_fd_sc_hd__conb_1
X_09017_ top0.CPU.register.registers\[151\] net567 vssd1 vssd1 vccd1 vccd1 _04802_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08190__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__B _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06229_ _02882_ _02885_ net780 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__mux2_1
XANTENNA__07994__A3 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 top0.CPU.register.registers\[488\] vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06629__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 top0.CPU.register.registers\[224\] vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
X_10603__255 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__inv_2
XANTENNA__07087__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 top0.CPU.register.registers\[495\] vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold172 top0.CPU.register.registers\[847\] vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08943__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 top0.CPU.register.registers\[706\] vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout641 _02383_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_2
Xfanout630 _02419_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06954__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net676 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_4
Xfanout652 _02368_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_8
X_09919_ _05411_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__xnor2_1
Xfanout663 net664 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_2
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07026__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_29_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05914__C1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11812_ net1504 _01451_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[305\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11743_ net1435 _01382_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[236\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ net1366 _01313_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08084__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427__79 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__inv_2
XANTENNA__06317__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12226_ net1918 _01865_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[719\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_12_0_clk_X clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ net1849 _01796_ net1029 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[650\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08934__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11289__941 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__inv_2
XANTENNA__08395__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05944__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12088_ net1780 _01727_ net1029 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06580_ top0.CPU.register.registers\[272\] top0.CPU.register.registers\[304\] top0.CPU.register.registers\[336\]
+ top0.CPU.register.registers\[368\] net931 net897 vssd1 vssd1 vccd1 vccd1 _03237_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05920__A2 _02553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06556__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08250_ net2865 net417 _04710_ net494 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a22o_1
XANTENNA__06881__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08181_ net506 net220 net619 net427 net2584 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a32o_1
X_07201_ _03005_ _03053_ net341 _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a22o_1
XFILLER_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07132_ net457 _03787_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__or2_1
XANTENNA__06363__X _03020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08622__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07063_ net449 _03719_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__or2_4
X_06014_ top0.CPU.register.registers\[774\] top0.CPU.register.registers\[806\] top0.CPU.register.registers\[838\]
+ top0.CPU.register.registers\[870\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02671_
+ sky130_fd_sc_hd__mux4_1
X_10441__93 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__inv_2
X_10938__590 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__inv_2
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07728__A3 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08386__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ top0.CPU.internalMem.pcOut\[9\] net641 net636 _04599_ vssd1 vssd1 vccd1 vccd1
+ _04600_ sky130_fd_sc_hd__o211a_2
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout382_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ net241 _05215_ _05216_ _05213_ _05214_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06916_ _03225_ net533 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09272__D _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07896_ top0.CPU.intMem_out\[20\] net627 _02854_ net591 net642 vssd1 vssd1 vccd1
+ vccd1 _04542_ sky130_fd_sc_hd__a221o_1
X_09635_ net3334 net605 net659 net3328 _05163_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06847_ net747 _03503_ _03498_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__a21oi_4
X_11082__734 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__inv_2
X_09566_ _02351_ _05113_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__xnor2_1
X_06778_ top0.CPU.register.registers\[142\] top0.CPU.register.registers\[174\] top0.CPU.register.registers\[206\]
+ top0.CPU.register.registers\[238\] net921 net887 vssd1 vssd1 vccd1 vccd1 _03435_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout814_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ top0.MMIO.WBData_i\[11\] net137 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05729_ top0.CPU.Op\[5\] _02379_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__nand2_4
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08517_ net161 net679 net386 net365 net2327 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a32o_1
X_08448_ net2977 net170 net375 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__mux2_1
X_11123__775 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__inv_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08379_ net175 net702 net390 net382 net2820 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a32o_1
XFILLER_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08613__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ clknet_leaf_59_clk _01038_ net1091 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10341_ net2237 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09169__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10272_ net144 _05158_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__nand2_1
XANTENNA__05978__A2 _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_12011_ net1703 _01650_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[504\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_105_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08140__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690__342 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__inv_2
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_2
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_2
Xfanout482 net484 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_2
Xfanout493 net496 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_2
XANTENNA__08144__A3 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987__639 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__inv_2
XFILLER_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731__383 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__inv_2
XANTENNA__10239__B2 top0.MMIO.WBData_i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ net767 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07104__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11726_ net1418 _01365_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[219\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ net1349 _01296_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[150\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08315__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08604__B2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11588_ net1280 _01227_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07407__A2 _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06615__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold919 top0.CPU.register.registers\[987\] vssd1 vssd1 vccd1 vccd1 net3141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold908 top0.CPU.register.registers\[765\] vssd1 vssd1 vccd1 vccd1 net3130 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06091__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06710__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08368__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ net1901 _01848_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07591__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ net451 _03758_ _04053_ _04404_ _04406_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__a311o_1
XFILLER_38_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07174__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066__718 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__inv_2
X_06701_ _03321_ _03322_ _03338_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__nand3_1
XANTENNA__08540__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ net454 _04268_ _04337_ _03719_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__a211o_1
XANTENNA__06777__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09420_ _05004_ _05008_ _05023_ _04948_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__o31ai_1
XFILLER_92_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07894__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06632_ top0.CPU.register.registers\[643\] top0.CPU.register.registers\[675\] top0.CPU.register.registers\[707\]
+ top0.CPU.register.registers\[739\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03289_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05703__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _04850_ _04863_ _04865_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__o21ba_1
X_06563_ net866 _03219_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__nor2_1
X_11107__759 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__inv_2
X_09282_ _04934_ _04938_ _04940_ top0.wishbone0.curr_state\[0\] vssd1 vssd1 vccd1
+ vccd1 _04942_ sky130_fd_sc_hd__o211ai_2
XANTENNA__06529__S0 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06518__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08302_ net3224 _04561_ net413 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
X_08233_ net509 net169 net685 net424 net2408 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a32o_1
X_06494_ _03134_ net447 vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__and2_1
XANTENNA__06303__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08164_ net3110 net426 _04682_ net501 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a22o_1
X_08095_ net504 net188 net694 net434 net2476 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a32o_1
X_07115_ net474 net457 net539 vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__or3_1
Xclkload70 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_16
X_07046_ net519 _03701_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__nor2_1
XANTENNA__08071__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload81 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_8
XANTENNA__08359__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload92 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__inv_16
X_10674__326 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__inv_2
XANTENNA__10166__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08997_ net171 net691 _04796_ net259 net3301 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ top0.CPU.internalMem.pcOut\[12\] net643 _04584_ _04585_ vssd1 vssd1 vccd1
+ vccd1 _04586_ sky130_fd_sc_hd__a22o_1
X_10715__367 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__inv_2
XFILLER_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout931_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ top0.CPU.internalMem.pcOut\[23\] net638 net633 _04527_ vssd1 vssd1 vccd1
+ vccd1 _04528_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ net577 _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__or2_1
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08196__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ top0.CPU.control.funct7\[2\] _05062_ net126 vssd1 vssd1 vccd1 vccd1 _01118_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05896__A1 top0.CPU.decoder.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05896__B2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09087__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05991__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10568__220 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__inv_2
X_12560_ clknet_leaf_54_clk _02199_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_11511_ net1203 _01150_ net970 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12491_ net2183 _02130_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[984\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08135__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11442_ clknet_leaf_60_clk _01090_ net1100 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10609__261 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__inv_2
XANTENNA__06940__S0 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06073__A1 top0.CPU.control.funct7\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ net2235 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ net3101 net117 net111 _05650_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
X_10186_ _04943_ _04942_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_72_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08770__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 _04749_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06759__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08522__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload6_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05887__A1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_17_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ net1401 _01348_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[202\]
+ sky130_fd_sc_hd__dfrtp_1
X_12689_ clknet_leaf_92_clk _02324_ net1082 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06931__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 top0.CPU.register.registers\[511\] vssd1 vssd1 vccd1 vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349__1001 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__inv_2
XFILLER_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold727 top0.CPU.register.registers\[59\] vssd1 vssd1 vccd1 vccd1 net2949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold705 top0.CPU.register.registers\[727\] vssd1 vssd1 vccd1 vccd1 net2927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07261__A0 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold738 top0.CPU.register.registers\[247\] vssd1 vssd1 vccd1 vccd1 net2960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 top0.CPU.register.registers\[888\] vssd1 vssd1 vccd1 vccd1 net2971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07737__X _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10411__63 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__inv_2
X_08920_ _04640_ net553 _04773_ net263 net3082 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__a32o_1
X_08851_ net191 net3125 net356 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__mux2_1
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07802_ net534 _03221_ net533 net525 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__and4_1
XANTENNA__07564__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05994_ net454 _02650_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__nor2_1
X_08782_ _04703_ net316 net290 net2718 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__a22o_1
XANTENNA__08287__Y _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ _03601_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07664_ _03563_ _04298_ _03445_ _03484_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08513__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_A _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06615_ net761 _03269_ net751 vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__a21o_1
X_09403_ top0.MMIO.WBData_i\[0\] net147 net143 top0.MISOtoMMIO\[0\] _05014_ vssd1
+ vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__o221a_1
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_36_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ net487 net531 net444 _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__o31a_1
XFILLER_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05973__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _04589_ _04976_ _04978_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__o31ai_1
X_06546_ net540 _03200_ _02812_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07619__A2 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1195_A top0.CPU.intMem_out\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _04922_ _04924_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__or2_1
X_06477_ _02852_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__xor2_1
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_clk_X clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08216_ _04549_ _04688_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nor2_1
X_11194__846 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__inv_2
X_09196_ top0.display.state\[2\] _04857_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__nand2_1
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ net224 net618 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__and2_1
XANTENNA__08044__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ net205 net693 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__and2_1
X_11235__887 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__inv_2
X_07029_ _02380_ _02447_ _02449_ _02452_ _02341_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout979_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__B1 _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__B _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__B1_N _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _05520_ _05523_ _05524_ _05526_ net238 vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__a311o_1
XFILLER_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08347__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 top0.CPU.register.registers\[15\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold21 top0.CPU.register.registers\[27\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold10 top0.CPU.register.registers\[14\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06989__S0 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 top0.CPU.register.registers\[811\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold43 top0.CPU.register.registers\[550\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
X_11088__740 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__inv_2
Xhold54 top0.CPU.register.registers\[160\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 top0.CPU.register.registers\[553\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 top0.CPU.register.registers\[552\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net1683 _01630_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[484\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold98 top0.CPU.register.registers\[609\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08504__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11129__781 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__inv_2
XANTENNA__05869__A1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05964__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06873__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12612_ clknet_leaf_80_clk _02247_ net1112 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08807__A1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12543_ clknet_leaf_78_clk _02182_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10843__495 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__inv_2
X_12474_ net2166 _02113_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[967\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ clknet_leaf_60_clk _01073_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08035__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06902__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ net3250 net119 net114 _05672_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a22o_1
XANTENNA__07794__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06141__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ net10 net656 net595 top0.MMIO.WBData_i\[17\] vssd1 vssd1 vccd1 vccd1 _02284_
+ sky130_fd_sc_hd__a22o_1
Xfanout1030 net1056 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08743__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1052 net1054 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
Xfanout1041 net1055 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_2
X_10169_ _04970_ _05604_ top0.display.delayctr\[28\] vssd1 vssd1 vccd1 vccd1 _05627_
+ sky130_fd_sc_hd__o21ai_1
Xfanout1063 net1065 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_4
Xfanout1074 net1088 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_2
XFILLER_66_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08510__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06400_ _03041_ _03053_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__nand2_1
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07380_ _04035_ _04036_ net345 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__mux2_1
X_06331_ top0.CPU.register.registers\[797\] top0.CPU.register.registers\[829\] top0.CPU.register.registers\[861\]
+ top0.CPU.register.registers\[893\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02988_
+ sky130_fd_sc_hd__mux4_1
X_09050_ _04673_ net279 net258 net2771 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__a22o_1
XANTENNA__06285__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06262_ net776 _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ net563 _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_116_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 top0.CPU.register.registers\[342\] vssd1 vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
X_06193_ net771 _02841_ _02845_ _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__o2bb2a_2
Xhold524 top0.CPU.register.registers\[779\] vssd1 vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 net79 vssd1 vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09395__A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold513 top0.CPU.register.registers\[443\] vssd1 vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 top0.CPU.register.registers\[649\] vssd1 vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08982__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ net238 _05444_ _05445_ net652 vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a31o_1
XANTENNA__06588__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 top0.CPU.register.registers\[564\] vssd1 vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 top0.CPU.register.registers\[725\] vssd1 vssd1 vccd1 vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 top0.CPU.register.registers\[515\] vssd1 vssd1 vccd1 vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ net720 net180 _04769_ net283 net3333 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__a32o_1
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09883_ top0.CPU.internalMem.pcOut\[18\] _05359_ top0.CPU.internalMem.pcOut\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout295_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__B2 _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05891__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 top0.MMIO.WBData_i\[15\] vssd1 vssd1 vccd1 vccd1 net3446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1213 net69 vssd1 vssd1 vccd1 vccd1 net3435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1202 top0.display.delayctr\[16\] vssd1 vssd1 vccd1 vccd1 net3424 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net224 net3299 net354 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1002_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ net688 _04738_ net292 net2604 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__a22o_1
XFILLER_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07362__B net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05977_ net772 _02633_ _02628_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__o21ai_4
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07716_ _03764_ net338 _03780_ _02577_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__a22o_1
X_08696_ _04481_ net2981 net360 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
XANTENNA__07930__X _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06199__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786__438 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__inv_2
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08501__A3 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_A _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07647_ net517 _03838_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ net443 _04166_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__a21oi_1
X_10530__182 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05946__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06529_ top0.CPU.register.registers\[274\] top0.CPU.register.registers\[306\] top0.CPU.register.registers\[338\]
+ top0.CPU.register.registers\[370\] net931 net897 vssd1 vssd1 vccd1 vccd1 _03186_
+ sky130_fd_sc_hd__mux4_1
X_09317_ _04967_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__or2_1
X_10827__479 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__inv_2
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08265__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06371__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _04088_ net233 net227 _02337_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a31o_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ net213 net669 net270 net247 net2310 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__a32o_1
XANTENNA__08017__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_12190_ net1882 _01829_ net1007 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[683\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08921__B net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_102_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10023_ top0.CPU.internalMem.pcOut\[30\] _05509_ vssd1 vssd1 vccd1 vccd1 _05511_
+ sky130_fd_sc_hd__or2_1
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07272__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ net1666 _01613_ net1122 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09150__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348__1000 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08256__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12526_ net2218 _02165_ net991 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1019\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06362__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ net2149 _02096_ net1074 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[950\]
+ sky130_fd_sc_hd__dfrtp_1
X_11408_ clknet_leaf_87_clk _01056_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05947__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12388_ net2080 _02027_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05873__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06880_ net761 _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__and2_1
X_05900_ _02376_ _02447_ _02450_ net734 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a31o_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05831_ _02486_ _02487_ net785 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10473__125 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__inv_2
XFILLER_67_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05762_ _02371_ _02372_ _02339_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__and3b_1
X_08550_ net166 net668 net389 net361 net2266 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a32o_1
X_08481_ net169 net621 net402 net372 net2434 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a32o_1
X_05693_ top0.CPU.internalMem.pcOut\[0\] vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__inv_2
X_07501_ _02790_ _03443_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nand2_1
X_10514__166 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__inv_2
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07432_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09444__A1 top0.MMIO.WBData_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ _02699_ net525 net444 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__or3_1
X_09102_ top0.CPU.register.registers\[90\] net564 vssd1 vssd1 vccd1 vccd1 _04826_
+ sky130_fd_sc_hd__or2_1
X_06314_ top0.CPU.register.registers\[156\] top0.CPU.register.registers\[188\] top0.CPU.register.registers\[220\]
+ top0.CPU.register.registers\[252\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02971_
+ sky130_fd_sc_hd__mux4_1
X_07294_ _03129_ net535 net467 vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__mux2_1
XANTENNA__06353__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09033_ top0.CPU.register.registers\[137\] net573 vssd1 vssd1 vccd1 vccd1 _04804_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout210_A _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06245_ top0.CPU.register.registers\[408\] top0.CPU.register.registers\[440\] top0.CPU.register.registers\[472\]
+ top0.CPU.register.registers\[504\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02902_
+ sky130_fd_sc_hd__mux4_1
Xhold310 top0.CPU.register.registers\[690\] vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07638__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06176_ net246 _02771_ _02791_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout308_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold332 top0.CPU.register.registers\[303\] vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06105__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 top0.CPU.register.registers\[1010\] vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 top0.CPU.register.registers\[353\] vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 top0.CPU.register.registers\[703\] vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 top0.CPU.register.registers\[810\] vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 top0.CPU.register.registers\[592\] vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 top0.CPU.register.registers\[866\] vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout812 net814 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_4
X_09935_ _05411_ _05422_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__nand2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout834 top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_2
Xfanout823 net825 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
Xfanout801 net805 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_4
Xhold398 top0.CPU.register.registers\[897\] vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
Xfanout845 net854 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_4
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _05354_ _05363_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__nand2_1
XFILLER_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1021 top0.CPU.register.registers\[399\] vssd1 vssd1 vccd1 vccd1 net3243 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net3365 _02396_ _04751_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__o21a_1
XFILLER_85_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08183__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1032 net78 vssd1 vssd1 vccd1 vccd1 net3254 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 top0.CPU.register.registers\[125\] vssd1 vssd1 vccd1 vccd1 net3232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 net891 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_2
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_4
Xhold1043 top0.CPU.register.registers\[76\] vssd1 vssd1 vccd1 vccd1 net3265 sky130_fd_sc_hd__dlygate4sd3_1
X_11347__999 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__inv_2
X_09797_ top0.CPU.internalMem.pcOut\[12\] _05280_ _05302_ vssd1 vssd1 vccd1 vccd1
+ _05303_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout844_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07804__C _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1076 top0.CPU.register.registers\[226\] vssd1 vssd1 vccd1 vccd1 net3298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 top0.CPU.register.registers\[1013\] vssd1 vssd1 vccd1 vccd1 net3287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 top0.CPU.register.registers\[405\] vssd1 vssd1 vccd1 vccd1 net3276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1098 top0.CPU.register.registers\[178\] vssd1 vssd1 vccd1 vccd1 net3320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08748_ _04686_ net316 net294 net2567 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__a22o_1
Xhold1087 top0.CPU.register.registers\[182\] vssd1 vssd1 vccd1 vccd1 net3309 sky130_fd_sc_hd__dlygate4sd3_1
X_08679_ net193 net698 net320 net299 net2594 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a32o_1
XANTENNA__09683__A1 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08486__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__C1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ net1382 _01329_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06436__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06249__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08789__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ net2003 _01950_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[804\]
+ sky130_fd_sc_hd__dfrtp_1
X_12242_ net1934 _01881_ net1054 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[735\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08946__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250__902 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__inv_2
XANTENNA__07749__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net1865 _01812_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10457__109 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__inv_2
XFILLER_77_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10006_ top0.CPU.internalMem.pcOut\[28\] net645 _05495_ vssd1 vssd1 vccd1 vccd1 _02205_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA__07714__C net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06280__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09123__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ net1649 _01596_ net972 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06032__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11888_ net1580 _01527_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08318__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ net2201 _02148_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1002\]
+ sky130_fd_sc_hd__dfrtp_1
X_06030_ top0.CPU.register.registers\[905\] top0.CPU.register.registers\[937\] top0.CPU.register.registers\[969\]
+ top0.CPU.register.registers\[1001\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02687_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06660__A1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08937__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07981_ _04127_ _04474_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__nor2_1
Xfanout119 net124 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
X_11034__686 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__inv_2
X_09720_ top0.CPU.internalMem.pcOut\[6\] net650 _05231_ vssd1 vssd1 vccd1 vccd1 _02183_
+ sky130_fd_sc_hd__o21a_1
X_06932_ top0.CPU.register.registers\[921\] top0.CPU.register.registers\[953\] top0.CPU.register.registers\[985\]
+ top0.CPU.register.registers\[1017\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03589_
+ sky130_fd_sc_hd__mux4_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07193__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net3383 top0.MISOtoMMIO\[2\] _05173_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06863_ _03507_ _03518_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06794_ net867 _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nor2_1
X_05814_ net744 _02470_ _02465_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09582_ _05122_ _05124_ top0.display.counter\[2\] vssd1 vssd1 vccd1 vccd1 _05126_
+ sky130_fd_sc_hd__a21o_1
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08602_ net3011 net329 net305 _04529_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a22o_1
X_08533_ _04717_ net408 net364 net2965 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05745_ net954 net950 net952 net947 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09114__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout258_A _04809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06023__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ _04681_ net395 net370 net2560 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a22o_1
X_07415_ _03406_ _04071_ _03405_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout425_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08395_ _04660_ net395 net378 net2870 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XFILLER_137_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _02730_ _03518_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_21_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_07_1133 vssd1 vssd1 vccd1 vccd1 team_07_1133/HI gpio_oeb[1] sky130_fd_sc_hd__conb_1
Xteam_07_1144 vssd1 vssd1 vccd1 vccd1 team_07_1144/HI gpio_out[10] sky130_fd_sc_hd__conb_1
Xteam_07_1166 vssd1 vssd1 vccd1 vccd1 team_07_1166/HI gpio_out[32] sky130_fd_sc_hd__conb_1
XANTENNA__08640__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ _03728_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__or2_1
Xteam_07_1177 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] team_07_1177/LO sky130_fd_sc_hd__conb_1
Xteam_07_1155 vssd1 vssd1 vccd1 vccd1 team_07_1155/HI gpio_out[21] sky130_fd_sc_hd__conb_1
Xteam_07_1188 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] team_07_1188/LO sky130_fd_sc_hd__conb_1
X_09016_ net3344 net350 _04801_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__a21o_1
X_10642__294 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__inv_2
XANTENNA_fanout794_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06228_ _02883_ _02884_ net731 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
Xhold151 top0.CPU.register.registers\[877\] vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 top0.CPU.register.registers\[456\] vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
X_06159_ _02814_ _02815_ net729 vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
Xhold140 top0.CPU.register.registers\[290\] vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07087__B _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold184 top0.CPU.register.registers\[869\] vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 top0.CPU.register.registers\[815\] vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 top0.CPU.register.registers\[70\] vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout631 _02418_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_2
Xfanout620 net623 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_4
X_09918_ _05400_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__and2_1
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_2
Xfanout653 net654 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_2
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout664 net667 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_2
X_10372__24 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__inv_2
Xfanout686 net687 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09849_ top0.CPU.internalMem.pcOut\[16\] net647 _05347_ _05350_ vssd1 vssd1 vccd1
+ vccd1 _02193_ sky130_fd_sc_hd__o22a_1
XANTENNA__07903__A1 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ net1503 _01450_ net1035 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[304\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06014__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08459__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ net1434 _01381_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[235\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__B _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08138__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11673_ net1365 _01312_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[166\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07419__A0 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06317__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ net1917 _01864_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[718\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09493__A _02355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net1848 _01795_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[649\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05724__A_N top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net1779 _01726_ net975 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[580\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06786__A1_N net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__B _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06005__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09004__Y _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10585__237 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__inv_2
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06556__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__A1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ net511 net181 net621 net428 net2773 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a32o_1
X_07200_ _03751_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__nand2_1
XANTENNA__08870__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ net457 _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626__278 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__inv_2
X_07062_ _02431_ _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or2_4
X_06013_ _02668_ _02669_ net728 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
XANTENNA__12574__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__A _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06820__A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479__131 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__inv_2
X_07964_ top0.CPU.intMem_out\[9\] net628 _04588_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_
+ sky130_fd_sc_hd__a22o_1
X_09703_ top0.CPU.internalMem.pcOut\[5\] _05207_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__or2_1
XANTENNA__09335__B1 _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07895_ _04432_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__and3_1
X_06915_ _03223_ _03224_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__nor2_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08689__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _03499_ _03500_ _03501_ _03502_ net760 net864 vssd1 vssd1 vccd1 vccd1 _03503_
+ sky130_fd_sc_hd__mux4_2
X_09634_ _04957_ _05162_ net662 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o21a_1
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06795__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ net632 _04631_ _05110_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout542_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout163_X net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ _03430_ _03431_ _03432_ _03433_ net765 net753 vssd1 vssd1 vccd1 vccd1 _03434_
+ sky130_fd_sc_hd__mux4_1
X_09496_ top0.MMIO.WBData_i\[19\] net140 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05728_ _02338_ _02380_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__nor2_2
X_08516_ net166 net679 net389 net365 net2397 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a32o_1
XANTENNA__07113__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08447_ net2914 net174 net374 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ net217 net706 net399 net383 net2704 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a32o_1
XANTENNA__09810__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ net482 _03953_ _03984_ _03841_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__a211o_1
X_10340_ net2244 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10271_ net3173 net120 net113 _05657_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ net1702 _01649_ net965 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[503\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout450 _02636_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06483__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout472 _02598_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout461 net466 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_2
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06235__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout494 net496 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12774_ net767 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08301__A1 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ net1417 _01364_ net958 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[218\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06312__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11656_ net1348 _01295_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[149\]
+ sky130_fd_sc_hd__dfrtp_1
X_11587_ net1279 _01226_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08604__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07407__A3 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06615__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold909 top0.CPU.register.registers\[894\] vssd1 vssd1 vccd1 vccd1 net3131 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06710__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__B1 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ net1900 _01847_ net1081 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[701\]
+ sky130_fd_sc_hd__dfrtp_1
X_10970__622 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__inv_2
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12139_ net1831 _01778_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[632\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09951__A top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06700_ _02579_ _02597_ _03356_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o21ai_2
XANTENNA__06226__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ _02554_ _03991_ _04336_ net448 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__o211a_1
XANTENNA__06777__S1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ _03286_ _03287_ net758 vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__mux2_1
XANTENNA__09096__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ _04991_ _04995_ _04996_ _04997_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.state_n\[1\]
+ sky130_fd_sc_hd__or4_1
X_11146__798 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__inv_2
X_06562_ _03217_ _03218_ net758 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
X_09281_ _02361_ top0.wishbone0.curr_state\[1\] top0.wishbone0.curr_state\[0\] _04941_
+ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XANTENNA__06529__S1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08301_ net2930 _04555_ net415 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
X_08232_ net504 net174 net684 net423 net2273 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a32o_1
X_06493_ net746 _03149_ _03142_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__a21oi_4
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_119_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ net204 net617 vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08056__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08094_ net515 net190 net699 net435 net2256 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a32o_1
X_07114_ net457 _03770_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__nand2_1
Xclkload60 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_8
Xclkload71 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_6
X_07045_ net519 _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1032_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_8
Xclkload82 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_16
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06909__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__A1 _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout492_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06465__S0 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ top0.CPU.register.registers\[166\] net566 net553 vssd1 vssd1 vccd1 vccd1
+ _04796_ sky130_fd_sc_hd__o21a_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07947_ top0.CPU.intMem_out\[12\] net626 _02768_ _02386_ net639 vssd1 vssd1 vccd1
+ vccd1 _04585_ sky130_fd_sc_hd__o221a_1
XFILLER_88_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout757_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ top0.CPU.intMem_out\[23\] net627 _04526_ net642 vssd1 vssd1 vccd1 vccd1 _04527_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _02516_ _05003_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__nand2_2
X_06829_ _03484_ _03485_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__nor2_1
XFILLER_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08196__B net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout924_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ top0.CPU.control.funct7\[1\] _05063_ net126 vssd1 vssd1 vccd1 vccd1 _01117_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09087__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ top0.MMIO.WBData_i\[23\] net137 vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_61_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11510_ net1202 _01149_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ net2182 _02129_ net984 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[983\]
+ sky130_fd_sc_hd__dfrtp_1
X_11441_ clknet_leaf_68_clk _01089_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08047__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire136 _05152_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06940__S1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06073__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954__606 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__inv_2
X_10323_ net2243 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09547__A0 top0.CPU.control.funct7\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10254_ _04938_ _05131_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__or2_1
X_10185_ top0.wishbone0.curr_state\[1\] top0.wishbone0.curr_state\[2\] _04942_ top0.wishbone0.curr_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_72_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_4
XANTENNA__06759__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10848__500 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__inv_2
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09078__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08825__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10093__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08286__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ net1400 _01347_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[201\]
+ sky130_fd_sc_hd__dfrtp_1
X_12688_ clknet_leaf_92_clk _02323_ net1082 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08038__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ net1331 _01278_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06931__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09946__A top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08053__A3 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__A2 top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 top0.CPU.register.registers\[797\] vssd1 vssd1 vccd1 vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold706 top0.CPU.register.registers\[507\] vssd1 vssd1 vccd1 vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 top0.CPU.register.registers\[728\] vssd1 vssd1 vccd1 vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07261__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09538__A0 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697__349 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__inv_2
Xhold739 top0.CPU.register.registers\[982\] vssd1 vssd1 vccd1 vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06695__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06370__A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09157__S net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _04581_ net3114 net355 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__mux2_1
X_07801_ net519 _03785_ _04456_ _04457_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__and4b_1
XANTENNA__07564__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ net196 net687 net325 net291 net2537 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__a32o_1
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05993_ top0.CPU.control.funct7\[0\] _02518_ _02649_ net581 vssd1 vssd1 vccd1 vccd1
+ _02650_ sky130_fd_sc_hd__a22o_2
X_07732_ _03582_ _03620_ _03618_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__o21ba_1
XANTENNA__05714__A top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _03563_ _04298_ _03484_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a21oi_1
X_06614_ net872 _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__and2_1
X_09402_ _05009_ net149 vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_36_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09333_ _04292_ net233 _04980_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a211o_1
XANTENNA__09069__A2 _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ net487 net531 net339 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__a21o_1
XANTENNA__08816__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06545_ net540 _02812_ _03200_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__nand3_1
XFILLER_61_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_126_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_138_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ _04916_ _04920_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__or2_1
XANTENNA__10084__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06545__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06476_ _02477_ _02496_ _02833_ _02869_ net543 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_134_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09195_ top0.display.state\[2\] _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and2_1
X_08215_ net3085 net423 _04700_ net508 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
X_08146_ net3131 net427 _04673_ net513 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout505_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ net2806 net433 _04661_ net492 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a22o_1
X_07028_ net747 _03684_ _03677_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07807__C net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout874_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold22 top0.CPU.register.registers\[10\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 top0.CPU.register.registers\[17\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06989__S1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08979_ _04556_ net698 _04790_ net260 net3320 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__a32o_1
Xhold55 top0.CPU.register.registers\[944\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 top0.CPU.register.registers\[2\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__B net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 top0.CPU.register.registers\[547\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 top0.CPU.register.registers\[680\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 top0.CPU.intMemAddr\[20\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 top0.CPU.register.registers\[996\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 top0.CPU.register.registers\[36\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net1682 _01629_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09701__B1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__A _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06610__S0 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_12611_ clknet_leaf_81_clk _02246_ net1112 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12542_ clknet_leaf_78_clk _02181_ net1107 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06279__C1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ net2165 _02112_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[966\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08283__A3 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ clknet_leaf_61_clk _01072_ net1100 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_8 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07243__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06677__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _04932_ net577 _05633_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__or3b_1
XANTENNA__07794__A2 _03882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10237_ net9 net653 net592 net3363 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__o22a_1
XFILLER_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09705__S net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1031 net1036 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__X _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1042 net1044 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
X_10168_ top0.display.delayctr\[28\] _04970_ _05604_ vssd1 vssd1 vccd1 vccd1 _05626_
+ sky130_fd_sc_hd__or3_1
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
Xfanout1097 net1106 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__buf_2
X_10099_ top0.display.delayctr\[15\] _05566_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__nand2_1
Xfanout1086 net1087 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
Xfanout1075 net1077 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06601__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_108_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08259__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06330_ _02985_ _02986_ net732 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__mux2_1
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__A3 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06261_ _02916_ _02917_ net724 vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08000_ _04292_ net233 net228 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_116_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06192_ net739 _02848_ net742 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__o21ai_1
Xhold536 top0.CPU.register.registers\[936\] vssd1 vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 top0.CPU.register.registers\[308\] vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09395__B _05006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 top0.CPU.register.registers\[214\] vssd1 vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 top0.CPU.register.registers\[321\] vssd1 vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 top0.CPU.register.registers\[556\] vssd1 vssd1 vccd1 vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ top0.CPU.internalMem.pcOut\[24\] _05426_ vssd1 vssd1 vccd1 vccd1 _05445_
+ sky130_fd_sc_hd__or2_1
Xhold547 top0.CPU.register.registers\[436\] vssd1 vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 top0.CPU.register.registers\[438\] vssd1 vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ top0.CPU.register.registers\[233\] net573 net559 vssd1 vssd1 vccd1 vccd1
+ _04769_ sky130_fd_sc_hd__o21a_1
X_09882_ top0.CPU.internalMem.pcOut\[19\] top0.CPU.internalMem.pcOut\[18\] _05359_
+ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__and3_1
XANTENNA__07537__A2 _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05891__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1203 top0.MMIO.WBData_i\[29\] vssd1 vssd1 vccd1 vccd1 net3425 sky130_fd_sc_hd__dlygate4sd3_1
X_08833_ net212 net3144 net355 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__mux2_1
Xhold1214 top0.CPU.internalMem.storeCt\[0\] vssd1 vssd1 vccd1 vccd1 net3436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout288_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ net946 net688 _04734_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__nand3_4
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05976_ _02629_ _02630_ _02631_ _02632_ net725 net776 vssd1 vssd1 vccd1 vccd1 _02633_
+ sky130_fd_sc_hd__mux4_2
XFILLER_73_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07715_ net341 _04131_ _04132_ net442 _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o221a_1
XANTENNA__08498__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ _02396_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__nand2_1
XANTENNA__09695__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161__813 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__inv_2
XFILLER_53_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07646_ _03895_ _04050_ _04161_ net441 _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__o221a_1
XFILLER_53_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout622_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ net449 net530 net339 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06528_ net865 _03180_ net860 vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o21ai_1
X_11202__854 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__inv_2
X_09316_ top0.display.delayctr\[12\] top0.display.delayctr\[13\] top0.display.delayctr\[14\]
+ top0.display.delayctr\[15\] vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__or4_1
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ top0.CPU.internalMem.pcOut\[2\] _04908_ net609 vssd1 vssd1 vccd1 vccd1 _04909_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06459_ _02497_ _02834_ net541 vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08670__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ net167 net3123 net250 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__mux2_1
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ net2919 net188 net430 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09525__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ top0.CPU.internalMem.pcOut\[30\] _05509_ vssd1 vssd1 vccd1 vccd1 _05510_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__05906__X _02563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__B _03092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08489__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ net1665 _01612_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07272__C net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810__462 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07161__A0 _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_12525_ net2217 _02164_ net958 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1018\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08661__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__S0 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12456_ net2148 _02095_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[949\]
+ sky130_fd_sc_hd__dfrtp_1
X_12387_ net2079 _02026_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[880\]
+ sky130_fd_sc_hd__dfrtp_1
X_11407_ clknet_leaf_87_clk _01055_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08413__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07216__B2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10378__30 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__inv_2
XFILLER_97_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05873__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06822__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05830_ top0.CPU.register.registers\[402\] top0.CPU.register.registers\[434\] top0.CPU.register.registers\[466\]
+ top0.CPU.register.registers\[498\] net846 net811 vssd1 vssd1 vccd1 vccd1 _02487_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_94_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05761_ top0.CPU.Op\[3\] _02378_ _02381_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__or3_1
XFILLER_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07500_ _02788_ _02789_ net528 vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__and3_1
XANTENNA__12599__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05692_ top0.CPU.internalMem.pcOut\[13\] vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__inv_2
X_08480_ net173 net615 net390 net371 net2501 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a32o_1
X_07431_ net342 _04074_ _04075_ _04086_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_46_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06807__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07362_ _02699_ net525 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__and2_1
XANTENNA__09444__A2 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06313_ net777 _02965_ _02968_ _02969_ net772 vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__o221ai_4
X_09101_ _04693_ net269 net251 net2712 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__a22o_1
XANTENNA__06889__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08652__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07293_ net536 net447 net467 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__mux2_1
XANTENNA__07455__A1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09032_ net182 net3311 net351 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06244_ _02899_ _02900_ net731 vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__mux2_1
XANTENNA__07919__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__B _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 top0.CPU.register.registers\[966\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ _02812_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__and2_1
Xhold311 top0.CPU.register.registers\[34\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 top0.CPU.register.registers\[116\] vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 top0.CPU.register.registers\[228\] vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__A2 _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 top0.CPU.register.registers\[700\] vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold366 top0.CPU.register.registers\[95\] vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 top0.CPU.register.registers\[40\] vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 net49 vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 top0.CPU.register.registers\[383\] vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
X_10753__405 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__inv_2
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
X_09934_ top0.CPU.internalMem.pcOut\[23\] net646 _05425_ _05428_ vssd1 vssd1 vccd1
+ vccd1 _02200_ sky130_fd_sc_hd__o22a_1
Xhold388 top0.CPU.register.registers\[596\] vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06969__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout802 net805 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_4
Xfanout824 net825 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout857 top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09865_ _05345_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nor2_1
Xfanout846 net854 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold1000 top0.CPU.register.registers\[180\] vssd1 vssd1 vccd1 vccd1 net3222 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__buf_4
XFILLER_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1220_A top0.CPU.intMem_out\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06813__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 top0.CPU.decoder.instruction\[18\] vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_8
X_08816_ net193 net675 _04736_ net287 top0.CPU.register.registers\[301\] vssd1 vssd1
+ vccd1 vccd1 _04751_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout572_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1011 net73 vssd1 vssd1 vccd1 vccd1 net3233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 top0.display.dataforOutput\[9\] vssd1 vssd1 vccd1 vccd1 net3255 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 top0.CPU.register.registers\[78\] vssd1 vssd1 vccd1 vccd1 net3244 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 net885 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_2
X_09796_ top0.CPU.internalMem.pcOut\[12\] _05280_ net240 vssd1 vssd1 vccd1 vccd1 _05302_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07930__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1066 top0.CPU.register.registers\[424\] vssd1 vssd1 vccd1 vccd1 net3288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06194__A1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1055 top0.CPU.register.registers\[820\] vssd1 vssd1 vccd1 vccd1 net3277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07804__D net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1044 top0.CPU.register.registers\[860\] vssd1 vssd1 vccd1 vccd1 net3266 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net198 net623 net325 net295 net2738 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 top0.CPU.register.registers\[176\] vssd1 vssd1 vccd1 vccd1 net3310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 top0.CPU.register.registers\[285\] vssd1 vssd1 vccd1 vccd1 net3299 sky130_fd_sc_hd__dlygate4sd3_1
X_05959_ net584 _02614_ _02615_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout837_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1099 top0.CPU.register.registers\[1018\] vssd1 vssd1 vccd1 vccd1 net3321 sky130_fd_sc_hd__dlygate4sd3_1
X_08678_ _04667_ net316 net298 net2805 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a22o_1
X_07629_ net489 _04040_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__nand2_1
XANTENNA__08486__A3 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__C_N top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08238__A3 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08643__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08424__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ net2002 _01949_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[803\]
+ sky130_fd_sc_hd__dfrtp_1
X_12241_ net1933 _01880_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[734\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10202__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ net1864 _01811_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330__982 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__inv_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10496__148 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__inv_2
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10005_ _05490_ _05491_ _05494_ _05110_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07851__X _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06280__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537__189 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__inv_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__A0 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ net1648 _01595_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08477__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06032__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07685__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ net1579 _01526_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08229__A3 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__C1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06119__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08634__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ net2200 _02147_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1001\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07988__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12439_ net2131 _02078_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[932\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08401__A3 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ net719 net505 net173 net547 net2340 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a32o_1
X_06931_ top0.CPU.register.registers\[793\] top0.CPU.register.registers\[825\] top0.CPU.register.registers\[857\]
+ top0.CPU.register.registers\[889\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03588_
+ sky130_fd_sc_hd__mux4_1
X_09650_ net3372 top0.MISOtoMMIO\[1\] _05173_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__mux2_1
XANTENNA__09392__C _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07193__B _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__inv_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08601_ net3182 net330 net314 _04523_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a22o_1
X_06793_ _03448_ _03449_ net766 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
X_05813_ _02466_ _02467_ _02468_ _02469_ net734 net781 vssd1 vssd1 vccd1 vccd1 _02470_
+ sky130_fd_sc_hd__mux4_2
X_09581_ net605 _05123_ _05125_ _05121_ net2901 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_124_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05744_ net954 net950 net952 net946 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__or4b_1
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08532_ _04716_ net400 net363 net2779 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a22o_1
XANTENNA__08468__A3 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06023__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _04680_ net385 net369 net2714 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
XANTENNA__06537__B _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ _03364_ _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__a21o_1
XANTENNA__08873__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__A2 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05782__S0 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08394_ _04659_ net386 net377 net2570 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout320_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07345_ _02730_ _03518_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08625__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1134 vssd1 vssd1 vccd1 vccd1 team_07_1134/HI gpio_oeb[3] sky130_fd_sc_hd__conb_1
Xteam_07_1145 vssd1 vssd1 vccd1 vccd1 team_07_1145/HI gpio_out[11] sky130_fd_sc_hd__conb_1
XANTENNA__07979__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05868__S net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ net484 _03719_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__or2_4
XFILLER_12_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11273__925 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__inv_2
XANTENNA__06636__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1167 vssd1 vssd1 vccd1 vccd1 team_07_1167/HI gpio_out[33] sky130_fd_sc_hd__conb_1
X_06227_ top0.CPU.register.registers\[278\] top0.CPU.register.registers\[310\] top0.CPU.register.registers\[342\]
+ top0.CPU.register.registers\[374\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02884_
+ sky130_fd_sc_hd__mux4_1
Xteam_07_1178 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] team_07_1178/LO sky130_fd_sc_hd__conb_1
Xteam_07_1156 vssd1 vssd1 vccd1 vccd1 team_07_1156/HI gpio_out[22] sky130_fd_sc_hd__conb_1
X_09015_ top0.CPU.register.registers\[152\] net568 net207 net613 vssd1 vssd1 vccd1
+ vccd1 _04801_ sky130_fd_sc_hd__o211a_1
Xteam_07_1189 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] team_07_1189/LO sky130_fd_sc_hd__conb_1
XANTENNA__09050__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 top0.CPU.register.registers\[584\] vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07936__X _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06158_ top0.CPU.register.registers\[528\] top0.CPU.register.registers\[560\] top0.CPU.register.registers\[592\]
+ top0.CPU.register.registers\[624\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02815_
+ sky130_fd_sc_hd__mux4_1
X_11314__966 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__inv_2
Xhold141 top0.CPU.register.registers\[194\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 top0.CPU.register.registers\[674\] vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 top0.CPU.register.registers\[79\] vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 top0.CPU.register.registers\[111\] vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
X_06089_ net784 _02743_ net738 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a21o_1
Xhold174 top0.CPU.register.registers\[832\] vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 top0.CPU.register.registers\[581\] vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ _05387_ _05392_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a21o_1
Xfanout632 _02418_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net677 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_2
XANTENNA_fanout954_A top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout643 _02382_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_2
XANTENNA__08156__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout687 net688 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
Xfanout698 net700 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ net236 _05348_ _05349_ net647 vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__o31ai_1
XFILLER_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ net857 net643 net590 _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ net1502 _01449_ net1047 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05914__B2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208__860 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__inv_2
X_11741_ net1433 _01380_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[234\]
+ sky130_fd_sc_hd__dfrtp_1
X_10881__533 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__inv_2
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06014__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ net1364 _01311_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[165\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
X_10922__574 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__inv_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08092__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ net1916 _01863_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[717\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12155_ net1847 _01794_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
X_12086_ net1778 _01725_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[579\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07233__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ net1631 _01578_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[432\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06005__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__A1 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257__909 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__inv_2
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_07130_ net518 net539 net475 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11001__653 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__inv_2
XANTENNA__08083__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08622__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06092__B _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07061_ _02428_ _03713_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__or2_1
X_06012_ top0.CPU.register.registers\[518\] top0.CPU.register.registers\[550\] top0.CPU.register.registers\[582\]
+ top0.CPU.register.registers\[614\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02669_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09478__A_N top0.MMIO.WBData_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05717__A top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ net561 _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_79_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09702_ top0.CPU.internalMem.pcOut\[5\] _05207_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nand2_1
X_06914_ _03488_ _03570_ _03566_ _03564_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__o211a_1
X_07894_ net3287 net549 net501 _04540_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XANTENNA__09886__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07897__A1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06845_ top0.CPU.register.registers\[267\] top0.CPU.register.registers\[299\] top0.CPU.register.registers\[331\]
+ top0.CPU.register.registers\[363\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03502_
+ sky130_fd_sc_hd__mux4_1
X_09633_ _02758_ _02766_ _05150_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__o21ba_2
XANTENNA__08689__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__inv_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout270_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08515_ net213 net680 net390 net365 net2849 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a32o_1
X_06776_ top0.CPU.register.registers\[526\] top0.CPU.register.registers\[558\] top0.CPU.register.registers\[590\]
+ top0.CPU.register.registers\[622\] net921 net887 vssd1 vssd1 vccd1 vccd1 _03433_
+ sky130_fd_sc_hd__mux4_1
X_10865__517 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__inv_2
X_09495_ top0.MMIO.WBData_i\[12\] net137 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05727_ _02339_ top0.CPU.Op\[2\] _02370_ _02371_ top0.CPU.Op\[5\] vssd1 vssd1 vccd1
+ vccd1 _02384_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout535_A _03173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ net3241 net177 net374 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__mux2_1
XFILLER_51_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906__558 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__inv_2
X_08377_ net179 net708 net401 net383 net2400 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_137_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout702_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ net244 _03972_ _03976_ net448 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08613__A3 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07259_ _03114_ _03915_ _03094_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09023__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432__84 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__inv_2
X_10270_ net144 _05156_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__nand2_1
XANTENNA__09594__A _02614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759__411 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__inv_2
XANTENNA__08377__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout440 _04637_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_6
XANTENNA__06483__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _02636_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_2
Xfanout462 net464 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
Xfanout484 _02555_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_2
XANTENNA__07337__A0 _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout473 net475 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05914__X _02571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06235__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_2
XFILLER_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12773_ net767 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06312__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11724_ net1416 _01363_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[217\]
+ sky130_fd_sc_hd__dfrtp_1
X_11655_ net1347 _01294_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09488__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11586_ net1278 _01225_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08065__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09014__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ net1899 _01846_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[700\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12138_ net1830 _01777_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[631\]
+ sky130_fd_sc_hd__dfrtp_1
X_12069_ net1761 _01708_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[562\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_10552__204 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__inv_2
XFILLER_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06226__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06630_ top0.CPU.register.registers\[771\] top0.CPU.register.registers\[803\] top0.CPU.register.registers\[835\]
+ top0.CPU.register.registers\[867\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03287_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_121_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08828__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ top0.CPU.register.registers\[17\] top0.CPU.register.registers\[49\] top0.CPU.register.registers\[81\]
+ top0.CPU.register.registers\[113\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03218_
+ sky130_fd_sc_hd__mux4_1
XFILLER_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08300_ net2842 _04550_ net416 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
X_09280_ _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__inv_2
XANTENNA__06303__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06492_ _03145_ _03148_ net753 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux2_1
XFILLER_33_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08231_ net504 net177 net683 net423 net2344 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a32o_1
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08162_ net2931 net426 _04681_ net500 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08056__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08093_ net514 net194 net697 net435 net2658 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a32o_1
X_07113_ net474 net538 _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__o21ai_1
Xclkload61 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_8
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_2
X_07044_ _03686_ _03700_ net583 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_132_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload72 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_8
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload83 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_4
XANTENNA__08359__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload94 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_2
XFILLER_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06465__S1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net176 net694 _04795_ net260 net3143 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__a32o_1
X_07946_ net561 _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__or2_1
XANTENNA__09308__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__A _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ net561 _04524_ _04525_ net625 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06828_ _03467_ _03468_ _03483_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__and3_1
X_09616_ top0.display.dataforOutput\[6\] net604 net658 net3304 _05149_ vssd1 vssd1
+ vccd1 vccd1 _01137_ sky130_fd_sc_hd__a221o_1
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_48_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05976__S0 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09547_ top0.CPU.control.funct7\[0\] _05082_ net125 vssd1 vssd1 vccd1 vccd1 _01116_
+ sky130_fd_sc_hd__mux2_1
X_06759_ top0.CPU.register.registers\[911\] top0.CPU.register.registers\[943\] top0.CPU.register.registers\[975\]
+ top0.CPU.register.registers\[1007\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03416_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__Y _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279__931 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__inv_2
XANTENNA__09087__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ top0.MMIO.WBData_i\[15\] net148 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_61_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11606__RESET_B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08429_ net2925 _04522_ net374 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
X_11440_ clknet_leaf_68_clk _01088_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08047__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06217__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__08598__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10322_ net2231 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__clkbuf_1
X_10993__645 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__inv_2
XFILLER_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08432__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ _04941_ _05639_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__nor2_1
XANTENNA__10263__A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B _03130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ top0.wishbone0.curr_state\[1\] top0.wishbone0.curr_state\[2\] _04942_ top0.wishbone0.curr_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__and4bb_1
XFILLER_94_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08770__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout292 _04749_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
Xfanout281 _04755_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_4
XFILLER_94_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout270 net272 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08387__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08522__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05967__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06188__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08286__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__A3 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10928__580 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__inv_2
X_11707_ net1399 _01346_ net1009 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[200\]
+ sky130_fd_sc_hd__dfrtp_1
X_12687_ clknet_leaf_91_clk _02322_ net1108 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06392__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08038__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ net1330 _01277_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06049__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11569_ net1261 _01208_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05966__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 top0.CPU.register.registers\[502\] vssd1 vssd1 vccd1 vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 top0.CPU.register.registers\[529\] vssd1 vssd1 vccd1 vccd1 net2940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 top0.CPU.register.registers\[523\] vssd1 vssd1 vccd1 vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
X_11072__724 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__inv_2
XANTENNA__06695__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__A3 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08780_ net201 net684 net319 net291 net2410 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__a32o_1
X_07800_ _03006_ _03022_ _03701_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o21a_1
XANTENNA__08761__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113__765 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__inv_2
XANTENNA__06797__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05992_ _02643_ _02648_ net743 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_4
X_07731_ _03715_ _04367_ _04379_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__o31ai_1
XFILLER_38_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05714__B top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ _04016_ _04044_ _04295_ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__or4_1
XANTENNA__08513__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06613_ top0.CPU.register.registers\[901\] top0.CPU.register.registers\[933\] top0.CPU.register.registers\[965\]
+ top0.CPU.register.registers\[997\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03270_
+ sky130_fd_sc_hd__mux4_1
X_09401_ net149 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__inv_2
XFILLER_111_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07593_ _03361_ _03363_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08277__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09332_ _04619_ _04623_ _04631_ _04976_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__or4_1
X_06544_ net540 _02812_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__and3_1
XANTENNA__08816__A3 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06826__A _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09263_ _04918_ _04920_ _04922_ _04924_ _04897_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__o2111ai_1
X_06475_ _03117_ _03130_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_134_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10680__332 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__inv_2
X_09194_ top0.display.state\[1\] top0.display.state\[0\] vssd1 vssd1 vccd1 vccd1 _04857_
+ sky130_fd_sc_hd__nor2_1
X_08214_ net223 net687 vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__and2_1
X_10977__629 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08145_ net212 net624 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__and2_1
XANTENNA__09777__A1 _03989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout400_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721__373 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__inv_2
X_08076_ net152 net690 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and2_1
X_07027_ _03680_ _03683_ net754 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__mux2_1
X_10402__54 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__inv_2
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07807__D net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 top0.CPU.register.registers\[19\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 top0.CPU.register.registers\[24\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 top0.CPU.register.registers\[940\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ top0.CPU.register.registers\[178\] net572 net559 vssd1 vssd1 vccd1 vccd1
+ _04790_ sky130_fd_sc_hd__o21a_1
Xhold56 top0.CPU.register.registers\[6\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 top0.CPU.register.registers\[822\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 top0.CPU.register.registers\[943\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 top0.CPU.register.registers\[236\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07929_ top0.CPU.intMem_out\[15\] net625 _02513_ _02386_ net638 vssd1 vssd1 vccd1
+ vccd1 _04570_ sky130_fd_sc_hd__o221a_1
Xhold89 top0.CPU.register.registers\[496\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05971__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05949__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06610__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ clknet_leaf_80_clk _02245_ net1113 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06736__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06295__X _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08268__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ clknet_leaf_78_clk _02180_ net1115 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10258__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ net2164 _02111_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[965\]
+ sky130_fd_sc_hd__dfrtp_1
X_11423_ clknet_leaf_60_clk _01071_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11056__708 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__inv_2
XFILLER_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06126__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__A1 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06471__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06677__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ net3327 net117 net111 _05629_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a22o_1
X_10236_ net8 net653 net592 net3446 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__o22a_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1021 net1056 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
Xfanout1010 net1011 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08743__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_2
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
Xfanout1032 net1036 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
X_10167_ _04957_ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__or2_1
Xfanout1065 net1088 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_2
Xfanout1098 net1100 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10098_ _04969_ _05548_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__or2_1
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_2
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06601__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06646__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664__316 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__inv_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06260_ top0.CPU.register.registers\[25\] top0.CPU.register.registers\[57\] top0.CPU.register.registers\[89\]
+ top0.CPU.register.registers\[121\] net825 net789 vssd1 vssd1 vccd1 vccd1 _02917_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705__357 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__inv_2
XANTENNA__06117__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06191_ _02846_ _02847_ net731 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
Xhold526 top0.CPU.register.registers\[595\] vssd1 vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold504 top0.CPU.register.registers\[606\] vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 top0.CPU.register.registers\[89\] vssd1 vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold559 net50 vssd1 vssd1 vccd1 vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08982__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ top0.CPU.internalMem.pcOut\[24\] _05426_ vssd1 vssd1 vccd1 vccd1 _05444_
+ sky130_fd_sc_hd__nand2_1
Xhold537 top0.CPU.register.registers\[954\] vssd1 vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 top0.CPU.register.registers\[729\] vssd1 vssd1 vccd1 vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
X_08901_ net720 net182 _04768_ net283 net3348 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__a32o_1
X_10558__210 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ _05377_ _05378_ net239 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a21o_1
XANTENNA__08734__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ net151 net3046 net355 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__mux2_1
Xhold1215 net61 vssd1 vssd1 vccd1 vccd1 net3437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1204 top0.display.delayctr\[25\] vssd1 vssd1 vccd1 vccd1 net3426 sky130_fd_sc_hd__dlygate4sd3_1
X_05975_ top0.CPU.register.registers\[260\] top0.CPU.register.registers\[292\] top0.CPU.register.registers\[324\]
+ top0.CPU.register.registers\[356\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02632_
+ sky130_fd_sc_hd__mux4_1
X_08763_ net155 net617 net314 net294 net2492 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_127_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout183_A _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07714_ _02962_ net521 net446 vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__or3_1
X_08694_ top0.CPU.decoder.instruction\[11\] _04668_ vssd1 vssd1 vccd1 vccd1 _04743_
+ sky130_fd_sc_hd__nor2_1
XFILLER_53_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout1092_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ _02769_ _03463_ net445 _04299_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout448_A _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A _04798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05731__Y _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ _03364_ _03382_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06527_ net752 _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nor2_1
X_09315_ top0.display.delayctr\[8\] top0.display.delayctr\[9\] top0.display.delayctr\[10\]
+ top0.display.delayctr\[11\] vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__or4_1
X_11241__893 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__inv_2
XANTENNA__06356__S0 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ top0.CPU.intMemAddr\[2\] _04623_ net769 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06458_ _03096_ net536 vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06990__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ net171 net669 _04848_ net249 net3221 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a32o_1
X_06389_ _03042_ _03043_ _03044_ _03045_ net765 net753 vssd1 vssd1 vccd1 vccd1 _03046_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__08422__A1 _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ net2729 net190 net431 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
X_08059_ net952 net950 net954 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_56_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_103_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08710__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net589 _04483_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a21o_1
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11692__RESET_B net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05922__X _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09150__A2 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net1664 _01611_ net988 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06595__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07161__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ net2216 _02163_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1017\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08661__A1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999__651 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__inv_2
XANTENNA__06898__S1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06472__Y _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ net2147 _02094_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[948\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06672__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ net2078 _02025_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[879\]
+ sky130_fd_sc_hd__dfrtp_1
X_11406_ clknet_leaf_87_clk _01054_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06405__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08177__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ _02359_ top0.wishbone0.prev_BUSY_O net655 vssd1 vssd1 vccd1 vccd1 _05647_
+ sky130_fd_sc_hd__and3_1
X_10393__45 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__inv_2
XANTENNA__06822__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05760_ top0.CPU.Op\[3\] net640 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__nor2_1
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11184__836 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__inv_2
XANTENNA__09677__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09141__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05691_ net784 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__inv_2
X_11225__877 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__inv_2
X_07430_ net452 _03933_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_46_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07361_ _03542_ _03558_ _03967_ net344 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a31o_1
XANTENNA__08101__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12568__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06312_ net727 _02966_ net736 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a21o_1
X_09100_ _04692_ net553 _04825_ net252 net3200 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a32o_1
XANTENNA__06889__S1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09031_ net187 net3112 net351 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__mux2_1
X_11078__730 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__inv_2
XFILLER_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07292_ net480 _03754_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o21a_1
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06243_ top0.CPU.register.registers\[24\] top0.CPU.register.registers\[56\] top0.CPU.register.registers\[88\]
+ top0.CPU.register.registers\[120\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02900_
+ sky130_fd_sc_hd__mux4_1
XFILLER_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold301 top0.CPU.register.registers\[458\] vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
X_06174_ net581 _02813_ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__o21ai_4
XANTENNA__12150__RESET_B net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold334 top0.CPU.register.registers\[457\] vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 top0.CPU.intMemAddr\[22\] vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
X_11119__771 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__inv_2
Xhold312 top0.CPU.register.registers\[216\] vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06510__S0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold378 top0.CPU.register.registers\[809\] vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 top0.CPU.register.registers\[366\] vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 top0.CPU.register.registers\[726\] vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top0.CPU.register.registers\[161\] vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout814 net819 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_2
XFILLER_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09933_ net235 _05426_ _05427_ net646 vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__o31ai_1
Xfanout803 net805 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08530__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 top0.CPU.register.registers\[470\] vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
X_10792__444 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__inv_2
Xfanout825 net834 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout847 net849 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_4
XFILLER_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ top0.CPU.internalMem.pcOut\[16\] _05343_ _05353_ vssd1 vssd1 vccd1 vccd1
+ _05364_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout398_A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_6
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07654__B net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net840 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_4
Xhold1012 top0.CPU.register.registers\[394\] vssd1 vssd1 vccd1 vccd1 net3234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1105_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08183__A3 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 net90 vssd1 vssd1 vccd1 vccd1 net3245 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _04719_ net316 net286 net2895 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__a22o_1
Xhold1001 top0.CPU.register.registers\[849\] vssd1 vssd1 vccd1 vccd1 net3223 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 top0.CPU.decoder.instruction\[17\] vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06813__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09795_ _05294_ _05297_ _05299_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__nor3_1
Xhold1056 top0.CPU.register.registers\[114\] vssd1 vssd1 vccd1 vccd1 net3278 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1067 top0.CPU.register.registers\[386\] vssd1 vssd1 vccd1 vccd1 net3289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 top0.CPU.register.registers\[156\] vssd1 vssd1 vccd1 vccd1 net3256 sky130_fd_sc_hd__dlygate4sd3_1
X_10833__485 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__inv_2
Xhold1045 top0.CPU.register.registers\[241\] vssd1 vssd1 vccd1 vccd1 net3267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 top0.CPU.register.registers\[138\] vssd1 vssd1 vccd1 vccd1 net3311 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net201 net620 _04747_ net295 net3332 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a32o_1
X_05958_ top0.CPU.decoder.instruction\[8\] _02448_ _02535_ net822 net583 vssd1 vssd1
+ vccd1 vccd1 _02615_ sky130_fd_sc_hd__a221o_1
Xhold1078 net48 vssd1 vssd1 vccd1 vccd1 net3300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08677_ net196 net697 net325 net299 net2526 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a32o_1
XANTENNA__06577__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05889_ top0.CPU.register.registers\[387\] top0.CPU.register.registers\[419\] top0.CPU.register.registers\[451\]
+ top0.CPU.register.registers\[483\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02546_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08340__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06286__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ _04283_ _04284_ net448 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ _04193_ _04203_ _04215_ _04175_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__o31ai_2
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08705__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ top0.CPU.internalMem.pcOut\[12\] top0.CPU.internalMem.pcOut\[11\] _04890_
+ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__or3_1
XANTENNA__06225__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ net1932 _01879_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[733\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08946__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ net1863 _01810_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06501__S0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05917__X _02574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold890 top0.CPU.register.registers\[139\] vssd1 vssd1 vccd1 vccd1 net3112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07845__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10004_ _05492_ _05493_ net645 vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09123__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07134__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ net1647 _01594_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[448\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12555__CLK clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11886_ net1578 _01525_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[379\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10438__90 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__inv_2
X_12507_ net2199 _02146_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1000\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06740__S0 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12438_ net2130 _02077_ net988 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[931\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08937__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10776__428 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__inv_2
X_12369_ net2061 _02008_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[862\]
+ sky130_fd_sc_hd__dfrtp_1
X_10520__172 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07474__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ _03585_ _03586_ net758 vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817__469 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__inv_2
X_06861_ _03512_ _03517_ net747 vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__mux2_4
XFILLER_95_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08600_ net2976 net329 net306 _04517_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a22o_1
X_05812_ top0.CPU.register.registers\[275\] top0.CPU.register.registers\[307\] top0.CPU.register.registers\[339\]
+ top0.CPU.register.registers\[371\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02469_
+ sky130_fd_sc_hd__mux4_1
X_06792_ top0.CPU.register.registers\[524\] top0.CPU.register.registers\[556\] top0.CPU.register.registers\[588\]
+ top0.CPU.register.registers\[620\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03449_
+ sky130_fd_sc_hd__mux4_1
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09580_ _05124_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05743_ net575 _02394_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__nand2_1
XANTENNA__09114__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08531_ _04715_ net396 net362 net2647 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a22o_1
XANTENNA__07125__A1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08322__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08462_ _04679_ net395 net370 net2750 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07413_ _03405_ _03406_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__and2b_1
XFILLER_51_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout146_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__Y _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ _04658_ net385 net377 net2509 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XANTENNA__05782__S1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ net486 _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08625__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1135 vssd1 vssd1 vccd1 vccd1 team_07_1135/HI gpio_oeb[4] sky130_fd_sc_hd__conb_1
X_07275_ net450 _03835_ _03925_ _03849_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a31o_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_07_1179 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] team_07_1179/LO sky130_fd_sc_hd__conb_1
Xteam_07_1146 vssd1 vssd1 vccd1 vccd1 team_07_1146/HI gpio_out[12] sky130_fd_sc_hd__conb_1
XANTENNA_fanout1055_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout313_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06731__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06226_ top0.CPU.register.registers\[406\] top0.CPU.register.registers\[438\] top0.CPU.register.registers\[470\]
+ top0.CPU.register.registers\[502\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02883_
+ sky130_fd_sc_hd__mux4_1
Xteam_07_1168 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] team_07_1168/LO sky130_fd_sc_hd__conb_1
Xteam_07_1157 vssd1 vssd1 vccd1 vccd1 team_07_1157/HI gpio_out[23] sky130_fd_sc_hd__conb_1
X_09014_ net208 net613 _04800_ net349 net3215 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__a32o_1
XANTENNA__08389__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06045__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 top0.CPU.register.registers\[880\] vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
X_06157_ top0.CPU.register.registers\[656\] top0.CPU.register.registers\[688\] top0.CPU.register.registers\[720\]
+ top0.CPU.register.registers\[752\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02814_
+ sky130_fd_sc_hd__mux4_1
Xhold142 top0.CPU.register.registers\[836\] vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 top0.CPU.register.registers\[163\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08928__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 top0.CPU.register.registers\[192\] vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold186 top0.CPU.register.registers\[837\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
X_06088_ net729 _02744_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__and2_1
Xhold164 top0.CPU.register.registers\[864\] vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 top0.CPU.register.registers\[579\] vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07039__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_4
Xfanout633 net634 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_2
X_09916_ _05386_ _05399_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__nand2_1
Xfanout600 _04859_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_2
XFILLER_59_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold197 net107 vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout655 _05646_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_2
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_2
Xfanout644 _02379_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
Xfanout688 net689 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
Xfanout677 _04704_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_8
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout947_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ top0.CPU.internalMem.pcOut\[15\] _05325_ top0.CPU.internalMem.pcOut\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09778_ top0.CPU.Op\[6\] top0.CPU.decoder.instruction\[7\] _02448_ _02518_ top0.CPU.control.funct7\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__a32o_1
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_29_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ net946 net624 _04734_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand3_4
XFILLER_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11740_ net1432 _01379_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[233\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06728__B _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ net1363 _01310_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[164\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08435__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463__115 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__inv_2
XANTENNA__08092__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12223_ net1915 _01862_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[716\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ net1846 _01793_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504__156 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363__15 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__inv_2
X_12085_ net1777 _01724_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[578\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08552__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11938_ net1630 _01577_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[431\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11869_ net1561 _01508_ net1024 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[362\]
+ sky130_fd_sc_hd__dfrtp_1
X_11296__948 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__inv_2
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11040__692 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__inv_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07060_ _03038_ _03669_ _03707_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06713__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06011_ top0.CPU.register.registers\[646\] top0.CPU.register.registers\[678\] top0.CPU.register.registers\[710\]
+ top0.CPU.register.registers\[742\] net830 net796 vssd1 vssd1 vccd1 vccd1 _02668_
+ sky130_fd_sc_hd__mux4_1
X_11337__989 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__inv_2
XANTENNA__11795__RESET_B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06660__Y _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__A3 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _05199_ _05204_ _05212_ net237 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__o31a_1
X_07962_ _04044_ net232 net227 vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__and3_1
XANTENNA__05717__B top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ _03505_ _03521_ _03541_ _03567_ _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__o41a_1
X_07893_ net723 net204 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and2_1
XANTENNA__08543__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ net3094 net605 net659 top0.display.dataforOutput\[11\] _05161_ vssd1 vssd1
+ vccd1 vccd1 _01141_ sky130_fd_sc_hd__a221o_1
X_06844_ top0.CPU.register.registers\[395\] top0.CPU.register.registers\[427\] top0.CPU.register.registers\[459\]
+ top0.CPU.register.registers\[491\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03501_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05733__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ net590 _02579_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__nor2_1
X_08514_ net169 net685 net402 net368 net2418 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a32o_1
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06775_ top0.CPU.register.registers\[654\] top0.CPU.register.registers\[686\] top0.CPU.register.registers\[718\]
+ top0.CPU.register.registers\[750\] net920 net887 vssd1 vssd1 vccd1 vccd1 _03432_
+ sky130_fd_sc_hd__mux4_1
X_09494_ top0.MMIO.WBData_i\[22\] net149 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__and2_1
X_05726_ _02378_ _02381_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout430_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net2933 net220 net375 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
X_10945__597 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__inv_2
X_08376_ net185 net708 net402 net383 net2645 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07327_ net488 _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ _03131_ _03152_ _03914_ _03151_ _03115_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a311o_1
X_10798__450 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__inv_2
XANTENNA__09023__A1 _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__A_N _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06209_ top0.CPU.register.registers\[20\] top0.CPU.register.registers\[52\] top0.CPU.register.registers\[84\]
+ top0.CPU.register.registers\[116\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02866_
+ sky130_fd_sc_hd__mux4_1
X_07189_ net451 _03748_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06503__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08190__C_N net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839__491 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__inv_2
XANTENNA__08782__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_4
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout452 _02635_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_2
XANTENNA__07337__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout496 net499 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
Xfanout485 net486 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06458__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12772_ net767 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11723_ net1415 _01362_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[216\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ net1346 _01293_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[147\]
+ sky130_fd_sc_hd__dfrtp_1
X_11024__676 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__inv_2
XFILLER_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408__60 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__inv_2
X_11585_ net1277 _01224_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08065__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08368__A3 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ net1898 _01845_ net991 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[699\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08773__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09009__B net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ net1829 _01776_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[630\]
+ sky130_fd_sc_hd__dfrtp_1
X_12068_ net1760 _01707_ net991 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[561\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07328__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08525__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591__243 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__inv_2
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08540__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10632__284 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__inv_2
X_06560_ top0.CPU.register.registers\[145\] top0.CPU.register.registers\[177\] top0.CPU.register.registers\[209\]
+ top0.CPU.register.registers\[241\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__mux4_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06491_ _03146_ _03147_ net764 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__mux2_1
X_08230_ net506 net219 net684 net423 net2330 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a32o_1
XANTENNA__10177__Y _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07199__B _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08161_ net205 net617 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07112_ net474 _03054_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__nand2_1
X_08092_ net2833 net436 _04667_ net502 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a22o_1
XANTENNA__05814__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07043_ net743 _03699_ _03693_ _03694_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__o2bb2a_4
Xclkload62 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_16
Xclkload51 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_4
Xclkload40 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_6
Xclkload73 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_132_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05728__A _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload95 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_8
Xclkload84 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__inv_16
XANTENNA__12622__Q net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08994_ top0.CPU.register.registers\[167\] net570 net557 vssd1 vssd1 vccd1 vccd1
+ _04795_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1018_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _04307_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__and3_1
XANTENNA__07662__B _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout478_A _02575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08516__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ net591 _02456_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__nand2_1
X_09615_ net142 _05148_ _04955_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06559__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06827_ _03467_ _03468_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a21oi_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_48_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05976__S1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06758_ top0.CPU.register.registers\[783\] top0.CPU.register.registers\[815\] top0.CPU.register.registers\[847\]
+ top0.CPU.register.registers\[879\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03415_
+ sky130_fd_sc_hd__mux4_1
X_09546_ net774 _05084_ net128 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
X_09477_ top0.MMIO.WBData_i\[10\] net148 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout812_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05709_ top0.CPU.internalMem.state\[2\] top0.CPU.internalMem.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _02366_ sky130_fd_sc_hd__or2_1
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ _03344_ _03345_ net870 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__mux2_1
XANTENNA__06565__Y _03222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08428_ net2853 _04516_ net373 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__mux2_1
XANTENNA__09244__A1 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload1 clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
X_08359_ _04641_ net388 net381 net2793 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a22o_1
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08713__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06058__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10321_ net2226 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10252_ net26 net654 net593 top0.MMIO.WBData_i\[31\] vssd1 vssd1 vccd1 vccd1 _02298_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08755__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08014__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10263__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ net2241 _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09544__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06230__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575__227 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__inv_2
XANTENNA__08507__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_4
Xfanout282 net284 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10616__268 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__inv_2
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09180__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05967__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06916__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ net1398 _01345_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[199\]
+ sky130_fd_sc_hd__dfrtp_1
X_10469__121 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__inv_2
X_12686_ clknet_leaf_92_clk _02321_ net1084 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06408__S net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06392__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09235__A1 top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11637_ net1329 _01276_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[130\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09786__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06049__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ net1260 _01207_ net1079 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[61\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold708 top0.CPU.register.registers\[786\] vssd1 vssd1 vccd1 vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08994__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold719 top0.CPU.register.registers\[640\] vssd1 vssd1 vccd1 vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
X_11499_ clknet_leaf_82_clk _01138_ net1108 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06143__S net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__B top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05982__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05991_ _02644_ _02645_ _02647_ _02646_ net784 net737 vssd1 vssd1 vccd1 vccd1 _02648_
+ sky130_fd_sc_hd__mux4_1
XFILLER_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07730_ _03847_ _04013_ _04383_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09171__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08865__Y _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _04307_ _04317_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__or2_1
XANTENNA__08513__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07721__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06612_ top0.CPU.register.registers\[773\] top0.CPU.register.registers\[805\] top0.CPU.register.registers\[837\]
+ top0.CPU.register.registers\[869\] net934 net900 vssd1 vssd1 vccd1 vccd1 _03269_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06080__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ _04897_ _05010_ _04893_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a21oi_1
X_07592_ _03361_ _03363_ net344 vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09331_ _04979_ _04589_ _04978_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__or3b_1
XFILLER_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_06543_ net246 _02771_ _02791_ _02831_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_36_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06288__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ top0.CPU.internalMem.pcOut\[9\] _04923_ net607 vssd1 vssd1 vccd1 vccd1 _04924_
+ sky130_fd_sc_hd__mux2_1
X_06474_ _03117_ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_134_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09193_ net604 vssd1 vssd1 vccd1 vccd1 top0.chipSelectTFT sky130_fd_sc_hd__inv_2
XANTENNA__08029__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08213_ net2888 net422 _04699_ net501 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
X_08144_ net512 net150 net622 net428 net2329 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a32o_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08985__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05729__Y _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399__51 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__inv_2
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ net3251 net436 _04660_ net500 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a22o_1
X_07026_ _03681_ _03682_ net762 vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
XANTENNA__06053__S net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08201__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__A3 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06212__A1 _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 top0.CPU.register.registers\[26\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08977_ _04665_ net560 _04789_ net262 net3093 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__a32o_1
Xhold24 top0.CPU.register.registers\[5\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A1 top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 top0.CPU.register.registers\[299\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 top0.CPU.register.registers\[464\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07960__X _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07928_ net562 _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or2_1
Xhold57 top0.CPU.register.registers\[806\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 top0.CPU.register.registers\[935\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xhold68 top0.CPU.register.registers\[960\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ net713 net209 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__and2_1
XANTENNA__06071__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05949__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ net955 _05080_ net125 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06279__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08268__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960__612 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__inv_2
XANTENNA__09112__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ clknet_leaf_79_clk _02179_ net1107 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06228__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12471_ net2163 _02110_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[964\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11095__747 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__inv_2
X_11422_ clknet_leaf_68_clk _01070_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08443__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07228__B1 _03882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06126__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08991__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136__788 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__inv_2
X_10304_ net3245 net118 net111 _05671_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
X_10235_ net7 net656 net595 top0.MMIO.WBData_i\[14\] vssd1 vssd1 vccd1 vccd1 _02281_
+ sky130_fd_sc_hd__a22o_1
Xfanout1022 net1024 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
Xfanout1011 net1018 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout1000 net1001 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_2
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_2
Xfanout1044 net1055 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_2
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1033 net1035 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10166_ _02970_ _02979_ net551 vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_89_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ net3371 net665 _05167_ _05568_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a211o_1
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
Xfanout1088 net1132 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_2
Xfanout1077 net1088 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_2
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09153__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06062__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07703__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09303__A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09022__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ clknet_leaf_91_clk _02304_ net1085 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
X_06190_ top0.CPU.register.registers\[277\] top0.CPU.register.registers\[309\] top0.CPU.register.registers\[341\]
+ top0.CPU.register.registers\[373\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02847_
+ sky130_fd_sc_hd__mux4_1
X_10744__396 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06117__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08967__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold516 top0.CPU.register.registers\[367\] vssd1 vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06381__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold505 top0.CPU.register.registers\[452\] vssd1 vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 top0.CPU.register.registers\[477\] vssd1 vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 top0.CPU.register.registers\[126\] vssd1 vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 top0.CPU.register.registers\[363\] vssd1 vssd1 vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
X_08900_ top0.CPU.register.registers\[234\] net573 net559 vssd1 vssd1 vccd1 vccd1
+ _04768_ sky130_fd_sc_hd__o21a_1
X_09880_ _05377_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nor2_1
XANTENNA__08195__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ top0.CPU.decoder.instruction\[11\] _02397_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _04752_ sky130_fd_sc_hd__or3_4
XANTENNA__08589__A top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1205 top0.CPU.intMem_out\[23\] vssd1 vssd1 vccd1 vccd1 net3427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 top0.CPU.intMem_out\[4\] vssd1 vssd1 vccd1 vccd1 net3438 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05974_ top0.CPU.register.registers\[388\] top0.CPU.register.registers\[420\] top0.CPU.register.registers\[452\]
+ top0.CPU.register.registers\[484\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02631_
+ sky130_fd_sc_hd__mux4_1
X_10638__290 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__inv_2
X_08762_ net158 net614 net306 net293 net2565 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__a32o_1
X_07713_ net450 _03975_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__and2_1
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09144__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ net155 net693 net316 net298 net2494 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_127_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09695__B2 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07644_ net488 _04243_ _04300_ _03841_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__a211o_1
XFILLER_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07575_ _02432_ _03712_ _04217_ _04230_ _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__o311a_1
XANTENNA__11920__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06526_ _03181_ _03182_ net871 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
X_09314_ _04962_ _04963_ _04964_ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout510_A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ top0.CPU.internalMem.pcOut\[3\] _04906_ net609 vssd1 vssd1 vccd1 vccd1 _04907_
+ sky130_fd_sc_hd__mux2_1
X_06457_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout608_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06681__A1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ top0.CPU.register.registers\[38\] net565 net553 vssd1 vssd1 vccd1 vccd1 _04848_
+ sky130_fd_sc_hd__o21a_1
X_06388_ top0.CPU.register.registers\[541\] top0.CPU.register.registers\[573\] top0.CPU.register.registers\[605\]
+ top0.CPU.register.registers\[637\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03045_
+ sky130_fd_sc_hd__mux4_1
X_08127_ net3054 _04581_ net430 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07955__X _04592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05867__S0 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08058_ net502 net154 net705 net440 net2290 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a32o_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
X_07009_ _03621_ _03659_ _03661_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout977_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
X_10020_ net589 _03009_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__nor2_1
XANTENNA__08186__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06511__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06292__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ net1663 _01610_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[464\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08489__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06044__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06595__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06747__A _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687__339 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__inv_2
XANTENNA__09438__A1 top0.MMIO.WBData_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12523_ net2215 _02162_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1016\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06672__A1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12454_ net2146 _02093_ net1127 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[947\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08949__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ clknet_leaf_87_clk _01053_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08413__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ net2077 _02024_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07865__X _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07584__Y _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08177__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10218_ net1 top0.wishbone0.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nand2_1
XANTENNA__05826__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ top0.display.delayctr\[24\] net663 _05141_ _05607_ _05610_ vssd1 vssd1 vccd1
+ vccd1 _02233_ sky130_fd_sc_hd__a221o_1
XANTENNA__06283__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09017__B net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06035__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05690_ net778 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07360_ _03558_ _03967_ _03542_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_46_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06311_ net782 _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__and2_1
X_09030_ _04586_ net3235 net352 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__mux2_1
XANTENNA__08652__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07291_ net347 _03923_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or2_1
XFILLER_31_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07860__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06242_ top0.CPU.register.registers\[152\] top0.CPU.register.registers\[184\] top0.CPU.register.registers\[216\]
+ top0.CPU.register.registers\[248\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02899_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08404__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06173_ net581 _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nand2_1
Xhold302 top0.CPU.register.registers\[710\] vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
X_10369__21 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__inv_2
XANTENNA__05849__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold313 top0.CPU.register.registers\[551\] vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 top0.CPU.register.registers\[340\] vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07000__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold335 top0.CPU.register.registers\[212\] vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold357 top0.CPU.register.registers\[447\] vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 top0.CPU.register.registers\[170\] vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ top0.CPU.internalMem.pcOut\[23\] _05416_ vssd1 vssd1 vccd1 vccd1 _05427_
+ sky130_fd_sc_hd__nor2_1
Xhold368 top0.CPU.register.registers\[718\] vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout815 net818 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08168__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold379 top0.CPU.register.registers\[377\] vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_4
XANTENNA__05736__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09863_ top0.CPU.internalMem.pcOut\[18\] _05362_ vssd1 vssd1 vccd1 vccd1 _05363_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout837 net840 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
Xfanout826 net828 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
X_08814_ net198 net675 net325 net287 net2554 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a32o_1
Xhold1013 top0.CPU.register.registers\[140\] vssd1 vssd1 vccd1 vccd1 net3235 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _05297_ _05299_ _05294_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1000_A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 top0.CPU.decoder.instruction\[19\] vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_8
Xhold1024 top0.CPU.register.registers\[988\] vssd1 vssd1 vccd1 vccd1 net3246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1002 top0.CPU.register.registers\[785\] vssd1 vssd1 vccd1 vccd1 net3224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 top0.CPU.register.registers\[510\] vssd1 vssd1 vccd1 vccd1 net3257 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ top0.CPU.register.registers\[368\] net572 _04736_ vssd1 vssd1 vccd1 vccd1
+ _04747_ sky130_fd_sc_hd__o21a_1
Xhold1046 top0.CPU.register.registers\[242\] vssd1 vssd1 vccd1 vccd1 net3268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1057 net94 vssd1 vssd1 vccd1 vccd1 net3279 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__A2 _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 top0.CPU.register.registers\[80\] vssd1 vssd1 vccd1 vccd1 net3290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1079 top0.CPU.register.registers\[166\] vssd1 vssd1 vccd1 vccd1 net3301 sky130_fd_sc_hd__dlygate4sd3_1
X_05957_ net741 _02605_ _02612_ _02613_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__08340__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ net200 net695 net319 net299 net2473 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a32o_1
X_05888_ top0.CPU.register.registers\[259\] top0.CPU.register.registers\[291\] top0.CPU.register.registers\[323\]
+ top0.CPU.register.registers\[355\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02545_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06577__S1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ net482 _04037_ _04117_ net337 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ _04209_ _04211_ _04214_ _04139_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__o31a_1
XANTENNA__06286__B _02942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08891__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06509_ top0.CPU.register.registers\[275\] top0.CPU.register.registers\[307\] top0.CPU.register.registers\[339\]
+ top0.CPU.register.registers\[371\] net939 net906 vssd1 vssd1 vccd1 vccd1 _03166_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_24_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08643__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ _03928_ _04142_ _04144_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__and4_1
X_09228_ top0.CPU.internalMem.pcOut\[15\] top0.CPU.internalMem.pcOut\[14\] top0.CPU.internalMem.pcOut\[13\]
+ top0.CPU.internalMem.pcOut\[31\] vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__or4_1
XANTENNA__07851__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09159_ _04716_ net279 net249 net2804 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a22o_1
XANTENNA__10202__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ net1862 _01809_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[663\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08946__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold891 net82 vssd1 vssd1 vccd1 vccd1 net3113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold880 top0.CPU.register.registers\[251\] vssd1 vssd1 vccd1 vccd1 net3102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ top0.CPU.internalMem.pcOut\[27\] _05467_ top0.CPU.internalMem.pcOut\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05917__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09108__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11954_ net1646 _01593_ net1097 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06342__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11885_ net1577 _01524_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[378\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06893__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_43_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08095__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08634__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__B _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ net2198 _02145_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[999\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06740__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ net2129 _02076_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[930\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12368_ net2060 _02007_ net1083 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[861\]
+ sky130_fd_sc_hd__dfrtp_1
X_11151__803 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__inv_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12299_ net1991 _01938_ net1072 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06151__S net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ _03513_ _03514_ _03515_ _03516_ net761 net864 vssd1 vssd1 vccd1 vccd1 _03517_
+ sky130_fd_sc_hd__mux4_1
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06256__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05811_ top0.CPU.register.registers\[403\] top0.CPU.register.registers\[435\] top0.CPU.register.registers\[467\]
+ top0.CPU.register.registers\[499\] net856 net821 vssd1 vssd1 vccd1 vccd1 _02468_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08570__A1 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ top0.CPU.register.registers\[652\] top0.CPU.register.registers\[684\] top0.CPU.register.registers\[716\]
+ top0.CPU.register.registers\[748\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03448_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_124_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05742_ net575 _02394_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__and2_4
X_08530_ net206 net3074 net362 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__mux2_1
XANTENNA__08322__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08461_ _04678_ net387 net369 net2694 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07412_ _04045_ _04046_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08873__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ _04657_ net388 net377 net2703 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XANTENNA__08086__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07343_ _03998_ _03999_ net347 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__mux2_1
Xteam_07_1136 vssd1 vssd1 vccd1 vccd1 team_07_1136/HI gpio_oeb[5] sky130_fd_sc_hd__conb_1
XANTENNA__08107__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ net442 _03928_ _03929_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__o211a_1
XANTENNA__06636__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1158 vssd1 vssd1 vccd1 vccd1 team_07_1158/HI gpio_out[24] sky130_fd_sc_hd__conb_1
XANTENNA__06731__S1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06225_ _02880_ _02881_ net731 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
Xteam_07_1147 vssd1 vssd1 vccd1 vccd1 team_07_1147/HI gpio_out[13] sky130_fd_sc_hd__conb_1
Xteam_07_1169 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] team_07_1169/LO sky130_fd_sc_hd__conb_1
X_09013_ top0.CPU.register.registers\[153\] net564 vssd1 vssd1 vccd1 vccd1 _04800_
+ sky130_fd_sc_hd__or2_1
Xhold110 top0.CPU.register.registers\[255\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 top0.CPU.register.registers\[812\] vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 top0.CPU.register.registers\[991\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06156_ net907 _02474_ _02472_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a21o_1
X_10800__452 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__inv_2
Xhold132 top0.CPU.register.registers\[323\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 top0.CPU.register.registers\[293\] vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
X_06087_ top0.CPU.register.registers\[269\] top0.CPU.register.registers\[301\] top0.CPU.register.registers\[333\]
+ top0.CPU.register.registers\[365\] net850 net815 vssd1 vssd1 vccd1 vccd1 _02744_
+ sky130_fd_sc_hd__mux4_1
Xhold165 top0.CPU.register.registers\[808\] vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 top0.CPU.register.registers\[689\] vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_2
Xhold187 top0.CPU.register.registers\[1002\] vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 top0.CPU.register.registers\[1007\] vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _04854_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_2
X_09915_ top0.CPU.internalMem.pcOut\[22\] _05409_ vssd1 vssd1 vccd1 vccd1 _05411_
+ sky130_fd_sc_hd__xor2_1
Xfanout601 _04859_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_2
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_2
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout634 _02395_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_4
X_09846_ top0.CPU.internalMem.pcOut\[15\] top0.CPU.internalMem.pcOut\[16\] _05325_
+ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and3_1
XFILLER_98_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout645 net649 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_2
Xfanout667 _04855_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08010__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 _04687_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08561__A1 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09777_ _03989_ net234 net229 net631 vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout842_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ top0.CPU.register.registers\[922\] top0.CPU.register.registers\[954\] top0.CPU.register.registers\[986\]
+ top0.CPU.register.registers\[1018\] net910 net876 vssd1 vssd1 vccd1 vccd1 _03646_
+ sky130_fd_sc_hd__mux4_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08728_ net155 net3116 net358 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ net155 net705 net316 net302 net2378 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08716__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ net1362 _01309_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09401__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06627__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06236__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09120__B net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09577__A0 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ net1914 _01861_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[715\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06760__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07588__C1 _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543__195 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__inv_2
XANTENNA__08451__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net1845 _01792_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06486__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12084_ net1776 _01723_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06238__S0 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08304__A1 _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06000__A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ net1629 _01576_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[430\]
+ sky130_fd_sc_hd__dfrtp_1
X_11868_ net1560 _01507_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[361\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08607__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11799_ net1491 _01438_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06713__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05985__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06010_ _02666_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__inv_2
XANTENNA__10178__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ net720 net509 net184 net547 net2409 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a32o_1
XFILLER_87_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09700_ _05199_ _05204_ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__o21ai_1
X_06912_ _03490_ net526 _03568_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a21o_1
X_07892_ top0.CPU.internalMem.pcOut\[21\] net640 net635 _04538_ vssd1 vssd1 vccd1
+ vccd1 _04539_ sky130_fd_sc_hd__o211a_2
XFILLER_110_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06843_ top0.CPU.register.registers\[11\] top0.CPU.register.registers\[43\] top0.CPU.register.registers\[75\]
+ top0.CPU.register.registers\[107\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03500_
+ sky130_fd_sc_hd__mux4_1
X_09631_ net142 _05160_ _04955_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05733__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ net652 net238 vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_4
X_06774_ top0.CPU.register.registers\[782\] top0.CPU.register.registers\[814\] top0.CPU.register.registers\[846\]
+ top0.CPU.register.registers\[878\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03431_
+ sky130_fd_sc_hd__mux4_1
X_05725_ _02378_ _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__nor2_1
X_08513_ net173 net683 net399 net367 net2675 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a32o_1
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _02355_ net139 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout256_A _04809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08444_ net2801 _04600_ net375 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__mux2_1
X_11320__972 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__inv_2
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486__138 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__inv_2
X_08375_ net186 net706 net398 net383 net2437 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a32o_1
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06056__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07326_ _03979_ _03982_ net345 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__mux2_1
X_07257_ _03246_ _03576_ _03132_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10527__179 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__inv_2
XANTENNA__09023__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06208_ top0.CPU.register.registers\[148\] top0.CPU.register.registers\[180\] top0.CPU.register.registers\[212\]
+ top0.CPU.register.registers\[244\] net833 net798 vssd1 vssd1 vccd1 vccd1 _02865_
+ sky130_fd_sc_hd__mux4_1
X_07188_ net450 _03806_ _03826_ _03830_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a2111o_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06139_ _02794_ _02795_ net726 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
Xfanout431 net432 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
Xfanout420 _04706_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 _03752_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
Xfanout453 _02635_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_2
Xfanout464 net466 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07337__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 _02598_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_2
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _05318_ _05323_ _05330_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__or3_1
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
Xfanout486 _02555_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_4
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06640__S0 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771_ net61 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11434__Q top0.CPU.intMem_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08446__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11722_ net1414 _01361_ net965 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[215\]
+ sky130_fd_sc_hd__dfrtp_1
X_11653_ net1345 _01292_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_120_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06474__B _03130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05808__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11584_ net1276 _01223_ net1030 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08470__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423__75 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09014__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ net1897 _01844_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[698\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ net1828 _01775_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[629\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_97_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12067_ net1759 _01706_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[560\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263__915 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__inv_2
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08828__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304__956 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__inv_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06490_ top0.CPU.register.registers\[21\] top0.CPU.register.registers\[53\] top0.CPU.register.registers\[85\]
+ top0.CPU.register.registers\[117\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03147_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_103_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ net3316 net425 _04680_ net491 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a22o_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09253__A2 top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08056__A3 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07111_ _03764_ _03767_ net347 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08091_ net221 net693 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and2_1
XANTENNA__08461__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07042_ _03695_ _03696_ _03697_ _03698_ net730 top0.CPU.control.rs2\[3\] vssd1 vssd1
+ vccd1 vccd1 _03699_ sky130_fd_sc_hd__mux4_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload52 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__inv_16
XANTENNA__06604__S net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload41 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__clkinv_8
Xclkload30 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_12
Xclkload74 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_132_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload63 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__inv_16
Xclkload96 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_12
XANTENNA__11945__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload85 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_16
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871__523 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__inv_2
X_08993_ net218 net695 net277 net260 net2596 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__B _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ net722 net514 net195 net547 net2349 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a32o_1
XANTENNA__05744__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _03939_ _04474_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__nor2_1
XFILLER_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10912__564 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__inv_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09614_ _02665_ _05007_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__or2_1
X_06826_ _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout373_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_48_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06757_ _03412_ _03413_ net762 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
X_09545_ net781 _05059_ net128 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XANTENNA__08819__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_129_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09476_ net130 net133 _05056_ net598 net3336 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__o32a_1
X_05708_ top0.CPU.internalMem.state\[2\] top0.CPU.internalMem.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _02365_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ top0.CPU.register.registers\[896\] top0.CPU.register.registers\[928\] top0.CPU.register.registers\[960\]
+ top0.CPU.register.registers\[992\] net921 net887 vssd1 vssd1 vccd1 vccd1 _03345_
+ sky130_fd_sc_hd__mux4_1
X_11047__699 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ net2871 _04510_ net373 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A3 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ _04640_ net392 net381 net3034 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a22o_1
Xclkload2 clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
X_08289_ net2889 net212 net415 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
X_07309_ net342 _03943_ _03944_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__a31o_1
XANTENNA__07255__A1 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06514__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ net2223 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09643__B1_N _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ net25 net656 net595 top0.MMIO.WBData_i\[30\] vssd1 vssd1 vccd1 vccd1 _02297_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09952__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ net663 net602 _05636_ top0.display.delayctr\[31\] vssd1 vssd1 vccd1 vccd1
+ _05637_ sky130_fd_sc_hd__o22a_1
Xfanout250 _04842_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_4
XFILLER_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_4
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout272 net281 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
Xfanout294 _04746_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09180__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06613__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ net1397 _01344_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[198\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08286__A3 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12685_ clknet_leaf_91_clk _02320_ net1084 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08691__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A3 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ net1328 _01275_ net961 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[129\]
+ sky130_fd_sc_hd__dfrtp_1
X_11567_ net1259 _01206_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07790__A1_N net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06424__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold709 top0.CPU.register.registers\[886\] vssd1 vssd1 vccd1 vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ clknet_leaf_82_clk net3305 net1108 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10855__507 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__inv_2
XFILLER_124_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05990_ top0.CPU.register.registers\[5\] top0.CPU.register.registers\[37\] top0.CPU.register.registers\[69\]
+ top0.CPU.register.registers\[101\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02647_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06852__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12119_ net1811 _01758_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[612\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ net343 _03941_ _04308_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a31o_1
XFILLER_38_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06611_ _03266_ _03267_ net761 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__mux2_1
X_10749__401 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__inv_2
XANTENNA__06080__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07591_ net342 _04233_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a21o_1
XFILLER_53_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10353__5 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09330_ _04604_ _04608_ _04612_ _04616_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__or4_1
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06542_ net246 _02771_ _02791_ net543 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_36_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08277__A3 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ top0.CPU.intMemAddr\[9\] _04597_ net770 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06288__A2 _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06395__A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08682__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06473_ net859 _03122_ _03128_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a21bo_1
X_08212_ net204 net682 vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__and2_1
X_09192_ top0.display.state\[0\] net666 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__and2b_1
XANTENNA__07003__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08143_ net946 _02399_ net624 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__nand3_4
XANTENNA_fanout121_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10241__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_A _04603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05739__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__A2 _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ net207 net693 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and2_1
X_07025_ top0.CPU.register.registers\[31\] top0.CPU.register.registers\[63\] top0.CPU.register.registers\[95\]
+ top0.CPU.register.registers\[127\] net936 net903 vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12633__Q top0.MMIO.WBData_i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05799__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold14 top0.CPU.register.registers\[12\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06843__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ top0.CPU.register.registers\[179\] net575 vssd1 vssd1 vccd1 vccd1 _04789_
+ sky130_fd_sc_hd__or2_1
Xhold47 top0.CPU.register.registers\[844\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold25 top0.CPU.register.registers\[11\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold36 top0.CPU.register.registers\[419\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 top0.CPU.register.registers\[44\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ _04354_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__and3_1
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05971__A1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 top0.CPU.register.registers\[291\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ top0.CPU.internalMem.pcOut\[26\] net638 net633 _04509_ vssd1 vssd1 vccd1
+ vccd1 _04510_ sky130_fd_sc_hd__o211a_4
XFILLER_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06071__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06809_ _03447_ net527 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__xnor2_1
X_07789_ _02750_ _03482_ net444 _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout922_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09528_ top0.CPU.Op\[6\] _05078_ net126 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_14_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ top0.MMIO.WBData_i\[23\] net146 net135 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08724__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ net2162 _02109_ net988 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[963\]
+ sky130_fd_sc_hd__dfrtp_1
X_11421_ clknet_leaf_68_clk _01069_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07228__B2 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10303_ _04938_ _05624_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__or2_1
XANTENNA__06244__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10234_ net6 net653 net592 net3401 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__o22a_1
Xfanout1012 net1018 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
XFILLER_79_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06834__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 net1004 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_2
X_10165_ net3374 net663 net602 _05623_ _05621_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a221o_1
XANTENNA__07400__B2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1045 net1047 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 net1132 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__clkbuf_2
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1089 net1092 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10096_ _05566_ _05567_ net601 vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
Xfanout1067 net1070 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08695__A _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06062__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__A2 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09303__B _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08259__A3 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08664__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12668_ clknet_leaf_91_clk _02303_ net1084 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XFILLER_128_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11619_ net1311 _01258_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08416__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12599_ clknet_leaf_89_clk _02234_ net1087 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06662__B _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold506 top0.CPU.register.registers\[605\] vssd1 vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 top0.CPU.register.registers\[311\] vssd1 vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 top0.CPU.register.registers\[632\] vssd1 vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 top0.CPU.register.registers\[568\] vssd1 vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08195__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07493__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269__921 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__inv_2
X_08830_ net155 net671 net314 net286 net2520 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_111_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1206 top0.display.delayctr\[21\] vssd1 vssd1 vccd1 vccd1 net3428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold1217 top0.display.delayctr\[3\] vssd1 vssd1 vccd1 vccd1 net3439 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ net162 net615 net309 net294 net2304 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__a32o_1
X_05973_ top0.CPU.register.registers\[4\] top0.CPU.register.registers\[36\] top0.CPU.register.registers\[68\]
+ top0.CPU.register.registers\[100\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02630_
+ sky130_fd_sc_hd__mux4_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12325__RESET_B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _03657_ _04367_ _03663_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07155__B1 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ net158 net690 net309 net297 net2432 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a32o_1
X_07643_ net483 _04237_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout169_A _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05741__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06396__Y _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983__635 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__inv_2
XFILLER_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07574_ _03710_ _03737_ _04216_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__or3_1
X_09313_ top0.display.delayctr\[4\] top0.display.delayctr\[7\] top0.display.delayctr\[16\]
+ top0.display.delayctr\[17\] vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__or4_1
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_A _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06525_ top0.CPU.register.registers\[914\] top0.CPU.register.registers\[946\] top0.CPU.register.registers\[978\]
+ top0.CPU.register.registers\[1010\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03182_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08655__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
X_09244_ top0.CPU.intMemAddr\[3\] _04619_ net769 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__mux2_1
X_06456_ _03096_ net536 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ net175 net669 net276 net249 net2260 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06387_ top0.CPU.register.registers\[669\] top0.CPU.register.registers\[701\] top0.CPU.register.registers\[733\]
+ top0.CPU.register.registers\[765\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03044_
+ sky130_fd_sc_hd__mux4_1
X_08126_ net3106 _04576_ net432 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout503_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05867__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ net493 _04630_ net701 net437 net2350 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a32o_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
X_07008_ _03660_ _03662_ _03638_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__o21bai_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_10918__570 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__inv_2
XFILLER_0_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08186__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06816__S0 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__A0 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ net150 net699 net280 net262 net2261 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06292__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ net1662 _01609_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08011__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06044__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07697__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08894__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062__714 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__inv_2
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08646__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_51_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07859__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ net2214 _02161_ net984 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1015\]
+ sky130_fd_sc_hd__dfrtp_1
X_11103__755 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__inv_2
XANTENNA__08962__B net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ net2145 _02092_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[946\]
+ sky130_fd_sc_hd__dfrtp_1
X_12384_ net2076 _02023_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[877\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09071__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ clknet_leaf_87_clk _01052_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09610__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08413__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07621__A1 _02578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07621__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ net1 top0.wishbone0.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__and2_1
XFILLER_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08202__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07924__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _05608_ _05609_ net600 vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06283__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967__619 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__inv_2
X_10079_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__nand2_1
XANTENNA__07137__A0 _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670__322 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__inv_2
XANTENNA__06035__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09033__B net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711__363 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08637__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
X_07290_ net490 _03719_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or2_1
X_06310_ top0.CPU.register.registers\[924\] top0.CPU.register.registers\[956\] top0.CPU.register.registers\[988\]
+ top0.CPU.register.registers\[1020\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02967_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08652__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06241_ net780 _02893_ _02896_ _02897_ net771 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__o221a_1
XANTENNA__07488__B _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06172_ net743 _02828_ _02820_ _02821_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__09062__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__X _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 top0.CPU.register.registers\[339\] vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05849__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold314 top0.CPU.register.registers\[555\] vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 top0.CPU.register.registers\[87\] vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09048__X _04809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold347 top0.CPU.intMemAddr\[2\] vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 top0.CPU.intMemAddr\[31\] vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ top0.CPU.internalMem.pcOut\[23\] _05416_ vssd1 vssd1 vccd1 vccd1 _05426_
+ sky130_fd_sc_hd__and2_1
Xhold369 top0.CPU.register.registers\[572\] vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 top0.CPU.register.registers\[686\] vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout816 net818 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08168__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06060__A2_N net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_2
XFILLER_131_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 net854 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09862_ _02495_ _04552_ net587 vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__mux2_1
X_10384__36 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__inv_2
Xfanout838 net840 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_2
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_4
XFILLER_112_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09793_ _05261_ _05274_ _05295_ _05298_ _05287_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a32o_1
Xhold1003 top0.CPU.register.registers\[173\] vssd1 vssd1 vccd1 vccd1 net3225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 top0.CPU.register.registers\[48\] vssd1 vssd1 vccd1 vccd1 net3236 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net200 net673 net319 net287 net2425 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_51_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1036 top0.CPU.register.registers\[45\] vssd1 vssd1 vccd1 vccd1 net3258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 top0.CPU.register.registers\[267\] vssd1 vssd1 vccd1 vccd1 net3280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1025 net75 vssd1 vssd1 vccd1 vccd1 net3247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 top0.CPU.register.registers\[154\] vssd1 vssd1 vccd1 vccd1 net3269 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _04685_ net307 net293 net2657 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22o_1
X_05956_ net735 _02608_ net772 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05752__A _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1069 top0.display.delayctr\[15\] vssd1 vssd1 vccd1 vccd1 net3291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout453_A _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _04666_ net308 net297 net2689 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a22o_1
X_05887_ net736 _02539_ _02542_ _02543_ net741 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a221o_2
XFILLER_81_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07626_ net462 _04254_ _04282_ net476 vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__o211a_1
XANTENNA__05785__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08628__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07557_ _04212_ _04213_ _04143_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__a21oi_1
X_06508_ net867 _03160_ _03163_ _03164_ net861 vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_33_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout718_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07679__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07488_ _02869_ _03129_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__xnor2_1
X_09227_ _04885_ _04886_ _04887_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__or4_1
X_06439_ _02888_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__xnor2_1
X_09158_ _04715_ net273 net248 net2740 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__a22o_1
X_08109_ net3132 _04481_ net431 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08800__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ net160 net615 net270 net255 net2263 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__a32o_1
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold870 top0.CPU.register.registers\[532\] vssd1 vssd1 vccd1 vccd1 net3092 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 top0.CPU.register.registers\[85\] vssd1 vssd1 vccd1 vccd1 net3103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 top0.CPU.register.registers\[269\] vssd1 vssd1 vccd1 vccd1 net3114 sky130_fd_sc_hd__dlygate4sd3_1
X_10654__306 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__inv_2
XFILLER_77_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08022__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__Q top0.CPU.intMem_out\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ top0.CPU.internalMem.pcOut\[28\] top0.CPU.internalMem.pcOut\[27\] _05467_
+ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and3_1
XFILLER_49_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06590__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08867__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ net1645 _01592_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06342__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08331__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11884_ net1576 _01523_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[377\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08619__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08095__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548__200 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__inv_2
XANTENNA__07842__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12505_ net2197 _02144_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[998\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12436_ net2128 _02075_ net961 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[929\]
+ sky130_fd_sc_hd__dfrtp_1
X_11190__842 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__inv_2
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12367_ net2059 _02006_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[860\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12298_ net1990 _01937_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[791\]
+ sky130_fd_sc_hd__dfrtp_1
X_11231__883 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__inv_2
XANTENNA__06256__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05810_ top0.CPU.register.registers\[19\] top0.CPU.register.registers\[51\] top0.CPU.register.registers\[83\]
+ top0.CPU.register.registers\[115\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02467_
+ sky130_fd_sc_hd__mux4_1
X_06790_ _02769_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_124_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05741_ _02394_ net634 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__nand2b_2
XFILLER_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ _04677_ net385 net369 net2671 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a22o_1
X_07411_ _04067_ _04055_ _04058_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__and3b_1
X_08391_ _04656_ net392 net377 net2566 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_15_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
X_07342_ net537 net536 net523 net522 net474 net457 vssd1 vssd1 vccd1 vccd1 _03999_
+ sky130_fd_sc_hd__mux4_1
X_10429__81 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__inv_2
XANTENNA__09283__B1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08086__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08625__A3 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ _02457_ _03092_ net341 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a21o_1
Xteam_07_1148 vssd1 vssd1 vccd1 vccd1 team_07_1148/HI gpio_out[14] sky130_fd_sc_hd__conb_1
Xteam_07_1159 vssd1 vssd1 vccd1 vccd1 team_07_1159/HI gpio_out[25] sky130_fd_sc_hd__conb_1
XFILLER_136_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ net209 net3269 net349 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
X_06224_ top0.CPU.register.registers\[22\] top0.CPU.register.registers\[54\] top0.CPU.register.registers\[86\]
+ top0.CPU.register.registers\[118\] net838 net803 vssd1 vssd1 vccd1 vccd1 _02881_
+ sky130_fd_sc_hd__mux4_1
Xteam_07_1137 vssd1 vssd1 vccd1 vccd1 team_07_1137/HI gpio_out[0] sky130_fd_sc_hd__conb_1
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08389__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 top0.CPU.register.registers\[971\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
X_06155_ _02810_ _02811_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__and2_1
Xhold133 top0.CPU.register.registers\[682\] vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 top0.CPU.register.registers\[876\] vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 top0.CPU.register.registers\[1003\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 top0.CPU.register.registers\[839\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold155 top0.CPU.register.registers\[938\] vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
X_06086_ top0.CPU.register.registers\[397\] top0.CPU.register.registers\[429\] top0.CPU.register.registers\[461\]
+ top0.CPU.register.registers\[493\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02743_
+ sky130_fd_sc_hd__mux4_1
Xhold166 top0.CPU.register.registers\[97\] vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 top0.CPU.register.registers\[800\] vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout624 _04670_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_4
Xfanout613 _04797_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_8
Xhold188 top0.CPU.register.registers\[336\] vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ top0.CPU.internalMem.pcOut\[22\] _05409_ vssd1 vssd1 vccd1 vccd1 _05410_
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1110_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_4
Xhold199 top0.CPU.register.registers\[481\] vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout657 _05645_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09653__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_4
X_09845_ _05342_ _05344_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__o21a_1
XANTENNA__07962__A _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net649 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08010__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989__641 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__inv_2
XANTENNA_fanout570_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net681 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_4
Xfanout668 net670 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
X_09776_ net647 _05281_ _05282_ _05110_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a31o_1
XFILLER_74_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06988_ top0.CPU.register.registers\[794\] top0.CPU.register.registers\[826\] top0.CPU.register.registers\[858\]
+ top0.CPU.register.registers\[890\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03645_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_29_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05939_ _02587_ _02595_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ net158 net3213 net357 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__mux2_1
X_08658_ net158 net701 net306 net301 net2433 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a32o_1
XFILLER_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07609_ net486 _04009_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ top0.CPU.decoder.instruction\[11\] _02397_ vssd1 vssd1 vccd1 vccd1 _04734_
+ sky130_fd_sc_hd__nor2_4
XANTENNA__06584__Y _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07824__B2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09026__A0 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174__826 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__inv_2
X_12221_ net1913 _01860_ net1024 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[714\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12152_ net1844 _01791_ net1029 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06486__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215__867 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12083_ net1775 _01722_ net1065 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[576\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06238__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08552__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068__720 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__inv_2
X_11936_ net1628 _01575_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[429\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_45_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11109__761 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__inv_2
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ net1559 _01506_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[360\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10782__434 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__inv_2
X_11798_ net1490 _01437_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10823__475 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__inv_2
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09568__A1 _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12419_ net2111 _02058_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10178__A2 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06162__S net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ top0.CPU.internalMem.pcOut\[10\] net641 net636 _04595_ vssd1 vssd1 vccd1
+ vccd1 _04596_ sky130_fd_sc_hd__o211a_4
XANTENNA__06251__A0 _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05854__X _02511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06911_ _03507_ _03518_ _03490_ net526 vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_4_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07891_ top0.CPU.intMem_out\[21\] net630 _04537_ net643 vssd1 vssd1 vccd1 vccd1 _04538_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__05988__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06842_ top0.CPU.register.registers\[139\] top0.CPU.register.registers\[171\] top0.CPU.register.registers\[203\]
+ top0.CPU.register.registers\[235\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03499_
+ sky130_fd_sc_hd__mux4_1
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09630_ _02532_ _05150_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__or2_1
XANTENNA__05733__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ net238 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__inv_2
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06773_ top0.CPU.register.registers\[910\] top0.CPU.register.registers\[942\] top0.CPU.register.registers\[974\]
+ top0.CPU.register.registers\[1006\] net921 net886 vssd1 vssd1 vccd1 vccd1 _03430_
+ sky130_fd_sc_hd__mux4_1
X_05724_ top0.CPU.Op\[4\] top0.CPU.Op\[5\] top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1
+ _02381_ sky130_fd_sc_hd__nand3b_2
X_08512_ net175 net683 net390 net367 net2477 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a32o_1
X_09492_ _02356_ net139 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__nor2_1
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout249_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ net3049 net185 net375 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__mux2_1
XFILLER_51_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08374_ net191 net710 net407 net384 net2496 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_63_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07325_ _03980_ _03981_ net458 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__mux2_1
XFILLER_32_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07957__A _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06165__S0 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ _03667_ net344 _03887_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout1060_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12592__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06207_ top0.CPU.register.registers\[404\] top0.CPU.register.registers\[436\] top0.CPU.register.registers\[468\]
+ top0.CPU.register.registers\[500\] net833 net798 vssd1 vssd1 vccd1 vccd1 _02864_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05912__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ _03834_ _03839_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06072__S net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06138_ top0.CPU.register.registers\[529\] top0.CPU.register.registers\[561\] top0.CPU.register.registers\[593\]
+ top0.CPU.register.registers\[625\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02795_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout785_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06069_ top0.CPU.register.registers\[138\] top0.CPU.register.registers\[170\] top0.CPU.register.registers\[202\]
+ top0.CPU.register.registers\[234\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02726_
+ sky130_fd_sc_hd__mux4_1
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08782__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout432 _04669_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
Xfanout421 _04689_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
Xfanout410 net412 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout952_A top0.CPU.decoder.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout443 _03751_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
Xfanout454 _02635_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09731__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ _05318_ _05323_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
Xfanout487 net488 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__A3 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ top0.CPU.internalMem.pcOut\[9\] _05254_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06640__S1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08298__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ net767 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11403__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766__418 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__inv_2
XANTENNA__05940__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08727__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11721_ net1413 _01360_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06247__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11652_ net1344 _01291_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[145\]
+ sky130_fd_sc_hd__dfrtp_1
X_10510__162 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__inv_2
XANTENNA__11450__Q top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807__459 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__inv_2
XANTENNA__09798__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11583_ net1275 _01222_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12773__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08970__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07273__A2 _03092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05903__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07078__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12204_ net1896 _01843_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[697\]
+ sky130_fd_sc_hd__dfrtp_1
X_12135_ net1827 _01774_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[628\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08773__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ net1758 _01705_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[559\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08525__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08210__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08289__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08828__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343__995 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__inv_2
XANTENNA__08864__C _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net1611 _01558_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[412\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08880__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07110_ _03765_ _03766_ net465 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__mux2_1
X_08090_ net513 net197 net697 net434 net2300 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__a32o_1
Xclkload20 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_8
X_07041_ top0.CPU.register.registers\[287\] top0.CPU.register.registers\[319\] top0.CPU.register.registers\[351\]
+ top0.CPU.register.registers\[383\] net852 net817 vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__mux4_1
Xclkload53 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_6
Xclkload42 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_2
Xclkload31 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinv_8
Xclkload75 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__clkinv_16
Xclkload64 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_8
Xclkload86 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__inv_4
Xclkload97 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_8
XANTENNA__07421__C1 _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ net180 net696 net277 net260 net2798 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__a32o_1
X_07943_ net634 _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__and2_1
XANTENNA__05744__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07874_ net2900 net549 net501 _04523_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
XANTENNA__08516__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06825_ net860 _03473_ _03477_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453__105 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__inv_2
X_09613_ net3355 net604 net658 net3359 _05147_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__a221o_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout366_A _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06756_ top0.CPU.register.registers\[527\] top0.CPU.register.registers\[559\] top0.CPU.register.registers\[591\]
+ top0.CPU.register.registers\[623\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03413_
+ sky130_fd_sc_hd__mux4_1
X_09544_ net787 _05074_ net127 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XANTENNA__08819__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09475_ top0.MMIO.WBData_i\[31\] net145 net135 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__o21a_1
X_05707_ top0.CPU.internalMem.state\[1\] top0.CPU.internalMem.state\[2\] top0.CPU.internalMem.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09232__A top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05760__A top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout533_A _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06687_ top0.CPU.register.registers\[768\] top0.CPU.register.registers\[800\] top0.CPU.register.registers\[832\]
+ top0.CPU.register.registers\[864\] net921 net887 vssd1 vssd1 vccd1 vccd1 _03344_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_61_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06386__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ net3217 net210 net373 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__mux2_1
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06862__Y _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_6
XANTENNA__06138__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ _04639_ net397 net382 net2789 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a22o_1
X_08288_ net2862 net151 net416 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
X_07308_ _02635_ _03956_ _03961_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__o211ai_2
X_07239_ _03839_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__and2b_1
X_10250_ net23 net653 net592 net3425 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__o22a_1
XANTENNA__07974__X _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ top0.display.delayctr\[30\] net663 _05630_ vssd1 vssd1 vccd1 vccd1 _05636_
+ sky130_fd_sc_hd__nor3_1
XANTENNA__06310__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11286__938 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__inv_2
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08507__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 _04783_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09704__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_4
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
Xfanout284 _04753_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_8
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_4
X_11030__682 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__inv_2
XFILLER_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09180__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08030__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06613__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11327__979 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__inv_2
X_11704_ net1396 _01343_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06377__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12684_ clknet_leaf_91_clk _02319_ net1085 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06129__S0 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11635_ net1327 _01274_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07246__A2 _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11566_ net1258 _01205_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ clknet_leaf_91_clk _01136_ net1085 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894__546 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__inv_2
XFILLER_108_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08746__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06301__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935__587 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__inv_2
XANTENNA__06852__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ net1810 _01757_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[611\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ net1741 _01688_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[542\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11396__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06610_ top0.CPU.register.registers\[517\] top0.CPU.register.registers\[549\] top0.CPU.register.registers\[581\]
+ top0.CPU.register.registers\[613\] net934 net900 vssd1 vssd1 vccd1 vccd1 _03267_
+ sky130_fd_sc_hd__mux4_1
X_07590_ _04241_ _04246_ _04236_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10788__440 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__inv_2
XFILLER_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06541_ _03196_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06368__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ top0.CPU.internalMem.pcOut\[8\] _04921_ net608 vssd1 vssd1 vccd1 vccd1 _04922_
+ sky130_fd_sc_hd__mux2_1
X_06472_ net858 _03122_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a21boi_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10829__481 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__inv_2
XANTENNA__05730__D net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ net3136 net422 _04698_ net500 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
X_09191_ top0.display.state\[2\] top0.display.state\[1\] vssd1 vssd1 vccd1 vccd1 _04855_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_134_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08142_ net951 _02389_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or2_1
XANTENNA__08434__A1 _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08985__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload120 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__05739__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07300__A _02578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ net2953 net433 _04659_ net493 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a22o_1
X_07024_ top0.CPU.register.registers\[159\] top0.CPU.register.registers\[191\] top0.CPU.register.registers\[223\]
+ top0.CPU.register.registers\[255\] net937 net903 vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_58_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08737__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _04664_ net554 _04788_ net259 net3222 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__a32o_1
Xhold15 top0.CPU.register.registers\[9\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 top0.CPU.register.registers\[13\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07926_ net719 net505 net199 net547 net2345 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_71_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014__666 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__inv_2
Xhold37 top0.CPU.register.registers\[865\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold59 top0.CPU.register.registers\[292\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 top0.CPU.register.registers\[672\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07857_ top0.CPU.intMem_out\[26\] net627 _04508_ net642 vssd1 vssd1 vccd1 vccd1 _04509_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08370__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__A1 _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06808_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__inv_2
X_07788_ _02750_ _03482_ net340 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a21o_1
X_09527_ top0.CPU.Op\[5\] _05087_ net127 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06739_ top0.CPU.register.registers\[134\] top0.CPU.register.registers\[166\] top0.CPU.register.registers\[198\]
+ top0.CPU.register.registers\[230\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03396_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06359__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07969__X _04603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ net132 net134 _05047_ _04948_ net3420 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__o32a_1
XFILLER_52_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08409_ net185 net696 net402 net379 net2355 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a32o_1
X_09389_ _02409_ _04988_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11420_ clknet_leaf_68_clk _01068_ net1101 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10581__233 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__inv_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07210__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ net3089 net118 net111 _05670_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10622__274 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__inv_2
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08189__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ net5 net653 net592 net3429 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__o22a_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07936__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1013 net1018 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
X_10164_ _04970_ _05604_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__o21ai_1
Xfanout1002 net1004 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
Xfanout1024 net1056 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
XANTENNA__06834__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10095_ top0.display.delayctr\[13\] _05562_ top0.display.delayctr\[14\] vssd1 vssd1
+ vccd1 vccd1 _05567_ sky130_fd_sc_hd__o21ai_1
Xfanout1079 net1087 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10299__A1 _02942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1057 net1059 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_4
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06598__S0 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09153__A2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08900__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06911__B2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07879__X _04528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ clknet_leaf_92_clk _02302_ net1082 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
X_11618_ net1310 _01257_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12598_ clknet_leaf_88_clk _02233_ net1078 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08967__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ net1241 _01188_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[42\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold507 top0.CPU.register.registers\[908\] vssd1 vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06522__S0 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold518 top0.CPU.register.registers\[53\] vssd1 vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 top0.CPU.register.registers\[345\] vssd1 vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06170__S net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 top0.MMIO.WBData_i\[12\] vssd1 vssd1 vccd1 vccd1 net3429 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05938__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05972_ top0.CPU.register.registers\[132\] top0.CPU.register.registers\[164\] top0.CPU.register.registers\[196\]
+ top0.CPU.register.registers\[228\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02629_
+ sky130_fd_sc_hd__mux4_1
Xhold1218 top0.display.delayctr\[29\] vssd1 vssd1 vccd1 vccd1 net3440 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08760_ net165 net616 net311 net293 net2733 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__a32o_1
X_07711_ _03657_ _03663_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__or3_1
XFILLER_66_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08691_ net162 net691 net309 net297 net2341 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a32o_1
XANTENNA__07155__A1 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09144__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07642_ _02769_ _03463_ net340 vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__a21o_1
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08352__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09312_ top0.display.delayctr\[28\] top0.display.delayctr\[29\] top0.display.delayctr\[30\]
+ top0.display.delayctr\[31\] vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__or4_1
X_07573_ _04050_ _04218_ _04222_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__o211a_1
XANTENNA__08104__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06524_ top0.CPU.register.registers\[786\] top0.CPU.register.registers\[818\] top0.CPU.register.registers\[850\]
+ top0.CPU.register.registers\[882\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03181_
+ sky130_fd_sc_hd__mux4_1
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ top0.CPU.internalMem.pcOut\[1\] _04904_ net611 vssd1 vssd1 vccd1 vccd1 _04905_
+ sky130_fd_sc_hd__mux2_1
X_06455_ net746 _03111_ _03103_ _03104_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__o2bb2a_2
X_10565__217 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__inv_2
X_09174_ net217 net673 net276 net249 net2599 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout329_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06386_ top0.CPU.register.registers\[797\] top0.CPU.register.registers\[829\] top0.CPU.register.registers\[861\]
+ top0.CPU.register.registers\[893\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03043_
+ sky130_fd_sc_hd__mux4_1
X_08125_ net2778 net197 net430 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
XANTENNA__06513__S0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10606__258 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__inv_2
XANTENNA__09656__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08560__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ net497 net161 net701 net437 net2562 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout698_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
X_07007_ _03657_ _03662_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and2b_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
X_10459__111 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__inv_2
XANTENNA__07918__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__A3 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06816__S1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07394__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _04732_ net949 net699 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__or3b_1
XANTENNA__09135__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ net562 _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or2_1
X_08889_ net719 _04556_ _04764_ net283 net3268 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__a32o_1
XANTENNA__08343__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08894__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142__794 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__inv_2
X_12521_ net2213 _02160_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1014\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12452_ net2144 _02091_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[945\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08036__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ clknet_leaf_87_clk _01051_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08949__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ net2075 _02022_ net1094 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06504__S0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07621__A2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ net3437 net123 net116 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a21o_1
XANTENNA__08177__A3 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10147_ top0.display.delayctr\[24\] _05604_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__nand2_1
XANTENNA__09126__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ top0.display.delayctr\[9\] _05551_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__nand2_1
XANTENNA__07137__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08334__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08637__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08101__A3 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_31_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06743__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06240_ net731 _02894_ net739 vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a21o_1
XFILLER_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07860__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06171_ _02824_ _02827_ net779 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux2_1
Xhold315 top0.CPU.register.registers\[335\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 top0.CPU.register.registers\[741\] vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 top0.CPU.register.registers\[431\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__A2 _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06321__A1_N net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07073__A0 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09930_ _05422_ _05423_ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__o21a_1
Xhold337 top0.CPU.intMemAddr\[29\] vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 top0.CPU.register.registers\[803\] vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 top0.CPU.register.registers\[697\] vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout806 top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05736__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09861_ top0.CPU.internalMem.pcOut\[17\] _05361_ net647 vssd1 vssd1 vccd1 vccd1 _02194_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07376__A1 _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950__602 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__inv_2
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_4
Xfanout828 net834 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_2
X_09792_ _05272_ _05288_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__nand2_1
Xhold1015 net92 vssd1 vssd1 vccd1 vccd1 net3237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1004 top0.CPU.register.registers\[96\] vssd1 vssd1 vccd1 vccd1 net3226 sky130_fd_sc_hd__dlygate4sd3_1
X_08812_ _04718_ net307 net285 net2975 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a22o_1
Xhold1026 top0.CPU.register.registers\[271\] vssd1 vssd1 vccd1 vccd1 net3248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 top0.CPU.register.registers\[112\] vssd1 vssd1 vccd1 vccd1 net3270 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net202 net620 net320 net295 net2360 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__a32o_1
XANTENNA__09117__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 top0.CPU.register.registers\[858\] vssd1 vssd1 vccd1 vccd1 net3259 sky130_fd_sc_hd__dlygate4sd3_1
X_05955_ net776 _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__nand2_1
X_11085__737 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__inv_2
Xhold1059 top0.CPU.register.registers\[172\] vssd1 vssd1 vccd1 vccd1 net3281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout279_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_A _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06848__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08674_ net202 net698 net320 net299 net2264 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a32o_1
XANTENNA__06567__C _03222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05886_ net782 _02540_ net777 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o21a_1
XANTENNA__08340__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07625_ net470 _03318_ _03725_ net462 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__o211ai_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08628__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126__778 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__inv_2
X_07556_ _02869_ _03130_ _04144_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__or3b_1
XANTENNA__05785__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06507_ net766 _03161_ net754 vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout613_A _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09226_ top0.CPU.internalMem.pcOut\[22\] top0.CPU.internalMem.pcOut\[19\] top0.CPU.internalMem.pcOut\[18\]
+ top0.CPU.internalMem.pcOut\[16\] vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__or4_1
XANTENNA__06734__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ _02852_ net447 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__xnor2_1
X_06438_ _02497_ _02834_ _02870_ net541 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06369_ _03024_ _03025_ net763 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__mux2_1
X_09157_ net205 net3120 net248 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__mux2_1
X_08108_ net545 _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__nor2_1
X_09088_ net164 net615 net270 net255 net2465 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a32o_1
XANTENNA__08290__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359__1011 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__inv_2
XANTENNA_fanout982_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ net222 net704 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold871 top0.CPU.register.registers\[179\] vssd1 vssd1 vccd1 vccd1 net3093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold860 top0.CPU.register.registers\[220\] vssd1 vssd1 vccd1 vccd1 net3082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 top0.CPU.register.registers\[558\] vssd1 vssd1 vccd1 vccd1 net3104 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08797__Y _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693__345 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__inv_2
Xhold893 top0.CPU.register.registers\[917\] vssd1 vssd1 vccd1 vccd1 net3115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ _05484_ _05489_ net235 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__o21a_1
XFILLER_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09108__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_4_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10734__386 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__inv_2
XANTENNA__08867__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11952_ net1644 _01591_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[445\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11453__Q top0.CPU.decoder.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12776__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11883_ net1575 _01522_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[376\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08619__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12504_ net2196 _02143_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[997\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10628__280 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__inv_2
XANTENNA__11851__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12435_ net2127 _02074_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[928\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12366_ net2058 _02005_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07892__X _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05837__B _02493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ net1989 _01936_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[790\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05740_ net575 net634 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__nand2_2
XANTENNA__10114__B1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07410_ net482 _04061_ _04066_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__a21oi_1
X_08390_ _04655_ net397 net378 net2630 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07341_ net447 net535 _03129_ net534 net459 net467 vssd1 vssd1 vccd1 vccd1 _03998_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06716__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07294__A0 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ _02457_ net537 net446 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__or3_1
Xteam_07_1149 vssd1 vssd1 vccd1 vccd1 team_07_1149/HI gpio_out[15] sky130_fd_sc_hd__conb_1
X_06223_ top0.CPU.register.registers\[150\] top0.CPU.register.registers\[182\] top0.CPU.register.registers\[214\]
+ top0.CPU.register.registers\[246\] net838 net803 vssd1 vssd1 vccd1 vccd1 _02880_
+ sky130_fd_sc_hd__mux4_1
X_09011_ net210 net3039 net349 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_07_1138 vssd1 vssd1 vccd1 vccd1 team_07_1138/HI gpio_out[2] sky130_fd_sc_hd__conb_1
XANTENNA__11592__RESET_B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444__96 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__inv_2
X_06154_ _02473_ _02792_ net581 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a21o_1
Xhold101 top0.CPU.register.registers\[545\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 top0.CPU.register.registers\[357\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold123 top0.CPU.register.registers\[1008\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 top0.CPU.register.registers\[676\] vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06085_ _02740_ _02741_ net730 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
Xhold145 top0.CPU.register.registers\[333\] vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 top0.CPU.register.registers\[688\] vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
X_10677__329 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__inv_2
Xhold156 top0.CPU.register.registers\[448\] vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 top0.CPU.register.registers\[965\] vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 top0.CPU.register.registers\[713\] vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _04858_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_2
X_09913_ net588 _04530_ _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a21o_1
XANTENNA__07349__A1 _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout614 net618 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
Xfanout647 net649 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_4
X_09844_ net239 _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__nor2_1
Xfanout636 net637 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_2
XANTENNA__08546__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 _05133_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_2
XANTENNA__07349__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05763__A top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net670 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1211_A top0.CPU.intMem_out\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ top0.CPU.internalMem.pcOut\[10\] top0.CPU.internalMem.pcOut\[9\] _05254_
+ top0.CPU.internalMem.pcOut\[11\] vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__a31o_1
XFILLER_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06987_ net862 _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ net162 net3289 net358 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05938_ _02590_ _02591_ _02594_ net739 net771 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_29_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_A _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05869_ net737 _02525_ net773 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__o21ai_1
X_08657_ net162 net702 net309 net302 net2642 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32o_1
XFILLER_27_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07521__B2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07521__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ net490 _04000_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__nand2_1
XANTENNA__06955__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ net2969 net153 net334 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__mux2_1
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ _04134_ _04194_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08077__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09209_ _04583_ _04868_ _04869_ _04870_ _04867_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__o41a_1
XANTENNA__07037__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ net1912 _01859_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[713\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08785__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ net1843 _01790_ net972 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[644\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12082_ net1774 _01721_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[575\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11448__Q top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold690 top0.CPU.register.registers\[817\] vssd1 vssd1 vccd1 vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08537__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08968__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09145__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A3 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ net1627 _01574_ net1097 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[428\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11866_ net1558 _01505_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[359\]
+ sky130_fd_sc_hd__dfrtp_1
X_11797_ net1489 _01436_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[290\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08208__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ net2110 _02057_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08776__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ net2041 _01988_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[842\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08791__A3 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06910_ _03524_ net525 _03558_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__o21a_1
XANTENNA__08528__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07890_ net561 _04535_ _04536_ net625 vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__o211a_1
X_06841_ net864 _03493_ _03496_ _03497_ net860 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__o221a_1
XANTENNA__06398__B _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05988__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09560_ top0.CPU.Op\[6\] _02448_ _05107_ net643 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a31oi_1
XFILLER_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06772_ _02790_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__xnor2_2
XFILLER_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09491_ top0.MMIO.WBData_i\[2\] net139 vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__or2_1
X_08511_ net217 net683 net400 net367 net2374 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a32o_1
X_05723_ _02374_ _02377_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__nand2_1
X_11358__1010 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__inv_2
XFILLER_64_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08442_ net2772 net188 net375 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
XANTENNA__06937__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06027__A2_N _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08373_ net194 net709 net401 net383 net2542 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_63_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11197__849 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__inv_2
XANTENNA__08833__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ net533 net529 net469 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__mux2_1
XANTENNA__06165__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07255_ _03720_ _03911_ _03903_ _03900_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o211a_1
XANTENNA__07019__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06206_ top0.CPU.register.registers\[276\] top0.CPU.register.registers\[308\] top0.CPU.register.registers\[340\]
+ top0.CPU.register.registers\[372\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02863_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout409_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout311_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05912__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__A2 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ net578 _03842_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__nor2_1
X_06137_ top0.CPU.register.registers\[657\] top0.CPU.register.registers\[689\] top0.CPU.register.registers\[721\]
+ top0.CPU.register.registers\[753\] net828 net793 vssd1 vssd1 vccd1 vccd1 _02794_
+ sky130_fd_sc_hd__mux4_1
X_06068_ top0.CPU.register.registers\[394\] top0.CPU.register.registers\[426\] top0.CPU.register.registers\[458\]
+ top0.CPU.register.registers\[490\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02725_
+ sky130_fd_sc_hd__mux4_1
XFILLER_105_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 net406 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08519__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _04689_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 net435 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_4
Xfanout444 net446 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_2
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_2
Xfanout466 _02616_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_2
X_09827_ top0.CPU.internalMem.pcOut\[15\] _05328_ vssd1 vssd1 vccd1 vccd1 _05330_
+ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout945_A top0.CPU.control.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 net516 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_2
Xfanout488 _02554_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout477 _02577_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
X_09758_ top0.CPU.internalMem.pcOut\[9\] _05254_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__nand2_1
X_08709_ _04548_ _04743_ _04745_ net360 net3319 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__a32o_1
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09689_ _05189_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__nor2_1
XANTENNA__06152__A1_N net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06928__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ net1412 _01359_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ net1343 _01290_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10846__498 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__inv_2
X_11582_ net1274 _01221_ net1007 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08028__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05808__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05939__Y _02596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05903__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08758__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__Q top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10699__351 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__inv_2
X_12203_ net1895 _01842_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[696\]
+ sky130_fd_sc_hd__dfrtp_1
X_12134_ net1826 _01773_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[627\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09574__S _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ net1757 _01704_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[558\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09183__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08930__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__X _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09322__B top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ net1610 _01557_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[411\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_103_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ net1541 _01488_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08997__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload10 clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_6
X_07040_ top0.CPU.register.registers\[415\] top0.CPU.register.registers\[447\] top0.CPU.register.registers\[479\]
+ top0.CPU.register.registers\[511\] net851 net816 vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06472__A1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload43 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_16
Xclkload21 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_11_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload32 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__inv_16
Xclkload76 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_8
Xclkload54 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__inv_16
XANTENNA__08749__B1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload65 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__clkinv_8
X_10414__66 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__inv_2
XANTENNA__08213__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload87 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_2
Xclkload98 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__inv_6
X_08991_ net182 net696 net277 net260 net2568 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__a32o_1
X_07942_ top0.CPU.internalMem.pcOut\[13\] net642 _04580_ vssd1 vssd1 vccd1 vccd1 _04581_
+ sky130_fd_sc_hd__a21o_2
XANTENNA__05744__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07873_ net717 net207 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__and2_1
X_06824_ net752 _03480_ net747 vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06083__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09612_ net141 _05146_ net660 vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a21oi_1
X_10492__144 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__inv_2
X_09543_ net821 _05066_ net127 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
X_06755_ top0.CPU.register.registers\[655\] top0.CPU.register.registers\[687\] top0.CPU.register.registers\[719\]
+ top0.CPU.register.registers\[751\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ net132 net134 _05055_ net599 net3349 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__o32a_1
XANTENNA__05760__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10533__185 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06686_ _03341_ _03342_ net765 vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12647__Q top0.MMIO.WBData_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06386__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08425_ net2955 net211 net373 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ _04638_ net405 net384 net2755 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout526_A _03504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08988__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinvlp_4
X_07307_ net452 _03963_ _03843_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06138__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08563__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ net545 _02401_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__B _03989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ _02578_ _03893_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout895_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07169_ _03720_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__nor2_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08755__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ top0.display.delayctr\[30\] net664 net602 _05635_ _05634_ vssd1 vssd1 vccd1
+ vccd1 _02239_ sky130_fd_sc_hd__a221o_1
XANTENNA__06310__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout241 _05108_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_4
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08507__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09165__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07990__X _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_4
Xfanout252 _04822_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_4
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
Xfanout296 _04746_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07715__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__09180__A3 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08912__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11695__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05821__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06377__S1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12683_ clknet_leaf_82_clk _02318_ net1108 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
X_11703_ net1395 _01342_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[196\]
+ sky130_fd_sc_hd__dfrtp_1
X_11634_ net1326 _01273_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08691__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08979__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06129__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11565_ net1257 _01204_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11496_ clknet_leaf_91_clk net3356 net1085 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05888__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A_N _05162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07403__A0 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06301__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310__962 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__inv_2
X_12117_ net1809 _01756_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[610\]
+ sky130_fd_sc_hd__dfrtp_1
X_10476__128 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__inv_2
XFILLER_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ net1740 _01687_ net1081 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[541\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09156__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06065__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__Y _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06059__A1_N top0.CPU.control.funct7\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05812__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10517__169 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__inv_2
XFILLER_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06540_ net534 _03194_ _03195_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06368__S1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06471_ net745 _03127_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nand2_1
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08682__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08210_ net205 net682 vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__and2_1
X_09190_ net609 vssd1 vssd1 vccd1 vccd1 top0.CPU.addrControl sky130_fd_sc_hd__inv_2
XANTENNA__05800__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ net951 _02389_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nor2_4
Xclkload110 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload121 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10241__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ _04516_ net692 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__and2_1
X_07023_ _03678_ _03679_ net873 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06631__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ top0.CPU.register.registers\[180\] net565 vssd1 vssd1 vccd1 vccd1 _04788_
+ sky130_fd_sc_hd__or2_1
XANTENNA__05956__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold27 top0.CPU.register.registers\[31\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07925_ net633 _04566_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 top0.CPU.register.registers\[7\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 top0.CPU.register.registers\[39\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A1 top0.CPU.control.funct7\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 top0.CPU.register.registers\[816\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08558__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ net561 _04506_ _04507_ net625 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__o211a_1
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07787_ _03465_ _04298_ _03486_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a21bo_1
X_06807_ _03447_ net527 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__nor2_1
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ top0.CPU.Op\[4\] _05073_ net127 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
X_06738_ net864 _03390_ _03393_ _03394_ net860 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__o221a_1
X_09457_ top0.MMIO.WBData_i\[22\] _05041_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__and2_1
XANTENNA__08122__A1 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout810_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ net188 net694 net398 net379 net2684 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout908_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06669_ top0.CPU.register.registers\[769\] top0.CPU.register.registers\[801\] top0.CPU.register.registers\[833\]
+ top0.CPU.register.registers\[865\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03326_
+ sky130_fd_sc_hd__mux4_1
X_09388_ _04988_ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__or2_1
XANTENNA__08293__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ net3029 net410 net394 _04577_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a22o_1
X_11253__905 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__inv_2
XANTENNA__06107__A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10301_ _04938_ _05620_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__or2_1
XFILLER_4_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08189__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ net4 net653 net592 net3445 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
X_10163_ top0.display.delayctr\[27\] _05617_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__nand2_1
Xfanout1047 net1055 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_2
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
Xfanout1036 net1041 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_2
Xfanout1014 net1018 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08976__B net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__Q top0.CPU.control.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06047__S0 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ top0.display.delayctr\[13\] top0.display.delayctr\[14\] _05562_ vssd1 vssd1
+ vccd1 vccd1 _05566_ sky130_fd_sc_hd__or3_1
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12779__A top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1058 net1060 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05681__A top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__10299__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__A2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06598__S1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07225__X _03882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06496__B _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08113__A1 _04504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861__513 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06124__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ clknet_leaf_93_clk _02301_ net1081 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
X_12597_ clknet_leaf_89_clk _02232_ net1079 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07401__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08416__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ net1309 _01256_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_11548_ net1240 _01187_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_10902__554 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__inv_2
XANTENNA__06522__S1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 top0.CPU.register.registers\[472\] vssd1 vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 top0.CPU.register.registers\[478\] vssd1 vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ clknet_leaf_80_clk top0.CPU.busy net1113 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.prev_busy_o
+ sky130_fd_sc_hd__dfrtp_1
X_11037__689 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__inv_2
XANTENNA__09328__A _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09129__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06038__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08886__B net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1219 top0.CPU.intMem_out\[24\] vssd1 vssd1 vccd1 vccd1 net3441 sky130_fd_sc_hd__dlygate4sd3_1
X_07710_ _03621_ _03659_ _03664_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__a21boi_1
Xhold1208 top0.display.delayctr\[5\] vssd1 vssd1 vccd1 vccd1 net3430 sky130_fd_sc_hd__dlygate4sd3_1
X_05971_ net735 _02623_ _02626_ _02627_ net741 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_53_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07155__A2 _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ net164 net692 net311 net297 net2258 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__a32o_1
XFILLER_38_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08352__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07641_ _03570_ _04296_ _03466_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a21o_1
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07572_ net484 _04065_ _04227_ net476 _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__a221o_1
X_06523_ _03178_ _03179_ net762 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__mux2_1
XFILLER_81_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09311_ top0.display.delayctr\[1\] top0.display.delayctr\[18\] top0.display.delayctr\[19\]
+ top0.display.delayctr\[0\] vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__or4b_1
XANTENNA__08104__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ top0.CPU.intMemAddr\[1\] _04627_ net770 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__mux2_1
XANTENNA__06210__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06454_ _03107_ _03110_ net753 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XANTENNA__08407__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ net179 net674 net278 net249 net2710 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__a32o_1
X_06385_ top0.CPU.register.registers\[925\] top0.CPU.register.registers\[957\] top0.CPU.register.registers\[989\]
+ top0.CPU.register.registers\[1021\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03042_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10214__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ net2973 _04566_ net430 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout224_A _04492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645__297 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__inv_2
XANTENNA__08841__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ net493 net165 net701 net437 net2468 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a32o_1
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07006_ _03638_ _03660_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout593_A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10498__150 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__inv_2
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07981__A _04127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05929__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout760_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ net155 net705 net273 net264 net2353 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__a32o_1
XANTENNA__08288__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ top0.CPU.register.registers\[242\] net571 net560 vssd1 vssd1 vccd1 vccd1
+ _04764_ sky130_fd_sc_hd__o21a_1
X_07908_ _04342_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__and3_1
X_10539__191 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__inv_2
XANTENNA__09540__A0 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07839_ net2905 net549 net503 _04493_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a22o_1
XFILLER_72_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09260__X _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09509_ _02336_ _02352_ top0.MMIO.WBData_i\[14\] top0.MMIO.WBData_i\[20\] net148
+ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__o41a_1
XANTENNA__08646__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06201__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ net2212 _02159_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1013\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ net2143 _02090_ net1013 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[944\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08036__B _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ clknet_leaf_86_clk _01050_ net1091 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09071__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ net2074 _02021_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[875\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10215_ net3238 net122 _05644_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a21o_1
XFILLER_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07385__A2 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ top0.display.delayctr\[24\] _05604_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__or2_1
XFILLER_0_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10077_ top0.display.delayctr\[9\] _05551_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__or2_1
XFILLER_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08885__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06440__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08098__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09611__A _02683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06743__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12649_ clknet_leaf_66_clk _02284_ net1104 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_06170_ _02825_ _02826_ net729 vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09062__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06970__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08270__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 top0.CPU.register.registers\[586\] vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 top0.CPU.register.registers\[831\] vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07073__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold327 top0.CPU.register.registers\[426\] vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold349 top0.CPU.register.registers\[71\] vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 top0.CPU.register.registers\[630\] vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
X_09860_ _05357_ _05358_ _05359_ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__o22ai_1
Xfanout807 net809 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06259__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08573__A1 _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net819 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05736__D net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout829 net831 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_4
X_09791_ _05246_ _05251_ _05263_ _05295_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__and4_1
X_08811_ net202 net673 net320 net287 net2797 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a32o_1
Xhold1005 top0.CPU.register.registers\[135\] vssd1 vssd1 vccd1 vccd1 net3227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08742_ _04684_ net328 net296 net2844 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__a22o_1
XANTENNA__09505__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1016 net58 vssd1 vssd1 vccd1 vccd1 net3238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 top0.CPU.register.registers\[66\] vssd1 vssd1 vccd1 vccd1 net3249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 top0.CPU.register.registers\[983\] vssd1 vssd1 vccd1 vccd1 net3260 sky130_fd_sc_hd__dlygate4sd3_1
X_05954_ _02609_ _02610_ net724 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
Xhold1049 top0.CPU.register.registers\[257\] vssd1 vssd1 vccd1 vccd1 net3271 sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ _04665_ net327 net300 net2676 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07128__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__C_N net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_A _04611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ _04277_ _04278_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__and3_1
X_05885_ net726 _02541_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__or2_1
XANTENNA__06431__S0 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ _02852_ _03150_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nand2b_1
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06506_ net873 _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout439_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__B _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07486_ _03928_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1083_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ top0.CPU.internalMem.pcOut\[21\] top0.CPU.internalMem.pcOut\[20\] top0.CPU.internalMem.pcOut\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__or3_1
XANTENNA__06734__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06437_ _03078_ net537 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout606_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06880__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06368_ top0.CPU.register.registers\[542\] top0.CPU.register.registers\[574\] top0.CPU.register.registers\[606\]
+ top0.CPU.register.registers\[638\] net937 net903 vssd1 vssd1 vccd1 vccd1 _03025_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07976__A _04106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__B2 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ _04714_ net269 net247 net3133 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a22o_1
XANTENNA__08571__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08107_ net954 net953 net951 net948 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__or4bb_1
XANTENNA__08800__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ net213 net615 net270 net255 net2602 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_110_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06299_ net735 _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__or2_1
XANTENNA__08143__Y _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08038_ net508 net203 net707 net438 net2441 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a32o_1
XANTENNA__06811__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08013__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold872 top0.display.dataforOutput\[10\] vssd1 vssd1 vccd1 vccd1 net3094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 net85 vssd1 vssd1 vccd1 vccd1 net3083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold850 top0.CPU.register.registers\[317\] vssd1 vssd1 vccd1 vccd1 net3072 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _05484_ _05489_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__nand2_1
Xhold883 top0.CPU.register.registers\[724\] vssd1 vssd1 vccd1 vccd1 net3105 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08564__A1 _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 top0.CPU.register.registers\[384\] vssd1 vssd1 vccd1 vccd1 net3116 sky130_fd_sc_hd__dlygate4sd3_1
X_10375__27 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__inv_2
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _05462_ _05473_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06670__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ net1643 _01590_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[444\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06120__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06422__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11882_ net1574 _01521_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[375\]
+ sky130_fd_sc_hd__dfrtp_1
X_11259__911 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__inv_2
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_43_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08095__A3 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ net2195 _02142_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[996\]
+ sky130_fd_sc_hd__dfrtp_1
X_12434_ net2126 _02073_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[927\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05958__X _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06790__A _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12365_ net2057 _02004_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06489__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973__625 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__inv_2
XFILLER_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ net1988 _01935_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_122_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08004__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06566__B1 _03222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _02850_ net551 vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10114__A1 _02493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06413__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07340_ net488 _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__nand2_1
XANTENNA__08086__A3 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06716__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908__560 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07271_ _02457_ _03092_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__xnor2_1
X_09010_ net211 net613 _04799_ net349 net3256 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__a32o_1
XANTENNA__08491__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07294__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1139 vssd1 vssd1 vccd1 vccd1 team_07_1139/HI gpio_out[5] sky130_fd_sc_hd__conb_1
X_06222_ net780 _02874_ _02878_ net771 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__o211a_1
X_06153_ net579 _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or2_1
Xhold113 top0.CPU.register.registers\[749\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 top0.CPU.register.registers\[328\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 top0.CPU.register.registers\[720\] vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 top0.CPU.register.registers\[870\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 top0.CPU.register.registers\[746\] vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_11052__704 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__inv_2
X_06084_ top0.CPU.register.registers\[13\] top0.CPU.register.registers\[45\] top0.CPU.register.registers\[77\]
+ top0.CPU.register.registers\[109\] net849 net814 vssd1 vssd1 vccd1 vccd1 _02741_
+ sky130_fd_sc_hd__mux4_1
Xhold157 top0.CPU.register.registers\[616\] vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 top0.CPU.register.registers\[850\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 top0.CPU.register.registers\[620\] vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net586 _02871_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__nor2_1
Xfanout604 _04856_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_4
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
XANTENNA__06699__X _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout637 _02395_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08420__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 net649 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09743__B1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _05338_ _05341_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a21boi_2
Xfanout626 _02420_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout291_A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _05133_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout389_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07036__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__inv_2
XANTENNA__06211__Y _02868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06986_ _03641_ _03642_ net756 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout556_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ net164 net3178 net358 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__mux2_1
XFILLER_39_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05937_ _02592_ _02593_ net731 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__mux2_1
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05868_ _02523_ _02524_ net784 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XANTENNA__06404__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ net164 net703 net310 net301 net2575 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a32o_1
XANTENNA__08566__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07521__A2 _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ _04261_ _04263_ net448 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__o21a_1
X_08587_ net2906 net159 net333 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__mux2_1
XANTENNA__06955__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05799_ net781 net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_81_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07538_ _02962_ _03637_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_40_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ _04113_ _04123_ _04125_ _04121_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__a211o_1
XANTENNA__08482__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ _04568_ _04573_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__or2_1
X_10660__312 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__inv_2
XANTENNA__07037__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957__609 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__inv_2
XANTENNA__08234__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ net164 net680 net270 net251 net2452 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__X _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12150_ net1842 _01789_ net995 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[643\]
+ sky130_fd_sc_hd__dfrtp_1
X_10701__353 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__inv_2
XANTENNA__06115__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12081_ net1773 _01720_ net1050 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[574\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_92_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 top0.CPU.register.registers\[480\] vssd1 vssd1 vccd1 vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 top0.CPU.register.registers\[780\] vssd1 vssd1 vccd1 vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06769__B net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11464__Q top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ net1626 _01573_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[427\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05960__Y _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11865_ net1557 _01504_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[358\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11796_ net1488 _01435_ net962 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[289\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08473__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07028__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08225__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net2109 _02056_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07579__A2 _03379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ net2040 _01987_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[841\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07984__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net1971 _01918_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[772\]
+ sky130_fd_sc_hd__dfrtp_1
X_06840_ net760 _03494_ net751 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a21o_1
XANTENNA__06539__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06771_ net246 _02771_ net543 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ top0.MMIO.WBData_i\[9\] net137 vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or2_1
X_08510_ net179 net685 net401 net368 net2471 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a32o_1
X_05722_ _02374_ _02377_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__and2_1
X_08441_ net2946 net192 net376 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__mux2_1
XANTENNA__05803__S net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06937__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07303__B _03173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08372_ _04651_ net394 net382 net2590 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
XANTENNA__08464__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07323_ net534 _03221_ net469 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__mux2_1
X_07254_ _03907_ _03910_ net487 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__mux2_1
XANTENNA__07019__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06205_ net777 _02857_ _02860_ _02861_ net772 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__o221a_1
X_07185_ net518 _03745_ _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o21a_1
XFILLER_105_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06136_ _02473_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__and2_1
XANTENNA__08231__A3 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06067_ top0.CPU.register.registers\[266\] top0.CPU.register.registers\[298\] top0.CPU.register.registers\[330\]
+ top0.CPU.register.registers\[362\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02724_
+ sky130_fd_sc_hd__mux4_1
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout412 _04721_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_4
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
Xfanout401 net403 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_4
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
XANTENNA_fanout673_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_2
Xfanout456 _02617_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_2
X_09826_ top0.CPU.internalMem.pcOut\[15\] _05328_ vssd1 vssd1 vccd1 vccd1 _05329_
+ sky130_fd_sc_hd__or2_1
XFILLER_100_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout478 _02575_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_2
Xfanout467 _02598_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_4
X_09757_ _05263_ _05264_ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__o21a_1
XFILLER_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06969_ _03624_ _03625_ net765 vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__mux2_1
X_08708_ top0.CPU.register.registers\[403\] net575 vssd1 vssd1 vccd1 vccd1 _04745_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout938_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08296__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180__832 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__inv_2
X_09688_ _05180_ _05182_ _05190_ _05179_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__o211a_1
XFILLER_82_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06928__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ _04648_ net312 net301 net2991 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11650_ net1342 _01289_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[143\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07988__X _04618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11581_ net1273 _01220_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_11221__873 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__inv_2
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08470__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08222__A3 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ net1894 _01841_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[695\]
+ sky130_fd_sc_hd__dfrtp_1
X_12133_ net1825 _01772_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[626\]
+ sky130_fd_sc_hd__dfrtp_1
X_12064_ net1756 _01703_ net1044 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05684__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout990 net992 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_121_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08219__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11917_ net1609 _01556_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[410\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_103_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07898__X _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11848_ net1540 _01487_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[341\]
+ sky130_fd_sc_hd__dfrtp_1
X_11779_ net1471 _01418_ net1035 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[272\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05859__A _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06962__B net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06454__S net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979__631 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__inv_2
Xclkload11 clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_8
XANTENNA__06026__Y _02683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload44 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__clkinv_16
Xclkload22 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_11_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload33 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__inv_16
Xclkload77 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_8
Xclkload55 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_16
Xclkload66 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_2
XANTENNA__06855__S0 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload99 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload88 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__inv_2
XANTENNA__08241__Y _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ net187 net694 _04794_ net260 net3081 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__a32o_1
X_07941_ net562 _04578_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__o21a_1
XANTENNA__10308__A1 _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ top0.CPU.internalMem.pcOut\[24\] net641 net635 _04521_ vssd1 vssd1 vccd1
+ vccd1 _04522_ sky130_fd_sc_hd__o211a_2
XANTENNA__07185__B1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06823_ _03478_ _03479_ net762 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
XANTENNA__06083__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _02683_ _05007_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__or2_1
XFILLER_56_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09542_ net856 _05068_ net127 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
X_06754_ _02515_ _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164__816 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__inv_2
X_05705_ top0.MISOtoMMIO\[4\] vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout254_A _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ top0.MMIO.WBData_i\[30\] net146 net135 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_90_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
X_11205__857 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06685_ top0.CPU.register.registers\[512\] top0.CPU.register.registers\[544\] top0.CPU.register.registers\[576\]
+ top0.CPU.register.registers\[608\] net921 net887 vssd1 vssd1 vccd1 vccd1 _03342_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08844__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ net2970 _04492_ net374 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__mux2_1
X_08355_ net151 net709 net404 net383 net2974 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a32o_1
Xclkload5 clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout519_A _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A _04689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ net489 _03953_ _03962_ _03948_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a22oi_2
XANTENNA__08145__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058__710 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__inv_2
X_08286_ net495 net153 net671 net417 net2399 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a32o_1
XANTENNA__07660__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07237_ net347 _03893_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__nor2_1
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07168_ _03816_ _03824_ net487 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__mux2_1
XFILLER_3_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout790_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06846__S0 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06119_ _02774_ _02775_ net733 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout888_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ net486 _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout220 _04603_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout231 _04471_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10772__424 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__inv_2
Xfanout253 net254 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout264 _04772_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_8
X_09809_ top0.CPU.internalMem.pcOut\[12\] _05280_ top0.CPU.internalMem.pcOut\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout286 _04750_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_8
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_4
XFILLER_47_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout275 net281 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
XANTENNA__08912__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10813__465 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__inv_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05821__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08676__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xclkbuf_leaf_81_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
X_12682_ clknet_leaf_82_clk _02317_ net1108 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
X_11702_ net1394 _01341_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[195\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08039__B net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11633_ net1325 _01272_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08691__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06274__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11564_ net1256 _01203_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11495_ clknet_leaf_91_clk _01134_ net1084 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05888__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07403__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12116_ net1808 _01755_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[609\]
+ sky130_fd_sc_hd__dfrtp_1
X_12047_ net1739 _01686_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[540\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07118__B net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06065__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09614__A _02665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05861__B _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05812__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07014__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_72_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
X_06470_ _03123_ _03124_ _03125_ _03126_ net759 net862 vssd1 vssd1 vccd1 vccd1 _03127_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07890__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08140_ net2683 net154 net432 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XANTENNA__09092__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06184__S net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload111 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__inv_16
Xclkload122 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__inv_8
XANTENNA__07642__A1 _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload100 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__clkinv_1
X_08071_ net2759 net433 _04658_ net491 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a22o_1
X_07022_ top0.CPU.register.registers\[415\] top0.CPU.register.registers\[447\] top0.CPU.register.registers\[479\]
+ top0.CPU.register.registers\[511\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__mux4_1
XFILLER_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10756__408 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__inv_2
XANTENNA__05956__A1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _04663_ net555 _04787_ net262 net3066 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__a32o_1
X_07924_ top0.CPU.internalMem.pcOut\[16\] net642 _04564_ _04565_ vssd1 vssd1 vccd1
+ vccd1 _04566_ sky130_fd_sc_hd__a22o_2
Xhold17 top0.CPU.register.registers\[16\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_71_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500__152 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__inv_2
Xhold28 top0.CPU.register.registers\[1\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 top0.CPU.register.registers\[191\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08839__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ net591 _02928_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__nand2_1
X_06806_ net748 _03462_ _03451_ _03455_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__o2bb2a_2
X_07786_ _03464_ _03486_ _04298_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or3b_1
XFILLER_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09525_ top0.CPU.Op\[3\] _05085_ net127 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06737_ net760 _03391_ net751 vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a21o_1
XANTENNA__08658__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ net132 net134 _05046_ net599 net3432 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_63_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout636_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ _03323_ _03324_ net756 vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__mux2_1
X_08407_ net192 net699 net407 net380 net2665 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ top0.CPU.control.funct3\[2\] _02409_ top0.CPU.control.funct3\[0\] vssd1 vssd1
+ vccd1 vccd1 _04999_ sky130_fd_sc_hd__mux2_1
X_06599_ top0.CPU.register.registers\[263\] top0.CPU.register.registers\[295\] top0.CPU.register.registers\[327\]
+ top0.CPU.register.registers\[359\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03256_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout803_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08338_ net721 net197 net404 net411 net2648 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a32o_1
XANTENNA__09083__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ net507 net199 net672 net419 net2271 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a32o_1
X_11292__944 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__inv_2
XANTENNA__08830__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06841__C1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ net3341 net118 net111 _05669_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
X_10231_ net3 net656 net595 top0.MMIO.WBData_i\[10\] vssd1 vssd1 vccd1 vccd1 _02277_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333__985 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__inv_2
XANTENNA__07936__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1004 net1132 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
X_10162_ _04957_ _05620_ net661 vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__o21a_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1026 net1030 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
Xfanout1015 net1017 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
X_10093_ top0.display.delayctr\[13\] net665 net603 _05565_ _05165_ vssd1 vssd1 vccd1
+ vccd1 _02222_ sky130_fd_sc_hd__a221o_1
Xfanout1048 net1050 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07653__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1060 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08897__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06047__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08361__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11472__Q top0.CPU.control.funct7\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06124__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07321__A0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__A1 top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12665_ clknet_leaf_92_clk _02300_ net1082 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
X_11616_ net1308 _01255_ net1030 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09613__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ clknet_leaf_89_clk _02231_ net1087 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09074__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08416__A3 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10941__593 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__inv_2
XANTENNA__08821__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11547_ net1239 _01186_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[40\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold509 top0.CPU.register.registers\[490\] vssd1 vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
X_11478_ clknet_leaf_77_clk top0.CPU.internalMem.state_n\[3\] net1123 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.state\[3\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09328__B _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06060__B1 top0.CPU.control.funct7\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05970_ net782 _02624_ net776 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__o21a_1
XANTENNA__05938__B2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1209 top0.display.delayctr\[26\] vssd1 vssd1 vccd1 vccd1 net3431 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06038__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08888__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _03466_ _03570_ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__nand3_1
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07571_ net337 _04224_ _03841_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_45_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06522_ top0.CPU.register.registers\[530\] top0.CPU.register.registers\[562\] top0.CPU.register.registers\[594\]
+ top0.CPU.register.registers\[626\] net931 net897 vssd1 vssd1 vccd1 vccd1 _03179_
+ sky130_fd_sc_hd__mux4_1
X_09310_ top0.display.delayctr\[2\] top0.display.delayctr\[3\] top0.display.delayctr\[5\]
+ top0.display.delayctr\[6\] vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__or4_1
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08655__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11276__928 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__inv_2
X_09241_ top0.CPU.internalMem.pcOut\[4\] _04902_ net609 vssd1 vssd1 vccd1 vccd1 _04903_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07863__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06210__S1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06453_ _03108_ _03109_ net764 vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
X_09172_ net183 net676 net277 net249 net2855 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a32o_1
X_06384_ _03005_ _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09065__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ net2890 _04561_ net431 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11020__672 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__inv_2
XANTENNA_fanout217_A _04603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317__969 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__inv_2
X_08054_ net497 net215 net702 net437 net2431 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a32o_1
XANTENNA__08812__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07005_ _03640_ net520 vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__nand2_1
XANTENNA__06642__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07918__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05929__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07394__A3 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ net157 net701 net267 net263 net2447 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a32o_1
X_07907_ net3059 net549 net515 _04551_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
X_08887_ _04551_ net560 _04763_ net284 net3208 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ net723 net224 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__and2_1
XANTENNA__08894__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05788__S0 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ top0.MMIO.WBData_i\[16\] net138 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_36_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07769_ _02869_ _03129_ net445 _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o31ai_1
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884__536 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09439_ net3405 net597 net130 _05035_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__o22a_1
XANTENNA__06201__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925__577 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__inv_2
X_12450_ net2142 _02089_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[943\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09056__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__C net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11401_ clknet_leaf_57_clk _01049_ net1092 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12381_ net2073 _02020_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[874\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08803__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10778__430 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__inv_2
XFILLER_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09148__B _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ net2872 net123 net116 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a21o_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10145_ _02906_ _05577_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__nor2_1
X_10819__471 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__inv_2
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10076_ net3369 net665 net136 _05553_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a211o_1
XFILLER_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08334__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05779__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06440__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07115__C net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ clknet_leaf_65_clk _02283_ net1102 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11004__656 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__inv_2
XANTENNA__09047__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ clknet_leaf_90_clk _02214_ net1085 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold306 top0.CPU.register.registers\[63\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08243__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__A _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold317 top0.CPU.register.registers\[329\] vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 top0.CPU.register.registers\[879\] vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 top0.CPU.intMemAddr\[8\] vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06259__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ _04717_ net328 net288 net2786 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a22o_1
Xfanout819 top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_2
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
Xhold1006 top0.CPU.register.registers\[133\] vssd1 vssd1 vccd1 vccd1 net3228 sky130_fd_sc_hd__dlygate4sd3_1
X_09790_ _05251_ _05263_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nand3_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06584__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1039 top0.CPU.register.registers\[83\] vssd1 vssd1 vccd1 vccd1 net3261 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _04683_ net321 net295 net2668 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a22o_1
Xhold1028 net93 vssd1 vssd1 vccd1 vccd1 net3250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 top0.CPU.register.registers\[721\] vssd1 vssd1 vccd1 vccd1 net3239 sky130_fd_sc_hd__dlygate4sd3_1
X_05953_ top0.CPU.register.registers\[257\] top0.CPU.register.registers\[289\] top0.CPU.register.registers\[321\]
+ top0.CPU.register.registers\[353\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02610_
+ sky130_fd_sc_hd__mux4_1
X_08672_ _04664_ net312 net297 net2769 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a22o_1
X_10571__223 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__inv_2
X_05884_ top0.CPU.register.registers\[899\] top0.CPU.register.registers\[931\] top0.CPU.register.registers\[963\]
+ top0.CPU.register.registers\[995\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02541_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08325__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ _03359_ net344 _04279_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout167_A _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_18_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06431__S1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07554_ _02889_ _03112_ _03928_ _04210_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a31o_1
X_10612__264 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__inv_2
X_06505_ top0.CPU.register.registers\[915\] top0.CPU.register.registers\[947\] top0.CPU.register.registers\[979\]
+ top0.CPU.register.registers\[1011\] net940 net906 vssd1 vssd1 vccd1 vccd1 _03162_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07836__A1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07485_ _04140_ _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__nand2b_1
X_09224_ top0.CPU.internalMem.pcOut\[30\] top0.CPU.internalMem.pcOut\[29\] top0.CPU.internalMem.pcOut\[28\]
+ top0.CPU.internalMem.pcOut\[27\] vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__or4_1
XANTENNA__09038__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06436_ _03078_ net537 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout334_A _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12555__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08852__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05942__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06367_ top0.CPU.register.registers\[670\] top0.CPU.register.registers\[702\] top0.CPU.register.registers\[734\]
+ top0.CPU.register.registers\[766\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03024_
+ sky130_fd_sc_hd__mux4_1
X_09155_ _04713_ net273 net248 net2541 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ net167 net621 net277 net257 net2510 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a32o_1
XFILLER_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06298_ _02953_ _02954_ net783 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__mux2_1
X_08106_ net502 net154 net693 net436 net2563 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a32o_1
X_08037_ net2968 net440 _04649_ net515 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a22o_1
Xhold873 _01141_ vssd1 vssd1 vccd1 vccd1 net3095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 net96 vssd1 vssd1 vccd1 vccd1 net3084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 top0.CPU.register.registers\[593\] vssd1 vssd1 vccd1 vccd1 net3073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold840 top0.CPU.register.registers\[641\] vssd1 vssd1 vccd1 vccd1 net3062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 top0.CPU.register.registers\[900\] vssd1 vssd1 vccd1 vccd1 net3117 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A top0.CPU.decoder.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold884 top0.CPU.register.registers\[910\] vssd1 vssd1 vccd1 vccd1 net3106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ top0.CPU.internalMem.pcOut\[27\] net645 _05478_ vssd1 vssd1 vccd1 vccd1 _02204_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08299__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08939_ _04651_ net274 net264 net3069 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__a22o_1
XANTENNA__06670__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ net1642 _01589_ net992 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09271__X _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06422__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ net1573 _01520_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[374\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08619__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11298__950 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09029__A0 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06186__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ net2194 _02141_ net988 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[995\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12433_ net2125 _02072_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[926\]
+ sky130_fd_sc_hd__dfrtp_1
X_11339__991 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__inv_2
XFILLER_8_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05687__A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08252__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12364_ net2056 _02003_ net984 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06489__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12295_ net1987 _01934_ net1038 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[788\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08004__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555__207 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__inv_2
XANTENNA__09606__B _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10128_ net3409 net667 _05141_ _05590_ _05593_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a221o_1
XANTENNA__06311__A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ _05539_ _05540_ net600 vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_50_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09622__A _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06413__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07270_ _03754_ _03926_ _03925_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__o21a_1
X_10449__101 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06221_ net739 _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__or2_1
XANTENNA__05924__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06152_ net741 _02808_ _02797_ _02801_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__o2bb2a_2
Xhold114 top0.CPU.register.registers\[767\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 top0.CPU.register.registers\[639\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
X_06083_ top0.CPU.register.registers\[141\] top0.CPU.register.registers\[173\] top0.CPU.register.registers\[205\]
+ top0.CPU.register.registers\[237\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02740_
+ sky130_fd_sc_hd__mux4_1
Xhold103 top0.CPU.register.registers\[1000\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11091__743 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__inv_2
Xhold136 top0.CPU.register.registers\[709\] vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 top0.CPU.register.registers\[959\] vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 top0.CPU.register.registers\[973\] vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ top0.CPU.internalMem.pcOut\[21\] _05407_ net647 vssd1 vssd1 vccd1 vccd1 _02198_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold169 top0.CPU.register.registers\[1004\] vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout605 _04856_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_2
XANTENNA__11948__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout649 net651 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_2
X_09842_ top0.CPU.internalMem.pcOut\[16\] _05343_ vssd1 vssd1 vccd1 vccd1 _05344_
+ sky130_fd_sc_hd__xor2_1
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_2
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_2
XANTENNA__08546__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 net618 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_2
X_11132__784 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__inv_2
X_09773_ top0.CPU.internalMem.pcOut\[11\] top0.CPU.internalMem.pcOut\[10\] top0.CPU.internalMem.pcOut\[9\]
+ _05254_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__and4_1
XFILLER_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06221__A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_A _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ net214 net3345 net357 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__mux2_1
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06985_ top0.CPU.register.registers\[538\] top0.CPU.register.registers\[570\] top0.CPU.register.registers\[602\]
+ top0.CPU.register.registers\[634\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03642_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_4_7_0_clk_X clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05936_ top0.CPU.register.registers\[0\] top0.CPU.register.registers\[32\] top0.CPU.register.registers\[64\]
+ top0.CPU.register.registers\[96\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02593_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09510__A4 top0.MMIO.WBData_i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05867_ top0.CPU.register.registers\[907\] top0.CPU.register.registers\[939\] top0.CPU.register.registers\[971\]
+ top0.CPU.register.registers\[1003\] net844 net809 vssd1 vssd1 vccd1 vccd1 _02524_
+ sky130_fd_sc_hd__mux4_1
X_08655_ net214 net702 net310 net302 net2727 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout451_A _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06404__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07606_ net337 _04093_ _04262_ net476 vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__a22o_1
X_08586_ net2924 net161 net333 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__mux2_1
X_05798_ _02447_ _02449_ _02452_ _02341_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_81_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07537_ _02909_ _03617_ _04135_ _02926_ _03600_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a32o_1
XFILLER_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06891__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _02650_ _04119_ _04124_ net443 vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__a22o_1
X_09207_ _04541_ _04557_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06419_ _03074_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__or2_1
X_07399_ _03905_ _03909_ net479 vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__mux2_1
XFILLER_6_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10996__648 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__inv_2
XANTENNA__08234__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ net3292 net251 _04839_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a21o_1
X_10435__87 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__inv_2
XANTENNA__08785__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07993__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ net202 _04670_ _04816_ net258 net3278 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__a32o_1
X_10740__392 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ net1772 _01719_ net1082 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[573\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11689__RESET_B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 top0.CPU.register.registers\[768\] vssd1 vssd1 vccd1 vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold670 top0.CPU.register.registers\[149\] vssd1 vssd1 vccd1 vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08537__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 top0.CPU.register.registers\[646\] vssd1 vssd1 vccd1 vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09145__C _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06131__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ net1625 _01572_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[426\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ net1556 _01503_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11795_ net1487 _01434_ net1065 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[288\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05906__S0 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10280__B2 _05168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07681__C1 _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ net2108 _02055_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[909\]
+ sky130_fd_sc_hd__dfrtp_1
X_11075__727 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__inv_2
XANTENNA__08776__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ net2039 _01986_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116__768 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__inv_2
X_12278_ net1970 _01917_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[771\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10356__8 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06770_ _03426_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__inv_2
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05721_ top0.CPU.Op\[0\] top0.CPU.Op\[1\] top0.CPU.Op\[2\] vssd1 vssd1 vccd1 vccd1
+ _02378_ sky130_fd_sc_hd__nand3_2
XFILLER_36_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08440_ net2882 _04581_ net375 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06187__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08371_ net197 net711 net404 net383 net2479 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_63_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10683__335 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__inv_2
X_07322_ _03977_ _03978_ net458 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__mux2_1
XFILLER_137_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07253_ _03908_ _03909_ net346 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__mux2_1
XANTENNA__06570__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06204_ net729 _02858_ net740 vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a21o_1
X_07184_ net450 _03742_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nand2_4
XANTENNA__09413__B1 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06135_ net873 _02474_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__nand2_1
XANTENNA__09964__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724__376 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__inv_2
XANTENNA__07975__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06066_ _02719_ _02720_ _02721_ _02722_ net728 net738 vssd1 vssd1 vccd1 vccd1 _02723_
+ sky130_fd_sc_hd__mux4_1
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
XANTENNA_fanout499_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08519__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_4
Xfanout424 _04689_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_4
X_09825_ _02513_ _04568_ net587 vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__mux2_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout446 _03739_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_2
Xfanout457 _02617_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout479 _02575_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_2
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
X_10618__270 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__inv_2
X_09756_ _05263_ _05264_ net241 vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08577__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ top0.CPU.register.registers\[539\] top0.CPU.register.registers\[571\] top0.CPU.register.registers\[603\]
+ top0.CPU.register.registers\[635\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03625_
+ sky130_fd_sc_hd__mux4_1
X_09687_ _05199_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__and2b_1
X_08707_ net223 net3285 net358 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_05919_ net480 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__inv_2
X_06899_ net747 _03555_ _03550_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _04647_ net315 net302 net3026 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a22o_1
XANTENNA__06389__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net3177 _04548_ net336 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11580_ net1272 _01219_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06561__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ net1893 _01840_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08758__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ net1824 _01771_ net991 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[625\]
+ sky130_fd_sc_hd__dfrtp_1
X_12063_ net1755 _01702_ net1102 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[556\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09183__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08930__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09608__B1_N _02649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ net1608 _01555_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[409\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10667__319 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ net1539 _01486_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ net1470 _01417_ net1047 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05859__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08997__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06552__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload12 clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload23 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_8
Xclkload34 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_11_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload56 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_8
Xclkload78 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_2
XANTENNA__08749__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload67 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_4
XANTENNA__10005__B2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload45 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload89 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__inv_4
XANTENNA__09066__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06855__S1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ top0.CPU.intMem_out\[13\] net625 _02734_ _02386_ net639 vssd1 vssd1 vccd1
+ vccd1 _04579_ sky130_fd_sc_hd__o221a_1
XFILLER_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10308__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09174__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ top0.CPU.intMem_out\[24\] net627 _04520_ net643 vssd1 vssd1 vccd1 vccd1 _04521_
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07185__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ top0.CPU.register.registers\[269\] top0.CPU.register.registers\[301\] top0.CPU.register.registers\[333\]
+ top0.CPU.register.registers\[365\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03479_
+ sky130_fd_sc_hd__mux4_1
X_09610_ top0.display.dataforOutput\[4\] net604 net658 net3355 _05145_ vssd1 vssd1
+ vccd1 vccd1 _01135_ sky130_fd_sc_hd__a221o_1
XFILLER_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09541_ net861 _05076_ net128 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XFILLER_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06753_ net246 _02771_ _02790_ net543 vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05704_ top0.CPU.internalMem.loadCt\[2\] vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__inv_2
X_09472_ net132 net134 _05054_ net599 net3433 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__o32a_1
X_11244__896 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__inv_2
XFILLER_64_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06684_ top0.CPU.register.registers\[640\] top0.CPU.register.registers\[672\] top0.CPU.register.registers\[704\]
+ top0.CPU.register.registers\[736\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03341_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_19_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ net3240 _04487_ net376 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__mux2_1
XANTENNA__06791__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ net949 net545 net711 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or3b_1
XANTENNA__08437__A1 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09021__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ net489 _03837_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__nor2_1
XANTENNA__08145__B net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload6 clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout414_A _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08285_ net491 net159 net668 net417 net2632 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a32o_1
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08860__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07236_ _03053_ net518 net538 net539 net456 net473 vssd1 vssd1 vccd1 vccd1 _03893_
+ sky130_fd_sc_hd__mux4_1
XFILLER_119_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07167_ _03819_ _03823_ net346 vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
X_10405__57 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__inv_2
XFILLER_133_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138__790 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__inv_2
X_06118_ top0.CPU.register.registers\[526\] top0.CPU.register.registers\[558\] top0.CPU.register.registers\[590\]
+ top0.CPU.register.registers\[622\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02775_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07329__X _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06846__S1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ _02428_ _02431_ _03710_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__or3_2
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
X_06049_ net728 _02703_ net737 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a21o_1
Xfanout210 _04504_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout221 _04576_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout254 _04822_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_4
XANTENNA_fanout950_A top0.CPU.decoder.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09165__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08373__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ top0.CPU.internalMem.pcOut\[13\] top0.CPU.internalMem.pcOut\[12\] _05280_
+ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__and3_1
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 net300 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_8
X_09739_ net631 _04601_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__o21bai_1
XFILLER_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06923__B2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_38_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12681_ clknet_leaf_92_clk _02316_ net1084 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
X_11701_ net1393 _01340_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[194\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11632_ net1324 _01271_ net1079 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06782__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08428__A1 _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09625__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ net1255 _01202_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ clknet_leaf_90_clk net3351 net1086 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07403__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__S1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ net1807 _01754_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[608\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_15_0_clk_X clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187__839 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__inv_2
X_12046_ net1738 _01685_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[539\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09156__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08364__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12492__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07014__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09630__A _02532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06773__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06525__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload112 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__clkinv_16
XANTENNA__07642__A2 _03463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload101 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_8
X_08070_ net209 net690 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__and2_1
X_07021_ top0.CPU.register.registers\[287\] top0.CPU.register.registers\[319\] top0.CPU.register.registers\[351\]
+ top0.CPU.register.registers\[383\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__mux4_1
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload123 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__clkinv_8
X_10795__447 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__inv_2
XANTENNA__07296__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ top0.CPU.register.registers\[181\] net568 vssd1 vssd1 vccd1 vccd1 _04787_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09147__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ top0.CPU.intMem_out\[16\] net625 _02813_ _02386_ net638 vssd1 vssd1 vccd1
+ vccd1 _04565_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_71_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836__488 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__inv_2
Xhold18 top0.CPU.register.registers\[4\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 top0.CPU.register.registers\[22\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07854_ _04388_ net231 net226 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__and3_1
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06805_ _03458_ _03461_ net867 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
XFILLER_56_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout364_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ net342 _04433_ _04434_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a31o_1
X_10689__341 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__inv_2
X_09524_ top0.CPU.Op\[2\] _05071_ net127 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XANTENNA__08855__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06736_ net871 _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and2_1
XFILLER_25_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09455_ top0.MMIO.WBData_i\[21\] net147 _05037_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__o21a_1
XFILLER_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06667_ top0.CPU.register.registers\[513\] top0.CPU.register.registers\[545\] top0.CPU.register.registers\[577\]
+ top0.CPU.register.registers\[609\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03324_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06764__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ net195 net697 net403 net379 net2674 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a32o_1
XANTENNA__07330__A1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09386_ net2558 _04475_ net606 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__mux2_1
X_06598_ _03251_ _03252_ _03253_ _03254_ net757 net749 vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07881__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08337_ net719 net201 net399 net411 net2328 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07995__A _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ net2912 net417 _04718_ net494 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
X_07219_ _03721_ _03724_ net455 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__mux2_1
X_10230_ net33 net653 net592 top0.MMIO.WBData_i\[9\] vssd1 vssd1 vccd1 vccd1 _02276_
+ sky130_fd_sc_hd__o22a_1
X_08199_ net3266 net421 _04692_ net499 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a22o_1
XANTENNA__08603__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__A3 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _02952_ _02960_ net551 vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__o21ba_1
XFILLER_126_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1027 net1029 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_4
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
Xfanout1005 net1007 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
Xfanout1038 net1041 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
X_10092_ top0.display.delayctr\[13\] _05562_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09138__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08346__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08897__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06109__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07857__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06755__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07321__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12664_ clknet_leaf_93_clk _02299_ net1081 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ net1307 _01254_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_12595_ clknet_leaf_90_clk _02230_ net1079 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ net1238 _01185_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10482__134 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__inv_2
XANTENNA__06832__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ clknet_leaf_80_clk top0.CPU.internalMem.state_n\[2\] net1111 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.state\[2\] sky130_fd_sc_hd__dfrtp_1
X_10523__175 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__inv_2
XFILLER_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10396__48 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09129__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06060__B2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ net1721 _01668_ net1029 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[522\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08337__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08352__A3 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ net462 _04225_ _04226_ _04170_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__o22a_1
X_06521_ top0.CPU.register.registers\[658\] top0.CPU.register.registers\[690\] top0.CPU.register.registers\[722\]
+ top0.CPU.register.registers\[754\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08104__A3 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ top0.CPU.intMemAddr\[4\] _04616_ net769 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__mux2_1
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06195__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06452_ top0.CPU.register.registers\[22\] top0.CPU.register.registers\[54\] top0.CPU.register.registers\[86\]
+ top0.CPU.register.registers\[118\] net923 net889 vssd1 vssd1 vccd1 vccd1 _03109_
+ sky130_fd_sc_hd__mux4_1
X_09171_ net186 net672 net276 net249 net2613 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a32o_1
X_06383_ net544 _02984_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nor2_1
X_08122_ net2821 _04555_ net431 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
XANTENNA__07076__A0 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05887__X _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ net509 net169 net709 net438 net2411 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a32o_1
X_07004_ _03657_ _03660_ _03638_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o21bai_2
XANTENNA_fanout112_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1021_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08040__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08955_ net163 net702 net270 net264 net2363 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__a32o_1
X_07906_ _02391_ _04549_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout579_A _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A _02575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08328__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ top0.CPU.register.registers\[243\] net575 vssd1 vssd1 vccd1 vccd1 _04763_
+ sky130_fd_sc_hd__or2_1
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06230__Y _02887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ top0.CPU.internalMem.pcOut\[29\] net641 net635 _04491_ vssd1 vssd1 vccd1
+ vccd1 _04492_ sky130_fd_sc_hd__o211a_2
XFILLER_57_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _02869_ _03129_ net340 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__a21o_1
XANTENNA__05788__S1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ top0.MMIO.WBData_i\[5\] net148 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09270__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06719_ top0.CPU.register.registers\[260\] top0.CPU.register.registers\[292\] top0.CPU.register.registers\[324\]
+ top0.CPU.register.registers\[356\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03376_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08500__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ _03796_ _03933_ _03947_ _03824_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout913_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09438_ top0.MMIO.WBData_i\[15\] net145 _05028_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__o21a_1
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ net2504 _04573_ net607 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
X_10466__118 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__inv_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300__952 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__inv_2
X_12380_ net2072 _02019_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[873\]
+ sky130_fd_sc_hd__dfrtp_1
X_11400_ clknet_leaf_59_clk _01048_ net1091 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07067__A0 _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10507__159 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__inv_2
XFILLER_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10213_ net2574 net117 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__and2_1
XANTENNA__08031__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10144_ net3385 net663 net661 _05603_ _05606_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a221o_1
XANTENNA__06788__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10075_ _05551_ _05552_ net601 vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05779__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06976__S0 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_26_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_12647_ clknet_leaf_65_clk _02282_ net1102 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05856__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09047__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043__695 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__inv_2
X_12578_ clknet_leaf_90_clk _02213_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08243__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold307 top0.CPU.register.registers\[229\] vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
X_11529_ net1221 _01168_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold318 top0.CPU.register.registers\[560\] vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 top0.CPU.register.registers\[612\] vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 net819 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_2
Xhold1018 top0.CPU.register.registers\[670\] vssd1 vssd1 vccd1 vccd1 net3240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1007 top0.CPU.register.registers\[61\] vssd1 vssd1 vccd1 vccd1 net3229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 top0.CPU.register.registers\[952\] vssd1 vssd1 vccd1 vccd1 net3251 sky130_fd_sc_hd__dlygate4sd3_1
X_08740_ _04682_ net315 net294 net2705 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__a22o_1
X_05952_ top0.CPU.register.registers\[385\] top0.CPU.register.registers\[417\] top0.CPU.register.registers\[449\]
+ top0.CPU.register.registers\[481\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02609_
+ sky130_fd_sc_hd__mux4_1
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08671_ _04663_ net315 net298 net2997 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a22o_1
X_05883_ top0.CPU.register.registers\[771\] top0.CPU.register.registers\[803\] top0.CPU.register.registers\[835\]
+ top0.CPU.register.registers\[867\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02540_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08730__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07622_ _03340_ _03358_ _03357_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06967__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ _02457_ _03092_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__and2b_1
XANTENNA__06719__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06504_ top0.CPU.register.registers\[787\] top0.CPU.register.registers\[819\] top0.CPU.register.registers\[851\]
+ top0.CPU.register.registers\[883\] net940 net906 vssd1 vssd1 vccd1 vccd1 _03161_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_66_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07484_ _02888_ _03112_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__nand2_1
XANTENNA__07297__B1 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09223_ top0.CPU.internalMem.pcOut\[26\] top0.CPU.internalMem.pcOut\[25\] top0.CPU.internalMem.pcOut\[24\]
+ top0.CPU.internalMem.pcOut\[23\] vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__or4_1
X_06435_ net745 _03091_ _03082_ _03086_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ _04712_ net268 net247 net2787 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a22o_1
XANTENNA__05942__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06366_ _03007_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__xnor2_1
X_08105_ net493 net159 net690 net433 net2424 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_4_3_0_clk_X clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout115_X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ net171 net616 net271 net255 net2445 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__a32o_1
X_06297_ top0.CPU.register.registers\[411\] top0.CPU.register.registers\[443\] top0.CPU.register.registers\[475\]
+ top0.CPU.register.registers\[507\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02954_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08153__B net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08261__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ net637 _04548_ net710 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__and3_2
XANTENNA__12595__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold830 top0.CPU.register.registers\[142\] vssd1 vssd1 vccd1 vccd1 net3052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold863 top0.CPU.register.registers\[852\] vssd1 vssd1 vccd1 vccd1 net3085 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 top0.CPU.register.registers\[566\] vssd1 vssd1 vccd1 vccd1 net3074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 top0.CPU.register.registers\[792\] vssd1 vssd1 vccd1 vccd1 net3063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09265__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05793__A top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 net81 vssd1 vssd1 vccd1 vccd1 net3096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 top0.CPU.register.registers\[950\] vssd1 vssd1 vccd1 vccd1 net3118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 top0.CPU.register.registers\[157\] vssd1 vssd1 vccd1 vccd1 net3107 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ _05475_ _05476_ _05477_ net235 net645 vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__o221ai_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851__503 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__inv_2
X_08938_ net196 net709 net278 net265 net2514 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ net3370 net284 _04756_ _04488_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06958__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ net1572 _01519_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[373\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05957__A1_N net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11027__679 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__inv_2
XANTENNA__11406__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05838__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06186__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12501_ net2193 _02140_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[994\]
+ sky130_fd_sc_hd__dfrtp_1
X_12432_ net2124 _02071_ net1081 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[925\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08788__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06416__X _03073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_97_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08252__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12363_ net2055 _02002_ net1072 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[856\]
+ sky130_fd_sc_hd__dfrtp_1
X_12294_ net1986 _01933_ net1128 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366__18 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__inv_2
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08004__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594__246 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08960__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05591_ _05592_ net600 vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__a21oi_1
X_10058_ top0.display.delayctr\[4\] _05536_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08712__A0 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10635__287 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__inv_2
XFILLER_63_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10488__140 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__inv_2
XANTENNA__06981__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08491__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06220_ _02875_ _02876_ net786 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
XANTENNA__05924__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10529__181 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__inv_2
XANTENNA__08779__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06151_ _02804_ _02807_ net777 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
X_06082_ _02735_ _02736_ _02737_ _02738_ net729 net738 vssd1 vssd1 vccd1 vccd1 _02739_
+ sky130_fd_sc_hd__mux4_2
Xhold104 top0.CPU.register.registers\[969\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 top0.CPU.register.registers\[754\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold115 top0.CPU.register.registers\[992\] vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 top0.CPU.register.registers\[748\] vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ net239 _05404_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__o21ai_1
Xhold148 top0.CPU.register.registers\[976\] vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 top0.CPU.register.registers\[611\] vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout606 net612 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload14_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ _02813_ _04563_ net587 vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__mux2_1
Xfanout639 _02383_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_2
Xfanout628 _02419_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08546__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_4
XANTENNA__08951__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08420__C net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ top0.CPU.internalMem.pcOut\[10\] net650 _05279_ vssd1 vssd1 vccd1 vccd1 _02187_
+ sky130_fd_sc_hd__o21a_1
XFILLER_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06984_ top0.CPU.register.registers\[666\] top0.CPU.register.registers\[698\] top0.CPU.register.registers\[730\]
+ top0.CPU.register.registers\[762\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03641_
+ sky130_fd_sc_hd__mux4_1
X_08723_ net168 net3220 net359 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__mux2_1
X_05935_ top0.CPU.register.registers\[128\] top0.CPU.register.registers\[160\] top0.CPU.register.registers\[192\]
+ top0.CPU.register.registers\[224\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02592_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout277_A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380__32 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08703__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ net167 net708 net322 net303 net2627 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a32o_1
X_05866_ top0.CPU.register.registers\[779\] top0.CPU.register.registers\[811\] top0.CPU.register.registers\[843\]
+ top0.CPU.register.registers\[875\] net844 net809 vssd1 vssd1 vccd1 vccd1 _02523_
+ sky130_fd_sc_hd__mux4_1
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09024__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05797_ _02447_ _02449_ _02452_ _02341_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a31oi_4
XANTENNA_fanout444_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ _04223_ _04225_ net458 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
X_08585_ net2790 net166 net333 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07052__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ _04187_ _04188_ _04192_ _04154_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__o31a_1
XANTENNA__08863__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout709_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ _04530_ _04546_ _04552_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__or3_1
XANTENNA__08482__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07467_ _02650_ net532 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06418_ _03059_ net538 vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__and2_1
X_07398_ net441 _04049_ _04050_ _04054_ _04048_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__o221a_1
XANTENNA__06493__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06349_ _02984_ _03005_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__nand2_1
X_09137_ top0.CPU.register.registers\[68\] net565 net213 net680 net553 vssd1 vssd1
+ vccd1 vccd1 _04839_ sky130_fd_sc_hd__o2111a_1
X_09068_ top0.CPU.register.registers\[114\] net571 net560 vssd1 vssd1 vccd1 vccd1
+ _04816_ sky130_fd_sc_hd__o21a_1
XANTENNA__08785__A3 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ net3246 net437 _04640_ net499 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a22o_1
Xhold660 top0.CPU.register.registers\[653\] vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 top0.CPU.register.registers\[494\] vssd1 vssd1 vccd1 vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 top0.CPU.register.registers\[901\] vssd1 vssd1 vccd1 vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08537__A3 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold682 top0.CPU.register.registers\[861\] vssd1 vssd1 vccd1 vccd1 net2904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08942__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05851__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06131__B _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ net1624 _01571_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[425\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06558__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ net1555 _01502_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11794_ net1486 _01433_ net1053 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08473__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05906__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08074__A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12415_ net2107 _02054_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[908\]
+ sky130_fd_sc_hd__dfrtp_1
X_12346_ net2038 _01985_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07433__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__A _02809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__B _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ net1969 _01916_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[770\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07418__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06322__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06095__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05842__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11399__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05720_ top0.CPU.Op\[0\] top0.CPU.Op\[1\] top0.CPU.Op\[2\] vssd1 vssd1 vccd1 vccd1
+ _02377_ sky130_fd_sc_hd__and3_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07153__A _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ net199 net707 net399 net383 net2357 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a32o_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_63_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ net527 net526 net469 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__mux2_1
XFILLER_118_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ _03808_ _03821_ net464 vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_1
XANTENNA__06570__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06203_ net783 _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__and2_1
X_07183_ net453 _03743_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__nor2_1
X_06134_ _02514_ _02790_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__and2_1
XANTENNA__07975__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06065_ top0.CPU.register.registers\[522\] top0.CPU.register.registers\[554\] top0.CPU.register.registers\[586\]
+ top0.CPU.register.registers\[618\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02722_
+ sky130_fd_sc_hd__mux4_1
XFILLER_132_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout403 net406 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09177__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 _04720_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09019__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08519__A3 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _04653_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_8
X_09824_ net648 _05327_ _05316_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06086__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout425 _04672_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_8
X_11249__901 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__inv_2
XANTENNA__08924__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 _03150_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08858__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 net461 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
Xfanout469 _02598_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
X_09755_ _05250_ _05252_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout561_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06967_ top0.CPU.register.registers\[667\] top0.CPU.register.registers\[699\] top0.CPU.register.registers\[731\]
+ top0.CPU.register.registers\[763\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03624_
+ sky130_fd_sc_hd__mux4_1
X_06898_ _03551_ _03552_ _03554_ _03553_ net871 net751 vssd1 vssd1 vccd1 vccd1 _03555_
+ sky130_fd_sc_hd__mux4_2
X_09686_ _05197_ _05198_ top0.CPU.internalMem.pcOut\[4\] vssd1 vssd1 vccd1 vccd1 _05200_
+ sky130_fd_sc_hd__a21o_1
X_05918_ _02573_ _02574_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__and2_1
X_08706_ net204 net3276 net358 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
XFILLER_27_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05849_ top0.CPU.register.registers\[143\] top0.CPU.register.registers\[175\] top0.CPU.register.registers\[207\]
+ top0.CPU.register.registers\[239\] net851 net816 vssd1 vssd1 vccd1 vccd1 _02506_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08152__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08637_ net705 _04739_ net302 net2611 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a22o_1
XANTENNA__06389__S1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963__615 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__inv_2
XFILLER_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout826_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ net3092 _04544_ net335 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XANTENNA__05910__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09101__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ _04700_ net400 net367 net2610 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__a22o_1
X_07519_ net455 _03810_ _03338_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__a21o_1
XANTENNA__05789__Y _02446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06561__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08207__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ net1892 _01839_ net1077 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[693\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08758__A3 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net1823 _01770_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[624\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net1754 _01701_ net1007 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold490 top0.CPU.register.registers\[91\] vssd1 vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07238__A _02578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07718__A1 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout970 net976 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07194__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05824__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
Xfanout992 net995 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1190 top0.CPU.intMem_out\[16\] vssd1 vssd1 vccd1 vccd1 net3412 sky130_fd_sc_hd__dlygate4sd3_1
X_11915_ net1607 _01554_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ net1538 _01485_ net1122 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09643__A1 _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11_0_clk_X clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11777_ net1469 _01416_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08915__C_N net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10747__399 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06552__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload13 clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_8
Xclkload24 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinv_8
Xclkload35 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_11_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload57 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_16
Xclkload68 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_4
XANTENNA__06604__X _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_6
Xclkload79 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__inv_4
X_12329_ net2021 _01968_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06090__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09159__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08251__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06068__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08906__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _02386_ _02907_ _04476_ _04518_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08382__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06987__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650__302 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__inv_2
X_06821_ top0.CPU.register.registers\[397\] top0.CPU.register.registers\[429\] top0.CPU.register.registers\[461\]
+ top0.CPU.register.registers\[493\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03478_
+ sky130_fd_sc_hd__mux4_1
X_09540_ net867 _05083_ net127 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
X_06752_ _03364_ _03383_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__a21oi_2
X_09471_ top0.MMIO.WBData_i\[29\] _05041_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and2_1
X_05703_ net1 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__inv_2
XFILLER_64_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08422_ net3149 _04481_ net375 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__mux2_1
XANTENNA__08685__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06683_ _03321_ _03322_ _03338_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_19_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06791__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ net717 net153 net394 net410 net2450 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a32o_1
X_07304_ _03720_ _03957_ _03960_ net441 _03959_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o221a_1
X_08284_ net497 net161 net668 net418 net2653 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a32o_1
X_07235_ _03799_ _03802_ net457 vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__mux2_1
Xclkload7 clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_8
XANTENNA_fanout407_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07166_ _03821_ _03822_ net464 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06117_ top0.CPU.register.registers\[654\] top0.CPU.register.registers\[686\] top0.CPU.register.registers\[718\]
+ top0.CPU.register.registers\[750\] net835 net801 vssd1 vssd1 vccd1 vccd1 _02774_
+ sky130_fd_sc_hd__mux4_1
X_07097_ net518 net457 net474 vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or3b_2
X_06048_ net784 _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__and2_1
XANTENNA__07058__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08161__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout776_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 _04498_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
Xfanout222 _04561_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06908__C1 _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_4
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
XANTENNA__08588__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _04772_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout288 _04750_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_4
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_8
X_09807_ _05309_ _05310_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout943_A top0.CPU.control.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07999_ net713 net497 net161 net546 net2296 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ top0.CPU.control.funct7\[3\] _02453_ net590 vssd1 vssd1 vccd1 vccd1 _05248_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__06923__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__B _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _05181_ _05183_ net237 vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__o21a_1
XANTENNA__08676__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06836__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ clknet_leaf_82_clk _02315_ net1108 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
X_11700_ net1392 _01339_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09625__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11631_ net1323 _01270_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06782__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07240__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ net1254 _01201_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ clknet_leaf_90_clk _01132_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire678 _04704_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_2
XANTENNA__06571__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08061__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12114_ net1806 _01753_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[607\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07403__A3 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12045_ net1737 _01684_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[538\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06470__S0 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__B _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11829_ net1521 _01468_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08419__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10226__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06525__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload113 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__clkinv_16
XFILLER_119_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload102 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__inv_12
X_07020_ net865 _03672_ _03675_ _03676_ net861 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__o221a_1
Xclkload124 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__inv_6
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08052__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170__822 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08971_ _04662_ net555 _04786_ net262 net3309 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__a32o_1
X_07922_ net561 _04563_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold19 top0.display.delayctr\[31\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
X_11211__863 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__inv_2
XANTENNA__09552__A0 top0.CPU.control.funct7\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07853_ net3033 net546 net494 _04505_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06804_ _03459_ _03460_ net766 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07784_ net451 _04289_ _04435_ _03848_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a221o_1
X_09523_ top0.CPU.Op\[1\] _05060_ net127 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
X_06735_ top0.CPU.register.registers\[902\] top0.CPU.register.registers\[934\] top0.CPU.register.registers\[966\]
+ top0.CPU.register.registers\[998\] net929 net895 vssd1 vssd1 vccd1 vccd1 _03392_
+ sky130_fd_sc_hd__mux4_1
XFILLER_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08658__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ net130 net133 _05045_ net597 net3376 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06666_ top0.CPU.register.registers\[641\] top0.CPU.register.registers\[673\] top0.CPU.register.registers\[705\]
+ top0.CPU.register.registers\[737\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03323_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_35_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06764__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ net2455 _04483_ net612 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__mux2_1
X_08405_ _04667_ net394 net378 net2580 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout524_A _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06597_ top0.CPU.register.registers\[519\] top0.CPU.register.registers\[551\] top0.CPU.register.registers\[583\]
+ top0.CPU.register.registers\[615\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03254_
+ sky130_fd_sc_hd__mux4_1
X_08336_ net3169 net409 net389 _04562_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
XANTENNA__09083__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ net222 net670 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__and2_1
XANTENNA__08830__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06841__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08198_ net211 net681 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__and2_1
X_07218_ net486 _03760_ _03865_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o31a_1
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout893_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ net347 _03756_ _03789_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__o31ai_1
XFILLER_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__B2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ net3431 net663 net661 _05616_ _05619_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
Xfanout1017 net1018 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_2
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
X_10091_ net3393 net665 net603 _05564_ _05163_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a221o_1
Xfanout1039 net1040 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08346__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08111__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10969__621 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08649__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06755__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ clknet_leaf_66_clk _02298_ net1119 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08066__B net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11614_ net1306 _01253_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_12594_ clknet_leaf_89_clk _02229_ net1079 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09074__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11545_ net1237 _01184_ net980 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08282__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05977__Y _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_131_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11476_ clknet_leaf_76_clk top0.CPU.internalMem.state_n\[1\] net1124 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.state\[1\] sky130_fd_sc_hd__dfrtp_1
X_11154__806 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06380__A1_N net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10289_ net3044 net120 net113 _05665_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__A0 top0.CPU.control.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ net1720 _01667_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08337__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08888__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048__700 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__inv_2
XANTENNA__06899__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09641__A _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06520_ _03157_ net535 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__xnor2_1
X_06451_ top0.CPU.register.registers\[150\] top0.CPU.register.registers\[182\] top0.CPU.register.registers\[214\]
+ top0.CPU.register.registers\[246\] net923 net889 vssd1 vssd1 vccd1 vccd1 _03108_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10762__414 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__inv_2
X_09170_ net191 net677 net280 net250 net2291 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__a32o_1
XANTENNA__09065__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06382_ _03023_ net539 vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__xor2_1
XANTENNA__08273__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08121_ net2848 _04548_ net432 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
XANTENNA__07076__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_122_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10803__455 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__inv_2
X_08052_ net504 net173 net706 net438 net2522 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a32o_1
XANTENNA__10080__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08812__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ _03623_ net521 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__nor2_1
XANTENNA__06999__X _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08954_ net164 net703 net270 net264 net2603 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09027__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__inv_2
XANTENNA__09525__A0 top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ _04545_ net554 _04762_ net282 net3137 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__a32o_1
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08879__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ _04476_ _04489_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a21o_1
XFILLER_56_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06434__S0 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net245 _04242_ _04423_ net448 vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__a22o_1
XANTENNA__06985__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _02358_ net138 vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout739_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06718_ top0.CPU.register.registers\[388\] top0.CPU.register.registers\[420\] top0.CPU.register.registers\[452\]
+ top0.CPU.register.registers\[484\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03375_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07839__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07698_ _03154_ _03914_ _03579_ _03115_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o211ai_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09437_ net3443 net597 net130 _05034_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06649_ top0.CPU.register.registers\[642\] top0.CPU.register.registers\[674\] top0.CPU.register.registers\[706\]
+ top0.CPU.register.registers\[738\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03306_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08454__X _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ net2716 _04578_ net607 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09056__A2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09299_ top0.CPU.addrControl _04951_ _04952_ vssd1 vssd1 vccd1 vccd1 top0.display.next_state\[0\]
+ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_113_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08319_ net2903 net154 net413 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08803__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546__198 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__inv_2
XANTENNA__08567__A1 _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ net2781 net123 net116 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a21o_1
XANTENNA__09285__X _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ _05604_ _05605_ net600 vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10074_ top0.display.delayctr\[8\] _05548_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09461__A top0.MMIO.WBData_i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06976__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08098__A3 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12646_ clknet_leaf_71_clk _02281_ net1119 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09047__A2 _04797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_104_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12577_ clknet_leaf_90_clk _02212_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold308 top0.CPU.register.registers\[428\] vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08270__A3 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11528_ net1220 _01167_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11459_ clknet_leaf_65_clk _01107_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold319 top0.CPU.register.registers\[56\] vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09636__A _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06018__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1019 top0.CPU.register.registers\[647\] vssd1 vssd1 vccd1 vccd1 net3241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1008 top0.CPU.register.registers\[857\] vssd1 vssd1 vccd1 vccd1 net3230 sky130_fd_sc_hd__dlygate4sd3_1
X_05951_ _02606_ _02607_ net724 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
XFILLER_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282__934 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__inv_2
X_08670_ net693 _04739_ net298 net2780 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a22o_1
X_05882_ _02537_ _02538_ net726 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
XANTENNA__08730__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07621_ _02578_ net245 _03877_ _04172_ net441 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__o32a_1
XANTENNA__06967__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07552_ _04206_ _04207_ _04208_ _04146_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o31a_1
X_06503_ _03158_ _03159_ net766 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__mux2_1
X_11323__975 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__inv_2
XANTENNA__08089__A3 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06719__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09140__D1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07483_ _02888_ net536 vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08494__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ net770 _04873_ _04876_ _04879_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a221o_1
XANTENNA__09038__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06434_ _03087_ _03088_ _03090_ _03089_ net869 net749 vssd1 vssd1 vccd1 vccd1 _03091_
+ sky130_fd_sc_hd__mux4_1
X_06365_ net583 _02454_ _03008_ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__o31a_2
X_09153_ _04711_ net267 net247 net2883 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a22o_1
XFILLER_108_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ net497 net162 net690 net433 net2488 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout222_A _04561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ net175 net615 net276 net257 net2487 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__a32o_1
X_06296_ top0.CPU.register.registers\[283\] top0.CPU.register.registers\[315\] top0.CPU.register.registers\[347\]
+ top0.CPU.register.registers\[379\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02953_
+ sky130_fd_sc_hd__mux4_1
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1131_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08035_ net3166 net439 _04648_ net498 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a22o_1
Xhold820 top0.CPU.register.registers\[279\] vssd1 vssd1 vccd1 vccd1 net3042 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 top0.CPU.register.registers\[158\] vssd1 vssd1 vccd1 vccd1 net3053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 top0.CPU.register.registers\[759\] vssd1 vssd1 vccd1 vccd1 net3075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 top0.CPU.register.registers\[398\] vssd1 vssd1 vccd1 vccd1 net3064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 top0.CPU.register.registers\[533\] vssd1 vssd1 vccd1 vccd1 net3086 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A3 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 net65 vssd1 vssd1 vccd1 vccd1 net3097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold897 top0.CPU.register.registers\[846\] vssd1 vssd1 vccd1 vccd1 net3119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 top0.CPU.register.registers\[440\] vssd1 vssd1 vccd1 vccd1 net3108 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ top0.CPU.internalMem.pcOut\[27\] _05467_ vssd1 vssd1 vccd1 vccd1 _05477_
+ sky130_fd_sc_hd__xnor2_1
X_10890__542 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__inv_2
XANTENNA_fanout856_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ net200 net707 _04778_ net265 net3324 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ top0.CPU.register.registers\[254\] _02396_ net559 vssd1 vssd1 vccd1 vccd1
+ _04756_ sky130_fd_sc_hd__o21a_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06407__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10931__583 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__inv_2
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _02387_ top0.CPU.Op\[4\] _02386_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__and3b_2
XANTENNA__06958__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ _04707_ net324 net287 net2896 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10220__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__D1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07513__B _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08485__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12500_ net2192 _02139_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[993\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ net2123 _02070_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[924\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08237__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12362_ net2054 _02001_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06894__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ net1985 _01932_ net1038 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05774__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ top0.display.delayctr\[20\] _05587_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__nand2_1
X_11266__918 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__inv_2
X_10057_ top0.display.delayctr\[4\] _05536_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11010__662 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__inv_2
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11307__959 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__inv_2
XANTENNA_clkload0_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08476__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07279__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ clknet_leaf_75_clk _02264_ net1124 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08228__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09440__A2 _05006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06150_ _02805_ _02806_ net726 vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
X_06081_ top0.CPU.register.registers\[525\] top0.CPU.register.registers\[557\] top0.CPU.register.registers\[589\]
+ top0.CPU.register.registers\[621\] net850 net815 vssd1 vssd1 vccd1 vccd1 _02738_
+ sky130_fd_sc_hd__mux4_1
Xhold116 top0.CPU.register.registers\[937\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07987__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 top0.CPU.register.registers\[578\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
X_10874__526 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__inv_2
Xhold127 top0.CPU.register.registers\[1005\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold138 top0.CPU.register.registers\[370\] vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 top0.CPU.intMemAddr\[19\] vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05894__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout607 net612 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
X_09840_ _05338_ _05341_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__nand2_1
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
Xfanout618 _04670_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06637__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ _05276_ _05277_ _05278_ net241 net652 vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__a221o_1
X_06983_ _02944_ _03639_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__xnor2_1
X_10915__567 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__inv_2
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08722_ net172 net3051 net357 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__mux2_1
X_05934_ net786 _02588_ net780 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_68_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05865_ net778 _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ net171 net703 net312 net302 net2700 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout172_A _04611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05796_ _02447_ _02449_ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__nand3_2
X_08584_ net2838 net215 net333 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__mux2_1
XFILLER_54_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__10161__B1_N net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768__420 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__inv_2
X_07604_ net482 _03996_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__and2_1
XANTENNA__08467__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07535_ _04165_ _04184_ _04191_ _04163_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__a2bb2o_1
X_07466_ _04115_ _04122_ _04118_ _04050_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout437_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09040__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ top0.CPU.intMemAddr\[19\] top0.CPU.intMemAddr\[18\] top0.CPU.intMemAddr\[17\]
+ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__or4_1
X_10809__461 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__inv_2
X_06417_ _03059_ net538 vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__nor2_1
XANTENNA__08482__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ _04012_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09136_ net167 net685 _04838_ net253 net3329 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__a32o_1
X_06348_ net580 _02455_ _03002_ _03004_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a31o_2
XANTENNA__08234__A3 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ _04684_ net560 _04815_ net258 net3001 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__a32o_1
XANTENNA__06876__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06279_ net776 _02931_ _02934_ _02935_ net772 vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__o221a_1
XANTENNA__09276__A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08018_ net211 net701 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__and2_1
Xhold650 net52 vssd1 vssd1 vccd1 vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 top0.CPU.register.registers\[1012\] vssd1 vssd1 vccd1 vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 top0.CPU.register.registers\[58\] vssd1 vssd1 vccd1 vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold694 top0.CPU.register.registers\[660\] vssd1 vssd1 vccd1 vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 top0.CPU.register.registers\[1021\] vssd1 vssd1 vccd1 vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__inv_2
XFILLER_92_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05851__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07524__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11931_ net1623 _01570_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[424\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_28_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06800__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11862_ net1554 _01501_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[355\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08458__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net1485 _01432_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[286\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08473__A3 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06574__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07130__A0 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07681__A1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08074__B net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10426__78 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__inv_2
X_10561__213 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__inv_2
X_12414_ net2106 _02053_ net1013 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[907\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08225__A3 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12345_ net2037 _01984_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07984__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10602__254 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__inv_2
X_12276_ net1968 _01915_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06619__S0 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__B _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06322__B _02978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06095__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09914__A top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ _02809_ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nor2_1
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05842__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08697__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07153__B _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08249__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07320_ net528 _03482_ net469 vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__mux2_1
XANTENNA__06484__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__A_N net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07251_ _03817_ _03822_ net455 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__mux2_1
XANTENNA__09648__X _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06202_ top0.CPU.register.registers\[916\] top0.CPU.register.registers\[948\] top0.CPU.register.registers\[980\]
+ top0.CPU.register.registers\[1012\] net833 net798 vssd1 vssd1 vccd1 vccd1 _02859_
+ sky130_fd_sc_hd__mux4_1
X_07182_ net452 _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__or2_1
XANTENNA__09413__A2 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06133_ _02788_ _02789_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__and2_2
XANTENNA__08621__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07975__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06072__X _02729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06064_ top0.CPU.register.registers\[650\] top0.CPU.register.registers\[682\] top0.CPU.register.registers\[714\]
+ top0.CPU.register.registers\[746\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02721_
+ sky130_fd_sc_hd__mux4_1
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
XFILLER_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440__92 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__inv_2
X_11288__940 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__inv_2
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
X_09823_ net235 _05325_ _05326_ _05323_ _05324_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__o32a_1
XANTENNA__06086__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07727__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout448 _02636_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout437 net439 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_4
Xfanout426 _04672_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10192__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout459 net461 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06935__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329__981 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__inv_2
X_09754_ _05260_ _05261_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__and2_1
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06966_ _02962_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06659__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ top0.CPU.internalMem.pcOut\[4\] _05197_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_
+ sky130_fd_sc_hd__and3_1
X_06897_ top0.CPU.register.registers\[8\] top0.CPU.register.registers\[40\] top0.CPU.register.registers\[72\]
+ top0.CPU.register.registers\[104\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03554_
+ sky130_fd_sc_hd__mux4_1
X_05917_ _02556_ _02557_ net583 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout554_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07344__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ net205 net3037 net358 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05848_ net778 _02500_ _02504_ net773 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__o211a_2
XANTENNA__07063__B _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08152__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08159__B net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08636_ _04645_ net305 net301 net2879 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a22o_1
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout819_A top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05910__A1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05779_ top0.CPU.register.registers\[791\] top0.CPU.register.registers\[823\] top0.CPU.register.registers\[855\]
+ top0.CPU.register.registers\[887\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02436_
+ sky130_fd_sc_hd__mux4_1
X_08567_ net3086 _04539_ net334 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
X_07518_ _04154_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__nand2_2
X_08498_ _04699_ net396 net366 net2817 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a22o_1
X_07449_ _04089_ _04090_ _04105_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__o21ai_4
XANTENNA__08860__A0 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ net196 net686 net278 net253 net2407 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_94_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08612__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12130_ net1822 _01769_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[623\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07966__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05977__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ net1753 _01700_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[554\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold480 top0.CPU.register.registers\[561\] vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 net47 vssd1 vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06926__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 net962 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08391__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05824__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout982 net1004 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout971 net976 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08679__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1191 top0.MMIO.WBData_i\[7\] vssd1 vssd1 vccd1 vccd1 net3413 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_84_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 top0.display.delayctr\[4\] vssd1 vssd1 vccd1 vccd1 net3402 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ net1606 _01553_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[407\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11081__733 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ net1537 _01484_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ net1468 _01415_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09643__A2 _02511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__B _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122__774 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__inv_2
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload14 clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload25 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_11_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload58 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_12
Xclkload69 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_12
Xclkload47 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__inv_2
Xclkload36 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_12
X_12328_ net2020 _01967_ net1077 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06333__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12259_ net1951 _01898_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[752\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06068__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ net864 _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__nor2_1
XFILLER_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07017__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ _03386_ _03405_ _03263_ _03384_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a211o_1
X_10986__638 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__inv_2
X_09470_ net130 net133 _05053_ net597 net3421 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_75_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
X_05702_ net3390 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__inv_2
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06682_ _03321_ _03322_ _03338_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__a21oi_1
X_08421_ net545 _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor2_1
X_10730__382 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__inv_2
XANTENNA__07342__A0 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__A2 _05162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06009__A1_N _02665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08352_ net713 net157 net386 net409 net2312 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a32o_1
X_07303_ _02477_ _03173_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07645__A1 _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ net495 net166 net670 net417 net2581 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a32o_1
X_07234_ _03791_ _03801_ net465 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__mux2_1
Xclkload8 clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_12
XANTENNA__06942__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1044_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout302_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07165_ net525 _03519_ net472 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__mux2_1
XANTENNA__07948__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06116_ _02473_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07096_ _03704_ net443 _03750_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05959__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06047_ top0.CPU.register.registers\[904\] top0.CPU.register.registers\[936\] top0.CPU.register.registers\[968\]
+ top0.CPU.register.registers\[1000\] net844 net809 vssd1 vssd1 vccd1 vccd1 _02704_
+ sky130_fd_sc_hd__mux4_1
Xfanout212 _04487_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout201 _04567_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout223 _04544_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _04471_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
Xfanout245 _03774_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
Xfanout256 _04809_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout671_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _05309_ _05310_ net236 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__o21a_1
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
X_07998_ net768 net640 net635 _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__o211a_2
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_8
Xfanout267 net269 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09737_ _04069_ net232 net227 net631 vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a31o_1
X_06949_ _03604_ _03605_ net764 vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065__717 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__inv_2
XFILLER_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09873__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ _05181_ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__nand2_1
XANTENNA__07802__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ net3354 net604 net658 net3358 _05137_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__a221o_1
X_08619_ net714 net175 net310 net329 net2636 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08109__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106__758 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__inv_2
XANTENNA__07550__A_N _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05895__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ net1322 _01269_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08833__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05990__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ net1253 _01200_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ clknet_leaf_90_clk _01131_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06153__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12113_ net1805 _01752_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[606\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673__325 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__inv_2
X_12044_ net1736 _01683_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[537\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09010__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout790 net799 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_2
X_10714__366 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_57_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06470__S1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_47_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__A0 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09077__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ net1520 _01467_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05886__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05981__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09616__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__A3 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08824__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ net1451 _01398_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[252\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload103 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__inv_6
XANTENNA__09639__A _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608__260 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__inv_2
Xclkload114 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__clkinv_16
Xclkload125 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__clkinv_16
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08052__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410__62 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__inv_2
X_08970_ top0.CPU.register.registers\[182\] net568 vssd1 vssd1 vccd1 vccd1 _04786_
+ sky130_fd_sc_hd__or2_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07921_ _04317_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__and3_1
XFILLER_69_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__09001__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08355__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07852_ net717 net210 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__and2_1
X_06803_ top0.CPU.register.registers\[268\] top0.CPU.register.registers\[300\] top0.CPU.register.registers\[332\]
+ top0.CPU.register.registers\[364\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03460_
+ sky130_fd_sc_hd__mux4_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
X_09522_ top0.CPU.Op\[0\] _05064_ net127 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
X_07783_ _04436_ _04437_ _04438_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__nand4_1
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06734_ top0.CPU.register.registers\[774\] top0.CPU.register.registers\[806\] top0.CPU.register.registers\[838\]
+ top0.CPU.register.registers\[870\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03391_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08658__A3 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ top0.MMIO.WBData_i\[20\] _05041_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__and2_1
X_06665_ net542 net471 net463 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout252_A _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08404_ net197 net697 net404 net379 net2351 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a32o_1
XANTENNA__09068__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ net2559 _04489_ net606 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__mux2_1
XANTENNA__05877__B1 top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08335_ net719 net203 net400 net411 net2348 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a32o_1
X_06596_ top0.CPU.register.registers\[647\] top0.CPU.register.registers\[679\] top0.CPU.register.registers\[711\]
+ top0.CPU.register.registers\[743\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03253_
+ sky130_fd_sc_hd__mux4_1
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07618__A1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05972__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ net508 net203 net673 net419 net2414 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a32o_1
XANTENNA__08291__A1 _04498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ net2904 net422 _04691_ net503 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08830__A3 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07217_ net477 _03866_ _03867_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a31o_1
X_07148_ _02555_ _03796_ _03800_ _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a211o_1
XANTENNA__08594__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout886_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657__309 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__inv_2
XFILLER_105_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ _03728_ _03735_ net487 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1018 net1056 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_2
Xfanout1007 net1011 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
X_10090_ _05562_ _05563_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__nand2_1
XFILLER_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06109__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07857__A1 top0.CPU.intMem_out\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12662_ clknet_leaf_66_clk _02297_ net1119 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08915__X _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11613_ net1305 _01252_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07609__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12593_ clknet_leaf_89_clk _02228_ net1079 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08806__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ net1236 _01183_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08282__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06435__X _03092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11475_ clknet_leaf_77_clk top0.CPU.internalMem.state_n\[0\] net1123 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.state\[0\] sky130_fd_sc_hd__dfstp_1
X_11193__845 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__inv_2
XANTENNA__08082__B net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234__886 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__inv_2
X_10288_ _02471_ _04958_ _04937_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08302__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12027_ net1719 _01666_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[520\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_120_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06348__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06757__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128__780 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__inv_2
XANTENNA__08257__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06450_ _03105_ _03106_ net870 vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06381_ _03023_ net539 vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__nor2_1
X_08120_ net2816 net223 net431 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XANTENNA__06492__S net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842__494 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__inv_2
X_08051_ net498 net177 net702 net437 net2458 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a32o_1
X_07002_ _03584_ net523 _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__a21o_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387__39 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__inv_2
XFILLER_89_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08025__B2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08953_ net214 net702 net271 net263 net2643 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__a32o_1
XANTENNA__11564__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ net637 _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__nand2_2
XANTENNA__08328__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1007_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__X _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ top0.CPU.register.registers\[244\] net565 vssd1 vssd1 vccd1 vccd1 _04762_
+ sky130_fd_sc_hd__or2_1
XFILLER_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07835_ top0.CPU.intMem_out\[29\] net627 _03003_ _02385_ net643 vssd1 vssd1 vccd1
+ vccd1 _04490_ sky130_fd_sc_hd__a221o_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06434__S1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ _03890_ _03910_ _02555_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__mux2_1
X_09505_ top0.MMIO.WBData_i\[3\] net149 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nand2b_1
X_06717_ top0.CPU.register.registers\[4\] top0.CPU.register.registers\[36\] top0.CPU.register.registers\[68\]
+ top0.CPU.register.registers\[100\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03374_
+ sky130_fd_sc_hd__mux4_1
X_09436_ top0.MMIO.WBData_i\[14\] _05026_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__and2_1
XANTENNA__08500__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07697_ net342 _04345_ _04346_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06648_ top0.CPU.register.registers\[770\] top0.CPU.register.registers\[802\] top0.CPU.register.registers\[834\]
+ top0.CPU.register.registers\[866\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03305_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05945__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ net2491 _04583_ net607 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
X_06579_ top0.CPU.register.registers\[400\] top0.CPU.register.registers\[432\] top0.CPU.register.registers\[464\]
+ top0.CPU.register.registers\[496\] net931 net897 vssd1 vssd1 vccd1 vccd1 _03236_
+ sky130_fd_sc_hd__mux4_1
X_11177__829 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__inv_2
XANTENNA_fanout801_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _04893_ _04925_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__or2_2
X_08318_ net2956 net159 net413 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__mux2_1
X_08249_ net210 net668 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10218__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06027__B1 _02683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06455__A1_N net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06122__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ net2577 net117 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__and2_1
XFILLER_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08122__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ top0.display.delayctr\[22\] _05596_ top0.display.delayctr\[23\] vssd1 vssd1
+ vccd1 vccd1 _05605_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07086__X _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ top0.display.delayctr\[8\] _05548_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__or2_1
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10785__437 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__inv_2
XANTENNA__06189__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05936__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ clknet_leaf_66_clk _02280_ net1102 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12576_ clknet_leaf_90_clk _02211_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10826__478 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__inv_2
X_11527_ net1219 _01166_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06266__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06361__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11458_ clknet_leaf_70_clk _01106_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10679__331 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__inv_2
Xhold309 top0.CPU.register.registers\[466\] vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
X_11389_ clknet_leaf_78_clk _01037_ net1111 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09636__B _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1009 net62 vssd1 vssd1 vccd1 vccd1 net3231 sky130_fd_sc_hd__dlygate4sd3_1
X_05950_ top0.CPU.register.registers\[1\] top0.CPU.register.registers\[33\] top0.CPU.register.registers\[65\]
+ top0.CPU.register.registers\[97\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02607_
+ sky130_fd_sc_hd__mux4_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05881_ top0.CPU.register.registers\[515\] top0.CPU.register.registers\[547\] top0.CPU.register.registers\[579\]
+ top0.CPU.register.registers\[611\] net828 net793 vssd1 vssd1 vccd1 vccd1 _02538_
+ sky130_fd_sc_hd__mux4_1
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07620_ net462 _03338_ net444 _04276_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__o31a_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07551_ _02477_ _03173_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__and2b_1
X_06502_ top0.CPU.register.registers\[531\] top0.CPU.register.registers\[563\] top0.CPU.register.registers\[595\]
+ top0.CPU.register.registers\[627\] net940 net906 vssd1 vssd1 vccd1 vccd1 _03159_
+ sky130_fd_sc_hd__mux4_1
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09140__C1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__X _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09691__B1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07482_ _04138_ _04134_ _04130_ _04135_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_45_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05927__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09221_ _02337_ _04882_ _04880_ top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 _04883_
+ sky130_fd_sc_hd__a211o_1
X_06433_ top0.CPU.register.registers\[23\] top0.CPU.register.registers\[55\] top0.CPU.register.registers\[87\]
+ top0.CPU.register.registers\[119\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03090_
+ sky130_fd_sc_hd__mux4_1
X_06364_ _02422_ _03020_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or2_1
X_09152_ _04710_ net274 net247 net2949 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a22o_1
XANTENNA__08246__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ net496 net165 net690 net433 net2472 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a32o_1
XFILLER_135_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09083_ net217 net620 net276 net257 net2402 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__a32o_1
X_06295_ net771 _02951_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__and2_2
X_08034_ net223 net703 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__and2_1
Xhold821 top0.CPU.register.registers\[989\] vssd1 vssd1 vccd1 vccd1 net3043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold810 top0.CPU.register.registers\[974\] vssd1 vssd1 vccd1 vccd1 net3032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 top0.CPU.register.registers\[909\] vssd1 vssd1 vccd1 vccd1 net3054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 net67 vssd1 vssd1 vccd1 vccd1 net3076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold843 net76 vssd1 vssd1 vccd1 vccd1 net3065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06009__B1 top0.CPU.control.funct7\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__Y _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold898 top0.CPU.register.registers\[54\] vssd1 vssd1 vccd1 vccd1 net3120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 top0.CPU.register.registers\[401\] vssd1 vssd1 vccd1 vccd1 net3109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 top0.CPU.register.registers\[921\] vssd1 vssd1 vccd1 vccd1 net3087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 top0.CPU.register.registers\[761\] vssd1 vssd1 vccd1 vccd1 net3098 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _05461_ _05466_ _05474_ net238 vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a31o_1
X_08936_ top0.CPU.register.registers\[208\] net570 net557 vssd1 vssd1 vccd1 vccd1
+ _04778_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout751_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ net722 net150 net280 net284 net2332 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09562__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06407__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__X _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _03785_ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__nor2_1
XFILLER_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08182__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472__124 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__inv_2
X_08798_ net677 _04738_ net288 net2829 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a22o_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10220__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__C1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07749_ net486 _04310_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a21oi_1
X_10513__165 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__inv_2
XFILLER_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09419_ _05009_ _05023_ net3406 _04949_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08237__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ net2122 _02069_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[923\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08788__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12361_ net2053 _02000_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[854\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06894__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12292_ net1984 _01931_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09737__A1 _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08960__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ top0.display.delayctr\[20\] _05587_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__or2_1
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10056_ net3439 net664 net602 _05538_ _05139_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_50_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08173__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346__998 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__inv_2
XANTENNA__07920__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11199__851 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__inv_2
X_12628_ clknet_leaf_93_clk _02263_ net1081 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
X_12559_ clknet_leaf_54_clk _02198_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08779__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06080_ top0.CPU.register.registers\[653\] top0.CPU.register.registers\[685\] top0.CPU.register.registers\[717\]
+ top0.CPU.register.registers\[749\] net850 net815 vssd1 vssd1 vccd1 vccd1 _02737_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07987__B1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold106 top0.CPU.register.registers\[752\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 top0.CPU.register.registers\[608\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top0.CPU.register.registers\[362\] vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05894__B _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 top0.CPU.register.registers\[961\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout608 net612 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_2
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06637__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456__108 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__inv_2
XANTENNA__08951__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ top0.CPU.internalMem.pcOut\[10\] _05267_ vssd1 vssd1 vccd1 vccd1 _05278_
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08697__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06982_ net544 _02927_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__nor2_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ net175 net3186 net357 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__mux2_1
X_05933_ net733 _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__or2_1
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ net175 net702 net310 net301 net2639 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_1_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05864_ _02519_ _02520_ net728 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ _04250_ _04253_ _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nand3b_2
X_08583_ net3134 net169 net336 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__mux2_1
X_05795_ top0.CPU.Op\[4\] _02424_ _02450_ _02376_ vssd1 vssd1 vccd1 vccd1 _02452_
+ sky130_fd_sc_hd__a22o_4
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout165_A _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07534_ _02534_ _03504_ _04164_ _04189_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__a221o_1
XFILLER_50_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ net337 _04035_ _04117_ net476 _03743_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__a221o_1
X_09204_ net770 top0.CPU.intMemAddr\[15\] top0.CPU.intMemAddr\[22\] top0.CPU.intMemAddr\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__or4_1
XANTENNA__06573__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06416_ net745 _03072_ _03066_ _03067_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_fanout1074_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__A2 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07396_ net485 _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nor2_1
X_09135_ top0.CPU.register.registers\[69\] net573 net559 vssd1 vssd1 vccd1 vccd1 _04838_
+ sky130_fd_sc_hd__o21a_1
X_06347_ net771 _03000_ _02992_ net584 vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__o211a_1
XFILLER_136_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ top0.CPU.register.registers\[115\] net576 vssd1 vssd1 vccd1 vccd1 _04815_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07442__A2 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06278_ net724 _02932_ net735 vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a21o_1
XANTENNA__06680__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06876__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__B2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09276__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout799_A top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ net3043 net440 _04639_ net503 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a22o_1
Xhold640 top0.CPU.register.registers\[799\] vssd1 vssd1 vccd1 vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold662 top0.CPU.register.registers\[625\] vssd1 vssd1 vccd1 vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 top0.CPU.register.registers\[473\] vssd1 vssd1 vccd1 vccd1 net2873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold673 top0.CPU.register.registers\[302\] vssd1 vssd1 vccd1 vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 top0.CPU.register.registers\[513\] vssd1 vssd1 vccd1 vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold695 top0.CPU.register.registers\[441\] vssd1 vssd1 vccd1 vccd1 net2917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08942__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _05459_ top0.CPU.internalMem.pcOut\[26\] vssd1 vssd1 vccd1 vccd1 _05460_
+ sky130_fd_sc_hd__and2b_1
XFILLER_77_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11033__685 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__inv_2
XANTENNA__07805__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ top0.CPU.register.registers\[220\] net566 vssd1 vssd1 vccd1 vccd1 _04773_
+ sky130_fd_sc_hd__or2_1
XFILLER_134_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ top0.CPU.internalMem.pcOut\[20\] _05396_ net647 vssd1 vssd1 vccd1 vccd1 _02197_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07083__Y _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ net1622 _01569_ net975 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[423\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371__23 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06800__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ net1553 _01500_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net1484 _01431_ net1083 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07130__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12413_ net2105 _02052_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[906\]
+ sky130_fd_sc_hd__dfrtp_1
X_12344_ net2036 _01983_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[837\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07969__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897__549 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__inv_2
X_12275_ net1967 _01914_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[768\]
+ sky130_fd_sc_hd__dfrtp_1
X_10641__293 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__inv_2
XANTENNA__06619__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ net577 net550 vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_108_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10039_ _05497_ _05512_ _05514_ _05525_ _05510_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__o311a_1
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07153__C _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07250_ _03905_ _03906_ net346 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_129_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06201_ top0.CPU.register.registers\[788\] top0.CPU.register.registers\[820\] top0.CPU.register.registers\[852\]
+ top0.CPU.register.registers\[884\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02858_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06307__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ net477 net518 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__nor2_1
XANTENNA__08621__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06132_ _02473_ _02772_ net582 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a21o_1
XANTENNA__06858__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06063_ top0.CPU.register.registers\[778\] top0.CPU.register.registers\[810\] top0.CPU.register.registers\[842\]
+ top0.CPU.register.registers\[874\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02720_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07543__C_N _03073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
XANTENNA__09177__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017__669 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__inv_2
Xfanout416 _04720_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_4
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_4
X_09822_ top0.CPU.internalMem.pcOut\[14\] _05313_ vssd1 vssd1 vccd1 vccd1 _05326_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08924__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__inv_2
Xfanout449 _02636_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_2
XANTENNA__06935__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06965_ _02927_ _02944_ net544 vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout282_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net152 net3286 net357 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__mux2_1
X_06896_ top0.CPU.register.registers\[136\] top0.CPU.register.registers\[168\] top0.CPU.register.registers\[200\]
+ top0.CPU.register.registers\[232\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03553_
+ sky130_fd_sc_hd__mux4_1
X_09684_ top0.CPU.decoder.instruction\[11\] _02448_ _02535_ net774 net590 vssd1 vssd1
+ vccd1 vccd1 _05198_ sky130_fd_sc_hd__a221o_1
X_05916_ net742 _02563_ _02571_ net584 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__o211ai_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05847_ net738 _02503_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__or2_1
XANTENNA__07896__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08635_ _04644_ net314 net302 net2730 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout547_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ net2942 net206 net334 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XANTENNA__09637__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ _04165_ _04167_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nor3_1
XANTENNA__09101__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05778_ top0.CPU.register.registers\[919\] top0.CPU.register.registers\[951\] top0.CPU.register.registers\[983\]
+ top0.CPU.register.registers\[1015\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02435_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08497_ _04698_ net395 net366 net2776 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a22o_1
X_10584__236 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__inv_2
XFILLER_50_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07448_ net448 _04104_ _04100_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__o21a_1
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ _03977_ _03981_ net456 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09118_ net200 net684 _04831_ net253 net3290 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a32o_1
XANTENNA__07359__X _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625__277 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09049_ net151 net624 net280 net258 net2638 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__a32o_1
X_12060_ net1752 _01699_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[553\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09168__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold470 net100 vssd1 vssd1 vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold481 top0.CPU.register.registers\[699\] vssd1 vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 top0.CPU.register.registers\[631\] vssd1 vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
X_10478__130 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__inv_2
Xfanout950 top0.CPU.decoder.instruction\[9\] vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_2
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08130__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout972 net976 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_2
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
Xhold1170 top0.MMIO.WBData_i\[25\] vssd1 vssd1 vccd1 vccd1 net3392 sky130_fd_sc_hd__dlygate4sd3_1
X_10519__171 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__inv_2
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1181 top0.display.delayctr\[10\] vssd1 vssd1 vccd1 vccd1 net3403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 top0.display.delayctr\[28\] vssd1 vssd1 vccd1 vccd1 net3414 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ net1605 _01552_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[406\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11844_ net1536 _01483_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ net1467 _01414_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__C net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload26 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_16
XTAP_TAPCELL_ROW_11_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11369__1021 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__inv_2
Xclkload15 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_2
Xclkload59 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_16
XANTENNA__06614__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload48 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_2
XANTENNA__08305__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload37 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_8
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ net2019 _01966_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[820\]
+ sky130_fd_sc_hd__dfrtp_1
X_12258_ net1950 _01897_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06090__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09159__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08367__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ net1881 _01828_ net1024 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[682\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07590__A1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07017__S1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _03263_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__nor2_1
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05701_ net767 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__inv_2
XANTENNA__07878__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06681_ net858 _03337_ _03330_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__o21ai_4
X_08420_ net954 net947 net952 net950 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__or4b_2
XFILLER_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06776__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ net713 net160 net391 net409 net2448 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a32o_1
X_08282_ net498 net215 net669 net417 net2482 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a32o_1
XANTENNA__07645__A2 _03463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07302_ _02477_ _03173_ net445 _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__o31a_1
X_07233_ _03888_ _03889_ net348 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__mux2_1
Xclkload9 clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_30_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05877__A2_N net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ net470 net524 _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a21bo_1
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06115_ net942 _02474_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07095_ _02416_ _03737_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__or2_1
XANTENNA__05959__A2 _02614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__X _05006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06046_ top0.CPU.register.registers\[776\] top0.CPU.register.registers\[808\] top0.CPU.register.registers\[840\]
+ top0.CPU.register.registers\[872\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02703_
+ sky130_fd_sc_hd__mux4_1
Xfanout202 _04556_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
Xfanout213 net216 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
XANTENNA_fanout497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net237 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout224 _04492_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_4
Xfanout279 net281 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ top0.CPU.internalMem.pcOut\[12\] _05293_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05310_ sky130_fd_sc_hd__a21o_1
X_07997_ top0.CPU.intMem_out\[2\] net630 _04588_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
X_09736_ _05226_ _05244_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a21oi_1
XFILLER_101_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06948_ top0.CPU.register.registers\[792\] top0.CPU.register.registers\[824\] top0.CPU.register.registers\[856\]
+ top0.CPU.register.registers\[888\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03605_
+ sky130_fd_sc_hd__mux4_1
X_09667_ _05114_ _05118_ _05117_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a21o_1
XANTENNA__06767__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout929_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ top0.CPU.register.registers\[265\] top0.CPU.register.registers\[297\] top0.CPU.register.registers\[329\]
+ top0.CPU.register.registers\[361\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03536_
+ sky130_fd_sc_hd__mux4_1
X_08618_ net718 net219 net318 net331 net2372 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__a32o_1
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout831_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07802__B _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _04957_ _05136_ net661 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__o21a_1
X_11145__797 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__inv_2
X_08549_ net216 net669 net390 net361 net2284 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a32o_1
XANTENNA__05895__A1 _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05990__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06418__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net1252 _01199_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08192__Y _04689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ clknet_leaf_90_clk _01130_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08125__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06153__B _02809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ net1804 _01751_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[605\]
+ sky130_fd_sc_hd__dfrtp_1
X_11039__691 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__inv_2
XFILLER_78_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08349__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ net1735 _01682_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[536\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10156__B1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07572__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_4
Xfanout791 net793 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09480__A top0.MMIO.WBData_i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08521__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ net1519 _01466_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05886__A1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05981__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ net1450 _01397_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload104 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__inv_6
X_11689_ net1381 _01328_ net1070 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[182\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload126 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__clkinv_16
Xclkload115 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__inv_8
XANTENNA__06344__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07260__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10953__605 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__inv_2
X_07920_ net3171 net548 net495 _04562_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09093__C _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ top0.CPU.internalMem.pcOut\[27\] net638 net633 _04503_ vssd1 vssd1 vccd1
+ vccd1 _04504_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_71_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_06802_ top0.CPU.register.registers\[396\] top0.CPU.register.registers\[428\] top0.CPU.register.registers\[460\]
+ top0.CPU.register.registers\[492\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03459_
+ sky130_fd_sc_hd__mux4_1
X_07782_ net487 net244 _04032_ _04087_ _04392_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__o32a_1
XANTENNA__08760__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ _05100_ _04864_ _02365_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__and3b_1
X_06733_ _03388_ _03389_ net760 vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__mux2_1
XANTENNA__08512__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__B2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ net131 net133 _05044_ net597 net3391 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__o32a_1
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06664_ net542 net471 net462 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_35_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09383_ net3003 _04494_ net606 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__mux2_1
XANTENNA__05877__B2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ net199 net695 net400 net379 net2389 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a32o_1
X_06595_ top0.CPU.register.registers\[775\] top0.CPU.register.registers\[807\] top0.CPU.register.registers\[839\]
+ top0.CPU.register.registers\[871\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03252_
+ sky130_fd_sc_hd__mux4_1
X_08334_ net3142 net412 net407 _04551_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XANTENNA__05972__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__X _03463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08265_ net3168 net420 _04717_ net516 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
X_08196_ net224 net689 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and2_1
X_07216_ net338 _03869_ _03872_ net485 net244 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a221o_1
X_07147_ net337 _03803_ _03719_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout781_A top0.CPU.control.rs2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout879_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ _03731_ _03734_ net346 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__mux2_1
X_10696__348 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__inv_2
XFILLER_10_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1019 net1021 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_4
Xfanout1008 net1011 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06029_ net454 _02650_ _02666_ _02684_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__or4b_2
XFILLER_113_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08346__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737__389 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__inv_2
XANTENNA__08751__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__C_N net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__C1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09719_ net241 _05227_ _05230_ _05110_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__o22ai_1
XFILLER_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08503__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368__1020 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__inv_2
XFILLER_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12661_ clknet_leaf_66_clk _02296_ net1104 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ net1304 _01251_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12592_ clknet_leaf_84_clk _02227_ net1107 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11543_ net1235 _01182_ net970 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_11474_ clknet_leaf_68_clk _01122_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct7\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07490__B1 _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08990__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10287_ net2757 net120 net113 _05664_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ net1718 _01665_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[519\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08742__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06979__S0 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06380_ net748 _03036_ _03027_ _03031_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__05897__B _02553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ net506 net219 net706 net438 net2314 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a32o_1
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07001_ _03584_ net523 _03603_ net522 vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__o22a_1
XANTENNA__09222__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08025__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net167 net708 _04782_ net265 net3306 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__a32o_1
XFILLER_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08981__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ _02386_ _02476_ net561 _04546_ _04547_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__o221a_4
XANTENNA__06013__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05890__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ _04540_ net555 _04761_ _04753_ net3021 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__a32o_1
X_07834_ _03886_ net231 net226 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__and3_1
XFILLER_69_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08733__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07765_ _03132_ _03246_ _03576_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout362_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ top0.MMIO.WBData_i\[24\] net149 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__and2_1
X_07696_ _04348_ _04349_ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__nand3_1
X_06716_ top0.CPU.register.registers\[132\] top0.CPU.register.registers\[164\] top0.CPU.register.registers\[196\]
+ top0.CPU.register.registers\[228\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03373_
+ sky130_fd_sc_hd__mux4_1
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07839__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09435_ net3395 net597 net131 _05033_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_84_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06647_ top0.CPU.register.registers\[898\] top0.CPU.register.registers\[930\] top0.CPU.register.registers\[962\]
+ top0.CPU.register.registers\[994\] net916 net882 vssd1 vssd1 vccd1 vccd1 _03304_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05945__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ net2634 _04589_ net608 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
X_06578_ _03233_ _03234_ net760 vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__mux2_1
XANTENNA__06536__X _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _04934_ top0.display.state\[2\] _04857_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__or3b_1
X_08317_ net3180 net161 net414 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__mux2_1
X_08248_ net2857 net417 _04709_ net499 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08179_ net509 net184 net621 net428 net2500 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a32o_1
X_10210_ net2713 net124 net116 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06027__B2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ _04971_ _05587_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__or2_2
XANTENNA__06122__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ net3396 net666 net602 _05550_ _05149_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a221o_1
XANTENNA__05881__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11160__812 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__inv_2
XFILLER_71_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06189__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05936__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12644_ clknet_leaf_65_clk _02279_ net1101 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_26_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201__853 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__inv_2
X_12575_ clknet_leaf_90_clk _02210_ net1079 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11526_ net1218 _01165_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06606__B _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06266__A1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06361__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ clknet_leaf_69_clk _01105_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct3\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06018__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05937__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ clknet_leaf_86_clk _01036_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08313__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ net2247 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08963__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05872__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__A0 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12009_ net1701 _01648_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05880_ top0.CPU.register.registers\[643\] top0.CPU.register.registers\[675\] top0.CPU.register.registers\[707\]
+ top0.CPU.register.registers\[739\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02537_
+ sky130_fd_sc_hd__mux4_1
XFILLER_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07453__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07172__B _03037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ _02496_ _03193_ _03960_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__and3b_1
X_06501_ top0.CPU.register.registers\[659\] top0.CPU.register.registers\[691\] top0.CPU.register.registers\[723\]
+ top0.CPU.register.registers\[755\] net940 net906 vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__mux4_1
X_09220_ top0.CPU.intMemAddr\[14\] top0.CPU.intMemAddr\[13\] _04867_ _04881_ vssd1
+ vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_66_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07481_ _04136_ _04137_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05927__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__D_N net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06432_ top0.CPU.register.registers\[151\] top0.CPU.register.registers\[183\] top0.CPU.register.registers\[215\]
+ top0.CPU.register.registers\[247\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03089_
+ sky130_fd_sc_hd__mux4_1
X_06363_ _03014_ _03019_ net743 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_2
XANTENNA__09443__A1 _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05701__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08246__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ net3382 net247 _04844_ _04709_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a22o_1
XANTENNA__09099__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ net179 net621 _04820_ net257 net3347 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__a32o_1
X_08102_ net497 net215 net691 net433 net2606 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a32o_1
X_10959__611 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__inv_2
X_10447__99 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__inv_2
X_06294_ _02947_ _02948_ _02949_ _02950_ net733 net739 vssd1 vssd1 vccd1 vccd1 _02951_
+ sky130_fd_sc_hd__mux4_1
X_08033_ net3187 net440 _04647_ net501 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a22o_1
Xhold800 top0.CPU.register.registers\[788\] vssd1 vssd1 vccd1 vccd1 net3022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 top0.CPU.register.registers\[1019\] vssd1 vssd1 vccd1 vccd1 net3033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout208_A _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 net80 vssd1 vssd1 vccd1 vccd1 net3044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06009__B2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 top0.CPU.register.registers\[922\] vssd1 vssd1 vccd1 vccd1 net3055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 top0.CPU.register.registers\[537\] vssd1 vssd1 vccd1 vccd1 net3077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 top0.CPU.register.registers\[181\] vssd1 vssd1 vccd1 vccd1 net3066 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 top0.CPU.register.registers\[654\] vssd1 vssd1 vccd1 vccd1 net3099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 top0.CPU.register.registers\[984\] vssd1 vssd1 vccd1 vccd1 net3088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 top0.CPU.register.registers\[885\] vssd1 vssd1 vccd1 vccd1 net3110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05863__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ _05461_ _05466_ _05474_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a21oi_1
Xhold899 top0.CPU.register.registers\[282\] vssd1 vssd1 vccd1 vccd1 net3121 sky130_fd_sc_hd__dlygate4sd3_1
X_08935_ _04650_ net269 net263 net2796 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__a22o_1
XANTENNA__08706__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _02403_ _04732_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__nor2_1
XANTENNA__09903__C1 top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ net946 net677 _04734_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__nand3_4
X_07817_ net233 net228 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__nand2_1
XFILLER_72_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ net338 _03888_ _03891_ _02577_ net244 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a221o_1
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ net484 _04333_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout911_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ net139 _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__nand2_1
XANTENNA__08194__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ _02338_ _04982_ _04984_ net629 _04973_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_23_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12360_ net2052 _01999_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08788__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12291_ net1983 _01930_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ _02868_ _05577_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10752__404 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__inv_2
X_10055_ _05536_ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__nand2_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09899__S net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09122__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08476__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__A1 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06031__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08308__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ clknet_leaf_75_clk _02262_ net1124 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12558_ clknet_leaf_54_clk _02197_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[20\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold107 top0.CPU.register.registers\[895\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
X_11509_ net1201 _01148_ net972 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12489_ net2181 _02128_ net1072 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[982\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold129 top0.CPU.register.registers\[687\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 top0.CPU.register.registers\[998\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06098__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08936__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 net610 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05845__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06981_ _03623_ net521 vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__and2_1
X_10495__147 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__inv_2
X_08720_ net219 net2922 net359 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__mux2_1
X_05932_ top0.CPU.register.registers\[384\] top0.CPU.register.registers\[416\] top0.CPU.register.registers\[448\]
+ top0.CPU.register.registers\[480\] net836 net801 vssd1 vssd1 vccd1 vccd1 _02589_
+ sky130_fd_sc_hd__mux4_1
X_08651_ net220 net706 net321 net303 net2384 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a32o_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05863_ top0.CPU.register.registers\[523\] top0.CPU.register.registers\[555\] top0.CPU.register.registers\[587\]
+ top0.CPU.register.registers\[619\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02520_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_1_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10536__188 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__inv_2
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07602_ _03841_ _03955_ _04258_ _04257_ net448 vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__a32o_1
XANTENNA__09113__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05794_ _02376_ _02450_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nand2_1
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08582_ net2861 net173 net335 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
XANTENNA__08467__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07533_ _03518_ _03973_ _02730_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nor3b_1
X_07464_ net339 _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nor2_1
XANTENNA__06022__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09203_ _04853_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__or2_1
XANTENNA__06527__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06415_ _03068_ _03069_ _03070_ _03071_ net759 net863 vssd1 vssd1 vccd1 vccd1 _03072_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ net171 net680 net271 net251 net2417 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1067_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07395_ _03893_ _04051_ net478 vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux2_1
X_06346_ _02455_ _03002_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__nand2_1
X_09065_ _04683_ net276 net257 net2544 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__a22o_1
X_06277_ net782 _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold630 top0.CPU.register.registers\[796\] vssd1 vssd1 vccd1 vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
X_08016_ net224 net712 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold663 top0.CPU.intMemAddr\[6\] vssd1 vssd1 vccd1 vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08927__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold652 top0.CPU.register.registers\[312\] vssd1 vssd1 vccd1 vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06262__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 top0.CPU.register.registers\[643\] vssd1 vssd1 vccd1 vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 top0.CPU.register.registers\[574\] vssd1 vssd1 vccd1 vccd1 net2918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 top0.CPU.register.registers\[318\] vssd1 vssd1 vccd1 vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 top0.CPU.register.registers\[781\] vssd1 vssd1 vccd1 vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout861_A top0.CPU.decoder.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ net585 _04506_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a21oi_2
XFILLER_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07805__B net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _04639_ net275 net264 net2831 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__a22o_1
X_09898_ _05395_ _05394_ _05393_ net236 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ net221 net3161 net354 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09104__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ net1552 _01499_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[353\]
+ sky130_fd_sc_hd__dfrtp_1
X_11791_ net1483 _01430_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08458__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07666__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07032__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12412_ net2104 _02051_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[905\]
+ sky130_fd_sc_hd__dfrtp_1
X_12343_ net2035 _01982_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[836\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272__924 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__inv_2
X_12274_ net1966 _01913_ net1054 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[767\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08630__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08918__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11313__965 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__inv_2
X_10107_ net3424 net665 net661 _05573_ _05576_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a221o_1
XANTENNA__08146__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _05523_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__12495__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06004__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ net1681 _01628_ net972 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10880__532 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06200_ _02855_ _02856_ net727 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XANTENNA__09658__A _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417__69 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__inv_2
X_07180_ net480 net518 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__nor2_1
XANTENNA__07409__B1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06131_ net579 _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__or2_1
XANTENNA__07449__Y _04106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06307__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921__573 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__inv_2
X_06062_ top0.CPU.register.registers\[906\] top0.CPU.register.registers\[938\] top0.CPU.register.registers\[970\]
+ top0.CPU.register.registers\[1002\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02719_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07178__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net408 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
Xfanout428 _04672_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_4
XANTENNA_clkload12_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ top0.CPU.internalMem.pcOut\[14\] _05313_ vssd1 vssd1 vccd1 vccd1 _05325_
+ sky130_fd_sc_hd__and2_1
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_4
X_09752_ _05258_ _05259_ top0.CPU.internalMem.pcOut\[9\] vssd1 vssd1 vccd1 vccd1 _05261_
+ sky130_fd_sc_hd__a21o_1
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07184__Y _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06964_ _03577_ _03578_ _03581_ _03601_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__a311o_2
X_08703_ net207 net3201 net358 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
XANTENNA__08137__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06895_ top0.CPU.register.registers\[392\] top0.CPU.register.registers\[424\] top0.CPU.register.registers\[456\]
+ top0.CPU.register.registers\[488\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03552_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09885__B2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _04248_ net232 net227 net632 vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a31o_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06021__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05915_ net742 _02563_ _02571_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout275_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05846_ _02501_ _02502_ net785 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06243__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _04643_ net306 net301 net2873 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a22o_1
X_05777_ _02416_ _02432_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__or2_1
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08565_ net3028 _04528_ net333 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
X_07516_ _04170_ _04171_ _04172_ _04169_ _04168_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__o2111ai_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ _04697_ net385 net365 net2673 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11256__908 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__inv_2
XANTENNA_fanout707_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ _03747_ _04102_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__o21a_1
XANTENNA__06320__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ _03978_ _04034_ net458 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__mux2_1
XFILLER_13_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_33_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11000__652 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__inv_2
X_09117_ top0.CPU.register.registers\[80\] net571 net557 vssd1 vssd1 vccd1 vccd1 _04831_
+ sky130_fd_sc_hd__o21a_1
X_06329_ top0.CPU.register.registers\[541\] top0.CPU.register.registers\[573\] top0.CPU.register.registers\[605\]
+ top0.CPU.register.registers\[637\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02986_
+ sky130_fd_sc_hd__mux4_1
X_09048_ net948 _04671_ _04732_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_94_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08612__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 top0.CPU.register.registers\[997\] vssd1 vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 top0.CPU.register.registers\[622\] vssd1 vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
X_10431__83 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__inv_2
XANTENNA__05809__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 top0.CPU.register.registers\[712\] vssd1 vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xhold493 top0.CPU.register.registers\[705\] vssd1 vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout951 top0.CPU.decoder.instruction\[9\] vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_2
Xfanout940 net941 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06482__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07027__S net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout973 net975 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout962 net1004 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_2
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_2
Xfanout995 net1004 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08679__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xhold1160 top0.CPU.register.registers\[60\] vssd1 vssd1 vccd1 vccd1 net3382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 top0.CPU.intMem_out\[9\] vssd1 vssd1 vccd1 vccd1 net3404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1193 top0.MISOtoMMIO\[5\] vssd1 vssd1 vccd1 vccd1 net3415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 top0.display.delayctr\[12\] vssd1 vssd1 vccd1 vccd1 net3393 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net1604 _01551_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[405\]
+ sky130_fd_sc_hd__dfrtp_1
X_11843_ net1535 _01482_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[336\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09242__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10864__516 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ net1466 _01413_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905__557 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__inv_2
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload16 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_8
Xclkload49 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__clkinv_8
Xclkload27 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_8
Xclkload38 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_16
X_12326_ net2018 _01965_ net1127 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[819\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758__410 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__inv_2
X_12257_ net1949 _01896_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[750\]
+ sky130_fd_sc_hd__dfrtp_1
X_12188_ net1880 _01827_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08119__A1 _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05700_ top0.MMIO.WBData_i\[29\] vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__inv_2
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06680_ _03333_ _03336_ net862 vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__mux2_1
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06776__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07180__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ net717 _04622_ net389 net409 net2297 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a32o_1
X_07301_ _02477_ _03173_ net340 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a21o_1
X_08281_ net510 net170 net674 net420 net2670 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a32o_1
X_07232_ _03793_ _03818_ net456 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__mux2_1
XFILLER_20_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07163_ net470 _03261_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__or2_1
XANTENNA__08055__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06114_ _02750_ _02769_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__and2_2
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07094_ _02416_ _03737_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__nor2_1
X_06045_ _02700_ _02701_ net728 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout203 _04556_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
XANTENNA__07636__A _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 net216 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
X_09804_ _05307_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__and2_1
Xfanout236 net237 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06540__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06908__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout247 _04842_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_8
Xfanout258 _04809_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07996_ net563 _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__or2_1
XFILLER_87_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06464__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout269 net281 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_4
X_09735_ _05221_ _05235_ _05234_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a21boi_1
X_06947_ top0.CPU.register.registers\[920\] top0.CPU.register.registers\[952\] top0.CPU.register.registers\[984\]
+ top0.CPU.register.registers\[1016\] net925 net891 vssd1 vssd1 vccd1 vccd1 _03604_
+ sky130_fd_sc_hd__mux4_1
X_10551__203 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__inv_2
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _05114_ _05118_ _05117_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06216__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06686__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06767__S1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06878_ top0.CPU.register.registers\[393\] top0.CPU.register.registers\[425\] top0.CPU.register.registers\[457\]
+ top0.CPU.register.registers\[489\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03535_
+ sky130_fd_sc_hd__mux4_1
X_08617_ net720 net179 net322 net331 net2466 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__a32o_1
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_38_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05829_ top0.CPU.register.registers\[274\] top0.CPU.register.registers\[306\] top0.CPU.register.registers\[338\]
+ top0.CPU.register.registers\[370\] net846 net811 vssd1 vssd1 vccd1 vccd1 _02486_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07802__C net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ _02572_ _05007_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout824_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ net169 net3060 net364 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07090__B net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05895__A2 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ net178 net619 net398 net371 net2422 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a32o_1
XANTENNA__09298__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11490_ clknet_leaf_83_clk top0.display.next_state\[2\] net1110 vssd1 vssd1 vccd1
+ vccd1 top0.display.state\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08046__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08061__A3 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ net1803 _01750_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[604\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09546__A0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net1734 _01681_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[535\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold290 top0.CPU.register.registers\[325\] vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10156__A1 _02942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09010__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout781 top0.CPU.control.rs2\[3\] vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_6
Xfanout770 top0.CPU.muxAddr.prev_control vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_2
XFILLER_93_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06758__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_47_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ net1518 _01465_ net1097 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[319\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09077__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ net1449 _01396_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[250\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08285__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278__930 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__inv_2
XANTENNA__08824__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11688_ net1380 _01327_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08316__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload127 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__clkinv_16
X_11319__971 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__inv_2
Xclkload116 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload105 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__inv_8
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08052__A3 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10992__644 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__inv_2
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ net2001 _01948_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09537__A0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09001__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ top0.CPU.intMem_out\[27\] net628 _04502_ net643 vssd1 vssd1 vccd1 vccd1 _04503_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_71_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06806__A1_N net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ _03456_ _03457_ net766 vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
X_07781_ net443 _04149_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nand2_1
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08760__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ _05094_ _05097_ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and3_1
X_06732_ top0.CPU.register.registers\[518\] top0.CPU.register.registers\[550\] top0.CPU.register.registers\[582\]
+ top0.CPU.register.registers\[614\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03389_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08287__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09451_ top0.MMIO.WBData_i\[19\] net146 net135 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__o21a_1
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06663_ _03303_ _03318_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_35_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09068__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09382_ net2564 _04500_ net606 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__mux2_1
X_06594_ top0.CPU.register.registers\[903\] top0.CPU.register.registers\[935\] top0.CPU.register.registers\[967\]
+ top0.CPU.register.registers\[999\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03251_
+ sky130_fd_sc_hd__mux4_1
X_08402_ _04666_ net389 net377 net2398 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08276__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08333_ net2920 net410 net392 _04545_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_125_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08264_ _04549_ _04705_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout238_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ net3018 net423 _04690_ net513 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
X_07215_ _03870_ _03871_ net346 vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__mux2_1
XANTENNA__09776__B1 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__X _04561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _03801_ _03802_ net465 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__mux2_1
X_07077_ _03732_ _03733_ net460 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__mux2_1
XANTENNA__06685__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071__723 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__inv_2
XANTENNA__09528__A0 top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06028_ _02650_ _02666_ _02684_ net449 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10401__53 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__inv_2
XANTENNA_fanout774_A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 net1011 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06701__C _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112__764 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07554__A2 _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _05228_ _05229_ net650 vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__o21a_1
X_07979_ top0.CPU.internalMem.pcOut\[6\] net640 net636 _04610_ vssd1 vssd1 vccd1 vccd1
+ _04611_ sky130_fd_sc_hd__o211a_4
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ net35 net3372 _05173_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12660_ clknet_leaf_66_clk _02295_ net1101 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ net1303 _01250_ net1009 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__11409__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ clknet_leaf_90_clk _02226_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_116_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08806__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08282__A3 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11542_ net1234 _01181_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ clknet_leaf_69_clk _01121_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct7\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10976__628 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10720__372 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__inv_2
XANTENNA__07793__A2 _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07276__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ _02493_ net550 _04937_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12268__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ net1717 _01664_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06979__S1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07215__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05876__A2_N _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06600__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ net1501 _01448_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[302\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_107_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08273__A3 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07000_ _03640_ net520 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nor2_1
X_11055__707 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__inv_2
XANTENNA__06667__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ top0.CPU.register.registers\[197\] net573 net559 vssd1 vssd1 vccd1 vccd1
+ _04782_ sky130_fd_sc_hd__o21a_1
XANTENNA__05795__A1 top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07186__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07902_ top0.CPU.internalMem.pcOut\[19\] net639 net625 top0.CPU.intMem_out\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o22a_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05890__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ top0.CPU.register.registers\[245\] net568 vssd1 vssd1 vccd1 vccd1 _04761_
+ sky130_fd_sc_hd__or2_1
X_07833_ net3164 net548 net514 _04488_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08729__B net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07764_ _04412_ _04413_ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o21ai_1
X_09503_ _02354_ net148 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nand2_1
X_06715_ _03368_ _03371_ net749 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__mux2_1
X_07695_ net448 _04350_ _04351_ _03757_ _03842_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__a32o_1
XANTENNA__08497__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ top0.MMIO.WBData_i\[13\] net145 _05028_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06646_ net478 _03283_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09365_ net2945 _04593_ net610 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
X_06577_ top0.CPU.register.registers\[16\] top0.CPU.register.registers\[48\] top0.CPU.register.registers\[80\]
+ top0.CPU.register.registers\[112\] net929 net895 vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__mux4_1
X_10663__315 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__inv_2
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ net2439 top0.CPU.internalMem.load2Ct_n\[0\] _04950_ vssd1 vssd1 vccd1 vccd1
+ top0.CPU.internalMem.load2Ct_n\[1\] sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08316_ net2993 net166 net413 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08247_ net211 net670 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704__356 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__inv_2
XANTENNA__08354__C_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ net506 net189 net619 net427 net2413 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout891_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09295__B _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06271__Y _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ _03039_ _03668_ net343 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07808__B _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10140_ _02446_ net551 net141 vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _05548_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__nand2_1
XANTENNA__05881__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__B1 top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07383__X _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08488__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06874__S net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07160__A0 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12643_ clknet_leaf_66_clk _02278_ net1104 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ clknet_leaf_90_clk _02209_ net1079 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11240__892 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__inv_2
XFILLER_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ net1217 _01164_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06897__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ clknet_leaf_67_clk _01104_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct3\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11387_ clknet_leaf_86_clk _01035_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10338_ net2236 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06974__B1 top0.CPU.decoder.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392__44 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__inv_2
XANTENNA__05872__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10269_ net2692 net120 net113 _05155_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
X_12008_ net1700 _01647_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[501\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06821__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08479__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06500_ net541 _02477_ _03116_ _03156_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__o22ai_4
X_07480_ _02908_ _03617_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_66_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06784__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06431_ top0.CPU.register.registers\[407\] top0.CPU.register.registers\[439\] top0.CPU.register.registers\[471\]
+ top0.CPU.register.registers\[503\] net910 net876 vssd1 vssd1 vccd1 vccd1 _03088_
+ sky130_fd_sc_hd__mux4_1
X_06362_ _03015_ _03016_ _03018_ _03017_ net785 net738 vssd1 vssd1 vccd1 vccd1 _03019_
+ sky130_fd_sc_hd__mux4_1
X_09150_ top0.CPU.register.registers\[60\] _02396_ net553 vssd1 vssd1 vccd1 vccd1
+ _04844_ sky130_fd_sc_hd__o21a_1
X_08101_ net510 net170 net697 net434 net2707 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a32o_1
X_09081_ top0.CPU.register.registers\[105\] net573 net559 vssd1 vssd1 vccd1 vccd1
+ _04820_ sky130_fd_sc_hd__o21a_1
XANTENNA__08651__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998__650 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__inv_2
X_06293_ top0.CPU.register.registers\[539\] top0.CPU.register.registers\[571\] top0.CPU.register.registers\[603\]
+ top0.CPU.register.registers\[635\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02950_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09396__A _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ net204 net712 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and2_1
XANTENNA__07909__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold812 top0.CPU.register.registers\[732\] vssd1 vssd1 vccd1 vccd1 net3034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold801 top0.CPU.register.registers\[410\] vssd1 vssd1 vccd1 vccd1 net3023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06091__Y _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 top0.CPU.register.registers\[790\] vssd1 vssd1 vccd1 vccd1 net3067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 top0.CPU.register.registers\[856\] vssd1 vssd1 vccd1 vccd1 net3056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 top0.CPU.register.registers\[249\] vssd1 vssd1 vccd1 vccd1 net3045 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__inv_2
Xhold878 net99 vssd1 vssd1 vccd1 vccd1 net3100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 net97 vssd1 vssd1 vccd1 vccd1 net3111 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06024__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold867 net89 vssd1 vssd1 vccd1 vccd1 net3089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 top0.CPU.register.registers\[629\] vssd1 vssd1 vccd1 vccd1 net3078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08934_ net202 net707 _04777_ net265 net3337 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__a32o_1
XANTENNA__06965__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1012_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05863__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _02398_ _02403_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_4_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06812__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ _03714_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__nand2_1
XANTENNA__07363__B net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06699__A1_N net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183__835 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__inv_2
X_08796_ net155 net682 net314 net290 net2443 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__a32o_1
X_07747_ _03738_ _04136_ _04138_ _03751_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11224__876 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__inv_2
XANTENNA__09682__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07678_ _02496_ net534 net445 _04334_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__o31a_1
XANTENNA__07142__A0 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08485__A3 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06694__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ top0.MMIO.WBData_i\[7\] _04933_ net143 top0.MISOtoMMIO\[7\] vssd1 vssd1 vccd1
+ vccd1 _05022_ sky130_fd_sc_hd__o22a_1
XANTENNA__08194__B net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06629_ top0.CPU.register.registers\[899\] top0.CPU.register.registers\[931\] top0.CPU.register.registers\[963\]
+ top0.CPU.register.registers\[995\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03286_
+ sky130_fd_sc_hd__mux4_1
X_09348_ _04863_ _04929_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06879__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08237__A3 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _02364_ _04929_ _04933_ _04862_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_97_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08642__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ net1982 _01929_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07538__B _03637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118__770 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__inv_2
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ net3410 net664 net662 _05586_ _05589_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10791__443 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__inv_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ top0.display.delayctr\[3\] _05533_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06803__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10832__484 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__inv_2
XANTENNA__07920__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07133__A0 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06031__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08881__B1 _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12626_ clknet_leaf_93_clk _02261_ net1081 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08228__A3 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ clknet_leaf_54_clk _02196_ net1041 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08633__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05948__S net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 top0.CPU.register.registers\[840\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
X_11508_ net1200 _01147_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12488_ net2180 _02127_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[981\]
+ sky130_fd_sc_hd__dfrtp_1
X_11439_ clknet_leaf_60_clk _01087_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold119 top0.CPU.register.registers\[418\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06098__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05845__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06980_ net746 _03636_ _03627_ _03631_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11167__819 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__inv_2
X_05931_ top0.CPU.register.registers\[256\] top0.CPU.register.registers\[288\] top0.CPU.register.registers\[320\]
+ top0.CPU.register.registers\[352\] net836 net801 vssd1 vssd1 vccd1 vccd1 _02588_
+ sky130_fd_sc_hd__mux4_1
X_08650_ net179 net708 net322 net303 net2556 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a32o_1
X_05862_ top0.CPU.register.registers\[651\] top0.CPU.register.registers\[683\] top0.CPU.register.registers\[715\]
+ top0.CPU.register.registers\[747\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02519_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07183__B _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08164__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07911__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_1_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07601_ _03744_ _03963_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nand2_1
XANTENNA__05922__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05922__B2 top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05793_ top0.CPU.Op\[3\] _02378_ _02381_ _02406_ vssd1 vssd1 vccd1 vccd1 _02450_
+ sky130_fd_sc_hd__or4_4
X_08581_ net2926 net178 net335 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07532_ _02717_ net524 _04021_ _03540_ _02698_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__a32o_1
XANTENNA__07470__Y _04127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07463_ _02650_ net532 vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__and2b_1
XANTENNA__06022__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08872__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ top0.CPU.internalMem.state\[0\] top0.CPU.internalMem.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _04864_ sky130_fd_sc_hd__and2b_1
X_06414_ top0.CPU.register.registers\[284\] top0.CPU.register.registers\[316\] top0.CPU.register.registers\[348\]
+ top0.CPU.register.registers\[380\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03071_
+ sky130_fd_sc_hd__mux4_1
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ net175 net680 net276 net253 net2571 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a32o_1
XANTENNA__07427__A1 _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05781__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07394_ net523 net522 net521 net520 net467 net456 vssd1 vssd1 vccd1 vccd1 _04051_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout318_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A _04603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06345_ top0.CPU.control.funct7\[4\] net644 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__nand2_1
XANTENNA__07427__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06276_ top0.CPU.register.registers\[922\] top0.CPU.register.registers\[954\] top0.CPU.register.registers\[986\]
+ top0.CPU.register.registers\[1018\] net825 net790 vssd1 vssd1 vccd1 vccd1 _02933_
+ sky130_fd_sc_hd__mux4_1
X_09064_ _04682_ net273 net256 net2573 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__a22o_1
XFILLER_135_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold620 top0.CPU.register.registers\[787\] vssd1 vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
X_08015_ net3323 net439 _04638_ net514 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10775__427 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__inv_2
Xhold653 top0.CPU.register.registers\[50\] vssd1 vssd1 vccd1 vccd1 net2875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 top0.CPU.register.registers\[644\] vssd1 vssd1 vccd1 vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold631 top0.CPU.register.registers\[665\] vssd1 vssd1 vccd1 vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold675 top0.CPU.register.registers\[520\] vssd1 vssd1 vccd1 vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 top0.CPU.register.registers\[907\] vssd1 vssd1 vccd1 vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 top0.CPU.register.registers\[538\] vssd1 vssd1 vccd1 vccd1 net2886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 top0.CPU.register.registers\[238\] vssd1 vssd1 vccd1 vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ net585 _02928_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nor2_1
XANTENNA__06689__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _04638_ net279 net266 net2612 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__a22o_1
X_09897_ top0.CPU.internalMem.pcOut\[20\] _05381_ net239 vssd1 vssd1 vccd1 vccd1 _05395_
+ sky130_fd_sc_hd__o21ai_1
X_10816__468 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__inv_2
XANTENNA__07805__C net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ net198 net3248 net355 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout854_A top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07902__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_28_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08779_ _04702_ net307 net289 net2841 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10669__321 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__inv_2
XANTENNA__07821__B net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ net1482 _01429_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06437__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09407__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12411_ net2103 _02050_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08615__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07969__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ net2034 _01981_ net988 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[835\]
+ sky130_fd_sc_hd__dfrtp_1
X_12273_ net1965 _01912_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08059__A_N net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08394__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ _05574_ _05575_ net601 vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a21oi_1
X_10362__14 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__inv_2
XANTENNA__08146__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ top0.CPU.internalMem.pcOut\[31\] _05522_ vssd1 vssd1 vccd1 vccd1 _05524_
+ sky130_fd_sc_hd__or2_1
XFILLER_88_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xclkbuf_leaf_87_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_108_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06628__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08319__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ net1680 _01627_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09004__A top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06004__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ clknet_leaf_81_clk _02244_ net1112 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07409__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10462__114 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__inv_2
X_06130_ net742 _02786_ _02777_ _02781_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__08621__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06061_ _02698_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__or2_1
XANTENNA__07178__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10503__155 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__inv_2
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09393__B _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _05320_ _05322_ net236 vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o21ai_1
Xfanout418 _04706_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
Xfanout429 net431 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06396__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09751_ top0.CPU.internalMem.pcOut\[9\] _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_
+ sky130_fd_sc_hd__nand3_1
X_06963_ _03618_ _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__or2_1
XANTENNA__06302__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_78_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_05914_ _02566_ _02567_ _02570_ net735 net772 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a221o_2
X_08702_ net208 net3274 net357 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
XANTENNA__08688__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06894_ top0.CPU.register.registers\[264\] top0.CPU.register.registers\[296\] top0.CPU.register.registers\[328\]
+ top0.CPU.register.registers\[360\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03551_
+ sky130_fd_sc_hd__mux4_1
X_09682_ top0.CPU.internalMem.pcOut\[3\] net651 _05193_ _05196_ vssd1 vssd1 vccd1
+ vccd1 _02180_ sky130_fd_sc_hd__o22a_1
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout170_A _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05845_ top0.CPU.register.registers\[911\] top0.CPU.register.registers\[943\] top0.CPU.register.registers\[975\]
+ top0.CPU.register.registers\[1007\] net851 net816 vssd1 vssd1 vccd1 vccd1 _02502_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07922__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06243__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ _04642_ net305 net301 net2664 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__a22o_1
X_05776_ _02416_ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__nor2_1
XANTENNA__09098__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ net2998 _04522_ net334 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08845__A0 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__A2 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07515_ net463 _03338_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08495_ _04696_ net395 net366 net2777 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a22o_1
XANTENNA__06825__X _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06320__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07446_ _03759_ _03789_ _03926_ _04101_ _03850_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o32a_1
X_11295__947 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__inv_2
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ _03519_ net525 net469 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__mux2_1
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_33_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06328_ top0.CPU.register.registers\[669\] top0.CPU.register.registers\[701\] top0.CPU.register.registers\[733\]
+ top0.CPU.register.registers\[765\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02985_
+ sky130_fd_sc_hd__mux4_1
X_09116_ _04702_ net269 net251 net2649 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__a22o_1
XANTENNA__08073__B2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11336__988 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__inv_2
X_09047_ net156 _04797_ _04808_ net350 net2911 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1132_X net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06259_ top0.CPU.register.registers\[153\] top0.CPU.register.registers\[185\] top0.CPU.register.registers\[217\]
+ top0.CPU.register.registers\[249\] net824 net790 vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__mux4_1
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 top0.CPU.register.registers\[223\] vssd1 vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 top0.CPU.register.registers\[633\] vssd1 vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 top0.CPU.register.registers\[896\] vssd1 vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 top0.CPU.intMemAddr\[13\] vssd1 vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold483 top0.CPU.register.registers\[373\] vssd1 vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout952 top0.CPU.decoder.instruction\[8\] vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_2
Xfanout941 top0.CPU.decoder.instruction\[15\] vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_8
Xfanout930 net938 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_4
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09949_ _05441_ _05442_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__nor2_1
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11189__841 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__inv_2
XFILLER_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07584__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout974 net975 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_4
Xfanout963 net965 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
Xfanout985 net995 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06482__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__X _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1150 top0.MISOtoMMIO\[0\] vssd1 vssd1 vccd1 vccd1 net3372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09523__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07336__A0 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1194 _02176_ vssd1 vssd1 vccd1 vccd1 net3416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 top0.MISOtoMMIO\[1\] vssd1 vssd1 vccd1 vccd1 net3383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 top0.CPU.intMem_out\[15\] vssd1 vssd1 vccd1 vccd1 net3405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 top0.CPU.intMem_out\[1\] vssd1 vssd1 vccd1 vccd1 net3394 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07832__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11911_ net1603 _01550_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[404\]
+ sky130_fd_sc_hd__dfrtp_1
X_11842_ net1534 _01481_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[335\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07551__B _03173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11773_ net1465 _01412_ net1024 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944__596 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__inv_2
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload17 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_8
X_12325_ net2017 _01964_ net1036 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[818\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload28 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_16
Xclkload39 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_16
XTAP_TAPCELL_ROW_11_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12256_ net1948 _01895_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08367__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12187_ net1879 _01826_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838__490 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__inv_2
XANTENNA__07575__B1 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07878__A1 top0.CPU.intMem_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09005__Y _04798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__A3 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05984__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07300_ _02578_ _03727_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__or2_1
XANTENNA__08827__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ net505 net174 net677 net419 net2279 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a32o_1
XFILLER_32_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07231_ _03790_ _03794_ _02617_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__mux2_1
X_11023__675 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__inv_2
X_07162_ _03817_ _03818_ net459 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__mux2_1
XANTENNA__08055__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06113_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__inv_2
XFILLER_8_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06161__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07093_ net519 _03701_ _03748_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06380__X _03037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06044_ top0.CPU.register.registers\[520\] top0.CPU.register.registers\[552\] top0.CPU.register.registers\[584\]
+ top0.CPU.register.registers\[616\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02701_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07636__B _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 _04539_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
X_09803_ _05305_ _05306_ _02350_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__o21ai_1
Xfanout237 _05109_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
Xfanout226 _04473_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07995_ _04275_ net233 net228 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__and3_1
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06464__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_4
Xfanout248 _04842_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
X_09734_ _05220_ _05236_ _05234_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__o21a_1
XFILLER_101_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10590__242 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__inv_2
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06946_ _02908_ _03602_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06877_ _03532_ _03533_ net760 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__mux2_1
X_09665_ net768 _05178_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__xor2_1
XANTENNA__06216__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887__539 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__inv_2
X_08616_ net720 net182 net323 net331 net2731 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05828_ net738 _02480_ _02483_ _02484_ net773 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_38_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07802__D net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ net2850 net604 net658 net3354 _05135_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__a221o_1
XANTENNA__05975__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631__283 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__inv_2
XANTENNA__08818__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05759_ _02413_ _02414_ _02412_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a21oi_2
X_08547_ net173 net672 net398 net363 net2265 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__a32o_1
X_08478_ net217 net619 net399 net371 net2379 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a32o_1
XFILLER_11_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ _04084_ _04085_ _04080_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__or3b_1
XANTENNA__08046__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08597__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ net1802 _01749_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[603\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 top0.CPU.register.registers\[486\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08349__A2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_12041_ net1733 _01680_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[534\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold291 top0.CPU.register.registers\[326\] vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10156__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net763 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06877__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout782 net787 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_4
Xfanout771 net775 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_4
Xfanout793 net799 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09849__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A _02578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08521__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_47_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11825_ net1517 _01464_ net1050 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[318\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08809__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08285__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007__659 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__inv_2
X_11756_ net1448 _01395_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[249\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ net1379 _01326_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[180\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06391__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08037__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload128 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload128/Y sky130_fd_sc_hd__clkinv_16
Xclkload106 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_6
Xclkload117 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_58_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12308_ net2000 _01947_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[801\]
+ sky130_fd_sc_hd__dfrtp_1
X_12239_ net1931 _01878_ net1001 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[732\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574__226 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__inv_2
X_06800_ top0.CPU.register.registers\[12\] top0.CPU.register.registers\[44\] top0.CPU.register.registers\[76\]
+ top0.CPU.register.registers\[108\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03457_
+ sky130_fd_sc_hd__mux4_1
XFILLER_110_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07780_ _03740_ _04148_ _04147_ net445 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08760__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ top0.CPU.register.registers\[646\] top0.CPU.register.registers\[678\] top0.CPU.register.registers\[710\]
+ top0.CPU.register.registers\[742\] net915 net882 vssd1 vssd1 vccd1 vccd1 _03388_
+ sky130_fd_sc_hd__mux4_1
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09450_ net130 net133 _05043_ net598 net3375 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__o32a_1
X_10615__267 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__inv_2
XANTENNA__08512__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06088__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ net203 net695 net406 net379 net2532 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a32o_1
XFILLER_64_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_06662_ _03303_ _03317_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__nor2_1
XANTENNA__06960__A1_N net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09381_ net2451 _04506_ net606 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__mux2_1
X_06593_ _02667_ _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09399__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ net2851 net410 net396 _04540_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
X_08263_ net3277 net419 _04716_ net508 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
X_10468__120 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ _03730_ _03765_ net459 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__mux2_1
X_10509__161 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__inv_2
X_08194_ net212 net688 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__and2_1
XANTENNA__09776__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07145_ net523 net520 net475 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__mux2_1
X_10398__50 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__inv_2
XANTENNA__07647__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ _03519_ net526 net468 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__mux2_1
XANTENNA__06551__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06027_ top0.CPU.control.funct7\[1\] _02518_ _02683_ net579 vssd1 vssd1 vccd1 vccd1
+ _02684_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__06685__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ top0.CPU.intMem_out\[6\] net629 _04588_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06697__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ top0.CPU.internalMem.pcOut\[5\] _05207_ top0.CPU.internalMem.pcOut\[6\] vssd1
+ vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12567__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06929_ top0.CPU.register.registers\[537\] top0.CPU.register.registers\[569\] top0.CPU.register.registers\[601\]
+ top0.CPU.register.registers\[633\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03586_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout934_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08503__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _02360_ top0.chipSelectTFT _05171_ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_
+ sky130_fd_sc_hd__or4_4
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ top0.display.counter\[1\] top0.display.counter\[0\] vssd1 vssd1 vccd1 vccd1
+ _05124_ sky130_fd_sc_hd__and2_1
XFILLER_43_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_100_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ clknet_leaf_83_clk _02225_ net1110 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11610_ net1302 _01249_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_11541_ net1233 _01180_ net972 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06278__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ clknet_leaf_67_clk _01120_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct7\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08019__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06125__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__B net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08990__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10285_ net3254 net119 net112 _05578_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a22o_1
XANTENNA__07276__B _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ net1716 _01663_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[517\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07844__X _04498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07950__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _02417_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07637__A_N _04106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload9_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06600__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11808_ net1500 _01447_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__S _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08258__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11739_ net1431 _01378_ net1009 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[232\]
+ sky130_fd_sc_hd__dfrtp_1
X_11094__746 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__inv_2
XANTENNA__08430__A1 _04528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ net171 net702 net271 net263 net2453 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__a32o_1
X_11135__787 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07901_ _03966_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__and3_2
X_08881_ _04534_ net555 _04760_ _04753_ net2963 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__a32o_1
X_07832_ net722 net212 vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__and2_1
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ top0.MMIO.WBData_i\[25\] net138 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or2_1
X_07763_ net452 _04419_ _04418_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o21a_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06714_ _03369_ _03370_ net757 vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__mux2_1
X_07694_ net483 _04079_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout250_A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ net3381 net597 net130 _05032_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_84_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11029__681 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__inv_2
X_06645_ _03285_ net531 vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nor2_1
X_09364_ net2631 _04597_ net608 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
X_06576_ top0.CPU.register.registers\[144\] top0.CPU.register.registers\[176\] top0.CPU.register.registers\[208\]
+ top0.CPU.register.registers\[240\] net929 net895 vssd1 vssd1 vccd1 vccd1 _03233_
+ sky130_fd_sc_hd__mux4_1
X_08315_ net2802 net215 net413 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__mux2_1
XFILLER_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ top0.CPU.internalMem.load2Ct\[1\] _04948_ top0.CPU.internalMem.load2Ct\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__and3b_1
XANTENNA__06355__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ net2910 net418 _04708_ net503 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a22o_1
X_08177_ net515 net190 net624 net428 net2366 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743__395 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09749__A1 _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ _03708_ net343 _03717_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__a31oi_4
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07808__C _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07059_ net544 _03714_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or2_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ top0.display.delayctr\[7\] _05545_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__nand2_1
XANTENNA__08700__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09921__A1 top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08185__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06220__S net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ clknet_leaf_66_clk _02277_ net1104 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06594__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07160__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ clknet_leaf_75_clk net767 net1125 vssd1 vssd1 vccd1 vccd1 top0.wishbone0.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06897__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11524_ net1216 _01163_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07999__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ clknet_leaf_69_clk _01103_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct3\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xwire243 _02890_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_1
X_11386_ clknet_leaf_86_clk _01034_ net1115 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06649__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ net2248 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06974__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08963__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10268_ net3100 net120 net113 _05656_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a22o_1
XANTENNA__08176__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ net1699 _01646_ net1000 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[500\]
+ sky130_fd_sc_hd__dfrtp_1
X_10199_ net3076 net122 _05644_ _04922_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XFILLER_66_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06821__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10286__A1 _02493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686__338 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__inv_2
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07151__A1 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06430_ top0.CPU.register.registers\[279\] top0.CPU.register.registers\[311\] top0.CPU.register.registers\[343\]
+ top0.CPU.register.registers\[375\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03087_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_66_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06361_ top0.CPU.register.registers\[30\] top0.CPU.register.registers\[62\] top0.CPU.register.registers\[94\]
+ top0.CPU.register.registers\[126\] net850 net815 vssd1 vssd1 vccd1 vccd1 _03018_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08100__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ net182 net622 net277 net257 net2427 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a32o_1
X_08100_ net505 net173 net694 net434 net2423 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a32o_1
X_06292_ top0.CPU.register.registers\[667\] top0.CPU.register.registers\[699\] top0.CPU.register.registers\[731\]
+ top0.CPU.register.registers\[763\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02949_
+ sky130_fd_sc_hd__mux4_1
X_10727__379 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__inv_2
X_08031_ net2961 net440 _04646_ net500 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
Xhold802 top0.CPU.register.registers\[500\] vssd1 vssd1 vccd1 vccd1 net3024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 top0.CPU.register.registers\[287\] vssd1 vssd1 vccd1 vccd1 net3046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 top0.CPU.register.registers\[524\] vssd1 vssd1 vccd1 vccd1 net3035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 top0.CPU.register.registers\[763\] vssd1 vssd1 vccd1 vccd1 net3068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 top0.CPU.register.registers\[760\] vssd1 vssd1 vccd1 vccd1 net3057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold868 top0.CPU.register.registers\[94\] vssd1 vssd1 vccd1 vccd1 net3090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 top0.CPU.register.registers\[766\] vssd1 vssd1 vccd1 vccd1 net3079 sky130_fd_sc_hd__dlygate4sd3_1
X_10368__20 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__inv_2
X_09982_ top0.CPU.internalMem.pcOut\[27\] _05472_ vssd1 vssd1 vccd1 vccd1 _05473_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__08954__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold879 net70 vssd1 vssd1 vccd1 vccd1 net3101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08933_ top0.CPU.register.registers\[210\] net574 net558 vssd1 vssd1 vccd1 vccd1
+ _04777_ sky130_fd_sc_hd__o21a_1
XANTENNA__07925__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net948 _02391_ _04732_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__or3_4
XANTENNA__06812__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06040__S net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__A3 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ _03703_ _03785_ _04456_ _04457_ _04469_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_4_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ net158 net679 net306 net289 net2725 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a32o_1
X_07746_ _02908_ net522 net341 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_38_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ net3368 _04949_ _05021_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__a21o_1
XANTENNA__06576__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07677_ _02496_ net534 net340 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a21o_1
XANTENNA__07142__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06628_ net484 _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ _04863_ _04994_ _04935_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__o21a_1
XFILLER_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06559_ net749 _03215_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__nor2_1
X_09278_ _02361_ net3444 _04939_ top0.wishbone0.curr_state\[0\] vssd1 vssd1 vccd1
+ vccd1 _00002_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06879__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ net511 net181 net685 net424 net2429 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a32o_1
XANTENNA__07819__B top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07850__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08945__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ _05587_ _05588_ net601 vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_128_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08430__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10053_ top0.display.delayctr\[3\] _05533_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__A3 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05916__C1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09122__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09261__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07133__A1 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_42_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ clknet_leaf_74_clk _02260_ net1125 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06892__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ clknet_leaf_54_clk _02195_ net1041 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06319__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06473__X _03130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ net1198 _01146_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12487_ net2179 _02126_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[980\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold109 top0.CPU.register.registers\[108\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ clknet_leaf_68_clk _01086_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08936__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05930_ net739 _02582_ _02585_ _02586_ net742 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a221o_1
X_05861_ _02452_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__nand2_4
X_08580_ net2897 net219 net335 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07372__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07600_ net482 _03983_ _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a21o_1
XANTENNA__09113__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05792_ _02338_ top0.CPU.Op\[4\] top0.CPU.Op\[3\] _02373_ vssd1 vssd1 vccd1 vccd1
+ _02449_ sky130_fd_sc_hd__or4_4
XFILLER_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07531_ _04160_ _04186_ _02515_ _03425_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a2bb2o_1
X_11247__899 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__inv_2
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07462_ net532 net444 vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__nor2_1
X_09201_ top0.CPU.internalMem.prev_busy_o _04861_ vssd1 vssd1 vccd1 vccd1 _04863_
+ sky130_fd_sc_hd__nand2_2
X_07393_ net454 _03742_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2_2
X_06413_ top0.CPU.register.registers\[412\] top0.CPU.register.registers\[444\] top0.CPU.register.registers\[476\]
+ top0.CPU.register.registers\[508\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03070_
+ sky130_fd_sc_hd__mux4_1
X_10351__3 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__inv_2
X_09132_ net3297 net253 _04837_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a21o_1
X_06344_ net771 _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__or2_1
XANTENNA__05781__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08624__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06275_ top0.CPU.register.registers\[794\] top0.CPU.register.registers\[826\] top0.CPU.register.registers\[858\]
+ top0.CPU.register.registers\[890\] net825 net790 vssd1 vssd1 vccd1 vccd1 _02932_
+ sky130_fd_sc_hd__mux4_1
X_09063_ _04681_ net273 net256 net2654 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__a22o_1
XANTENNA__06635__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ net212 net711 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__and2_1
Xhold610 top0.CPU.register.registers\[528\] vssd1 vssd1 vccd1 vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 net45 vssd1 vssd1 vccd1 vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 top0.CPU.register.registers\[784\] vssd1 vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold643 top0.CPU.register.registers\[827\] vssd1 vssd1 vccd1 vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 top0.CPU.register.registers\[379\] vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150__802 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__inv_2
Xhold687 top0.CPU.register.registers\[947\] vssd1 vssd1 vccd1 vccd1 net2909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top0.CPU.register.registers\[926\] vssd1 vssd1 vccd1 vccd1 net2898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07655__A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 top0.CPU.register.registers\[893\] vssd1 vssd1 vccd1 vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout582_A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ top0.CPU.internalMem.pcOut\[25\] net645 _05457_ vssd1 vssd1 vccd1 vccd1 _02202_
+ sky130_fd_sc_hd__o21ba_1
Xhold698 top0.CPU.register.registers\[756\] vssd1 vssd1 vccd1 vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07038__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net150 net710 net280 net266 net2672 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a32o_1
X_09896_ top0.CPU.internalMem.pcOut\[20\] _05381_ vssd1 vssd1 vccd1 vccd1 _05394_
+ sky130_fd_sc_hd__and2_1
XFILLER_112_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07942__X _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _04566_ net3189 net355 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ net202 net684 net319 net291 net2629 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__a32o_1
XFILLER_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ net442 _04133_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06549__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ net2102 _02049_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08615__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08425__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10256__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ net2033 _01980_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[834\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12272_ net1964 _01911_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08379__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08918__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09764__B top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ top0.display.delayctr\[16\] _05569_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__nand2_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09343__A2 top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ top0.CPU.internalMem.pcOut\[31\] _05522_ vssd1 vssd1 vccd1 vccd1 _05523_
+ sky130_fd_sc_hd__nand2_1
XFILLER_76_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10949__601 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__inv_2
XANTENNA__08551__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11987_ net1679 _01626_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07657__A2 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12608_ clknet_leaf_81_clk _02243_ net1112 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
X_12539_ clknet_leaf_83_clk _02178_ net1110 vssd1 vssd1 vccd1 vccd1 top0.display.reading_flag
+ sky130_fd_sc_hd__dfrtp_1
X_06060_ _02715_ net579 top0.CPU.control.funct7\[3\] _02518_ vssd1 vssd1 vccd1 vccd1
+ _02717_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06712__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10542__194 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__inv_2
Xfanout408 _04722_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_4
Xfanout419 net420 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
XANTENNA__08385__A3 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ top0.CPU.control.funct7\[4\] _02453_ net590 vssd1 vssd1 vccd1 vccd1 _05259_
+ sky130_fd_sc_hd__a21o_1
X_06962_ _03603_ net522 vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__and2_1
XANTENNA__08790__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ net241 _05194_ _05195_ net652 vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a31o_1
X_05913_ _02568_ _02569_ net725 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__mux2_1
X_08701_ net209 net3023 net357 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
X_06893_ net864 _03545_ _03548_ _03549_ net860 vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__o221a_1
XANTENNA__08542__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06779__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _04641_ net307 net301 net2809 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a22o_1
X_05844_ top0.CPU.register.registers\[783\] top0.CPU.register.registers\[815\] top0.CPU.register.registers\[847\]
+ top0.CPU.register.registers\[879\] net851 net816 vssd1 vssd1 vccd1 vccd1 _02501_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11386__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05775_ _02423_ _02427_ _02430_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout163_A _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ net3077 net208 net333 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__mux2_1
X_07514_ net471 _03356_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__nor2_1
X_08494_ _04695_ net387 net365 net2655 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a22o_1
XFILLER_35_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ _03833_ _03962_ _04101_ net489 vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout428_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout330_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06951__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ _03719_ _03877_ _03926_ _03933_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_33_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ net202 net689 _04830_ net253 net3313 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06327_ _02927_ _02944_ _02962_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__and4_1
XANTENNA__08073__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ top0.CPU.register.registers\[128\] net568 vssd1 vssd1 vccd1 vccd1 _04808_
+ sky130_fd_sc_hd__or2_1
X_06258_ _02911_ _02912_ _02913_ _02914_ net724 net736 vssd1 vssd1 vccd1 vccd1 _02915_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout797_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 top0.CPU.register.registers\[683\] vssd1 vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 top0.CPU.register.registers\[679\] vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 top0.CPU.register.registers\[599\] vssd1 vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ top0.CPU.register.registers\[405\] top0.CPU.register.registers\[437\] top0.CPU.register.registers\[469\]
+ top0.CPU.register.registers\[501\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02846_
+ sky130_fd_sc_hd__mux4_1
Xhold484 top0.CPU.register.registers\[591\] vssd1 vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold495 top0.CPU.register.registers\[231\] vssd1 vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 top0.CPU.register.registers\[324\] vssd1 vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08781__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout942 top0.CPU.control.funct3\[2\] vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
Xfanout931 net938 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
X_09948_ _05437_ _05440_ net235 vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__o21ai_1
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_4
Xfanout953 top0.CPU.decoder.instruction\[8\] vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_1
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_2
XFILLER_58_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout964 net968 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
Xfanout986 net988 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1151 _02171_ vssd1 vssd1 vccd1 vccd1 net3373 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ top0.CPU.internalMem.pcOut\[18\] _05362_ _05365_ _05366_ vssd1 vssd1 vccd1
+ vccd1 _05378_ sky130_fd_sc_hd__o2bb2a_1
Xhold1140 top0.display.delayctr\[11\] vssd1 vssd1 vccd1 vccd1 net3362 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout997 net1001 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07336__A1 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11910_ net1602 _01549_ net1119 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[403\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1173 top0.CPU.intMem_out\[13\] vssd1 vssd1 vccd1 vccd1 net3395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _02172_ vssd1 vssd1 vccd1 vccd1 net3384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1184 top0.CPU.intMem_out\[7\] vssd1 vssd1 vccd1 vccd1 net3406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07832__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07887__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1195 top0.CPU.intMem_out\[26\] vssd1 vssd1 vccd1 vccd1 net3417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11841_ net1533 _01480_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[334\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11772_ net1464 _01411_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[265\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10485__137 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__inv_2
Xclkload29 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_11_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12324_ net2016 _01963_ net995 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[817\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload18 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_6
X_10526__178 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__inv_2
X_12255_ net1947 _01894_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[748\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09494__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422__74 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__inv_2
XFILLER_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12186_ net1878 _01825_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[679\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08772__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08524__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05814__Y _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net652 _05503_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__o31a_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05984__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08827__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07230_ _03076_ _03666_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__and2_1
X_07161_ _03482_ net528 net468 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08055__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06112_ net582 _02768_ _02767_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__o21bai_4
XFILLER_9_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06161__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07092_ _03703_ _03738_ _03740_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06043_ top0.CPU.register.registers\[648\] top0.CPU.register.registers\[680\] top0.CPU.register.registers\[712\]
+ top0.CPU.register.registers\[744\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02700_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07636__C _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _04533_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
X_09802_ _02350_ _05305_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__or3_1
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
Xfanout238 net240 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
Xfanout216 _04618_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08763__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_4
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07994_ net716 net493 net165 net546 net2440 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout280_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ net650 _05242_ _05243_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a21oi_1
X_06945_ _02457_ net243 _02433_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08515__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__A1 _02578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ top0.CPU.register.registers\[9\] top0.CPU.register.registers\[41\] top0.CPU.register.registers\[73\]
+ top0.CPU.register.registers\[105\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03533_
+ sky130_fd_sc_hd__mux4_1
X_09664_ net768 _05178_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__nor2_1
X_11262__914 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__inv_2
XANTENNA_fanout378_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05827_ net785 _02481_ net778 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a21o_1
X_08615_ net718 net186 net318 net331 net2744 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a32o_1
X_09595_ _04957_ _05134_ net661 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout545_A _02400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05975__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05758_ _02339_ _02371_ _02373_ _02407_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__or4_1
X_08546_ net178 net672 net398 net363 net2535 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a32o_1
X_11303__955 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__inv_2
X_08477_ net179 net621 net401 net372 net2318 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a32o_1
X_05689_ net773 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07428_ _03835_ _03925_ net451 _03745_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__a211oi_1
X_07359_ net342 _03990_ _04006_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__a211o_2
XANTENNA__07099__B _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08703__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ _04581_ net3188 net351 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__mux2_1
XANTENNA__08349__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 top0.CPU.register.registers\[352\] vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ net1732 _01679_ net1077 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[533\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08754__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 top0.CPU.register.registers\[207\] vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
X_10870__522 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__inv_2
Xhold281 top0.CPU.register.registers\[203\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout750 net755 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_2
XANTENNA__08506__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout761 net763 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07309__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout772 net775 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_8
Xfanout783 net787 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout794 net796 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10911__563 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__inv_2
XANTENNA__08521__A3 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_47_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11824_ net1516 _01463_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11046__698 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ net1447 _01394_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[248\]
+ sky130_fd_sc_hd__dfrtp_1
X_11686_ net1378 _01325_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06391__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08037__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload107 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__clkinv_16
Xclkload118 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08993__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ net1999 _01946_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[800\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238_ net1930 _01877_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08745__B1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12169_ net1861 _01808_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11660__RESET_B net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06508__C1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ _02684_ _03248_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09170__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08512__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__inv_2
XFILLER_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _04665_ net407 net380 net2868 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
XFILLER_92_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_86_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09380_ net2721 _04512_ net606 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__mux2_1
X_06592_ _02651_ _02684_ _03247_ net542 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a31o_1
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08331_ net3303 net410 net395 _04534_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
X_08262_ net223 net673 vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__and2_1
XANTENNA__06287__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06308__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07213_ _03761_ _03766_ net456 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
X_08193_ net512 net150 net687 net424 net2753 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout126_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A0 _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ net537 net522 net473 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__mux2_1
XFILLER_106_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07075_ net524 net525 net468 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux2_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08984__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06026_ net741 _02682_ _02675_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a21oi_2
X_10854__506 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__inv_2
XANTENNA__08736__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05882__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A3 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ net562 _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__or2_1
XANTENNA__06211__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ top0.CPU.internalMem.pcOut\[6\] top0.CPU.internalMem.pcOut\[5\] _05207_ vssd1
+ vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__and3_1
X_06928_ top0.CPU.register.registers\[665\] top0.CPU.register.registers\[697\] top0.CPU.register.registers\[729\]
+ top0.CPU.register.registers\[761\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03585_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09161__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05970__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06859_ top0.CPU.register.registers\[266\] top0.CPU.register.registers\[298\] top0.CPU.register.registers\[330\]
+ top0.CPU.register.registers\[362\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03516_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ top0.display.counter\[4\] top0.display.counter\[3\] vssd1 vssd1 vccd1 vccd1
+ _05172_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06070__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ top0.display.counter\[1\] top0.display.counter\[0\] vssd1 vssd1 vccd1 vccd1
+ _05123_ sky130_fd_sc_hd__or2_1
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10748__400 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__inv_2
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08529_ _04714_ net388 net361 net3004 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a22o_1
XANTENNA__06278__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06285__Y _02942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ net1232 _01179_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ clknet_leaf_60_clk _01119_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct7\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08019__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08433__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06125__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05884__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ net3016 net120 net113 _05663_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a22o_1
X_12023_ net1715 _01662_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[516\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597__249 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06888__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06738__C1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_53_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07950__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout591 _02385_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_2
Xfanout580 _02422_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_53_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09152__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_46_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07702__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ net1499 _01446_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[300\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08258__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11738_ net1430 _01377_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[231\]
+ sky130_fd_sc_hd__dfrtp_1
X_11669_ net1361 _01308_ net970 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[162\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06652__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07900_ net2894 net548 net498 _04545_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a22o_1
X_08880_ top0.CPU.register.registers\[246\] net568 vssd1 vssd1 vccd1 vccd1 _04760_
+ sky130_fd_sc_hd__or2_1
X_07831_ top0.CPU.internalMem.pcOut\[30\] net638 net633 _04486_ vssd1 vssd1 vccd1
+ vccd1 _04487_ sky130_fd_sc_hd__o211a_1
XANTENNA__07941__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ top0.MMIO.WBData_i\[13\] net138 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__or2_1
X_07762_ _03881_ _03947_ _04112_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09143__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06713_ top0.CPU.register.registers\[516\] top0.CPU.register.registers\[548\] top0.CPU.register.registers\[580\]
+ top0.CPU.register.registers\[612\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03370_
+ sky130_fd_sc_hd__mux4_1
X_07693_ net485 _03924_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__nand2_1
X_09432_ top0.MMIO.WBData_i\[12\] net145 _05028_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__o21a_1
XANTENNA__06052__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06644_ net859 _03300_ _03293_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__o21ai_1
X_09363_ net2561 _04601_ net608 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
X_06575_ _03228_ _03231_ net864 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__mux2_1
XANTENNA__05731__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07422__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ net2867 net170 net416 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__mux2_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09294_ net2227 _04949_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.load2Ct_n\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06355__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ net224 net671 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout410_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ net510 net195 net622 net427 net2373 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout508_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07127_ _03720_ _03736_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08957__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07808__D _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05866__S0 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ net544 _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__nor2_1
X_06009_ _02665_ net579 top0.CPU.control.funct7\[2\] _02518_ vssd1 vssd1 vccd1 vccd1
+ _02666_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268__920 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__inv_2
XFILLER_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309__961 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__inv_2
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09134__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06291__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06043__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06499__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982__634 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__inv_2
XANTENNA__08428__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ clknet_leaf_66_clk _02276_ net1104 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06594__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06456__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_26_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ clknet_leaf_75_clk _00002_ net1124 vssd1 vssd1 vccd1 vccd1 top0.wishbone0.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07999__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ net1215 _01162_ net1017 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11454_ clknet_leaf_67_clk _01102_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09259__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08948__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ clknet_leaf_86_clk _01033_ net1115 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10336_ net2232 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
X_10267_ net144 _05148_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_12006_ net1698 _01645_ net1122 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07923__A1 top0.CPU.intMem_out\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__B2 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ _04912_ net129 net122 net3145 net115 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a221o_1
XFILLER_78_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__09125__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06282__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05934__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06034__S0 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10286__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061__713 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__inv_2
XFILLER_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06360_ top0.CPU.register.registers\[158\] top0.CPU.register.registers\[190\] top0.CPU.register.registers\[222\]
+ top0.CPU.register.registers\[254\] net853 net815 vssd1 vssd1 vccd1 vccd1 _03017_
+ sky130_fd_sc_hd__mux4_1
XFILLER_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08651__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102__754 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__inv_2
X_06291_ top0.CPU.register.registers\[795\] top0.CPU.register.registers\[827\] top0.CPU.register.registers\[859\]
+ top0.CPU.register.registers\[891\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02948_
+ sky130_fd_sc_hd__mux4_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
X_08030_ net205 net705 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__and2_1
Xhold803 top0.CPU.register.registers\[88\] vssd1 vssd1 vccd1 vccd1 net3025 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08939__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold836 net86 vssd1 vssd1 vccd1 vccd1 net3058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 top0.CPU.register.registers\[124\] vssd1 vssd1 vccd1 vccd1 net3047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 top0.CPU.register.registers\[184\] vssd1 vssd1 vccd1 vccd1 net3036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ net589 _04500_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a21o_1
Xhold869 top0.CPU.register.registers\[276\] vssd1 vssd1 vccd1 vccd1 net3091 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold858 top0.CPU.register.registers\[413\] vssd1 vssd1 vccd1 vccd1 net3080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 top0.CPU.register.registers\[206\] vssd1 vssd1 vccd1 vccd1 net3069 sky130_fd_sc_hd__dlygate4sd3_1
X_08932_ _04649_ net560 _04776_ net266 net3315 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__a32o_1
XANTENNA__07925__B _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10383__35 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__inv_2
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08863_ net155 net3155 net354 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__mux2_1
X_07814_ _04458_ _04470_ net544 vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o21ai_1
X_08794_ net162 net680 net310 net290 net2597 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a32o_1
XANTENNA__06273__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966__618 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__inv_2
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07745_ _03582_ _03620_ _03716_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__o21a_1
XANTENNA__07390__A2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09415_ top0.MMIO.WBData_i\[6\] _04933_ net143 top0.MISOtoMMIO\[6\] _05014_ vssd1
+ vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__o221a_1
X_10710__362 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__inv_2
XANTENNA__06576__S1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _03795_ _03819_ net346 vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06627_ net478 net471 net463 net542 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a31o_1
X_09346_ top0.CPU.internalMem.storeCt\[2\] _04993_ vssd1 vssd1 vccd1 vccd1 _04994_
+ sky130_fd_sc_hd__nor2_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06558_ _03213_ _03214_ net869 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
X_09277_ _04934_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06489_ top0.CPU.register.registers\[149\] top0.CPU.register.registers\[181\] top0.CPU.register.registers\[213\]
+ top0.CPU.register.registers\[245\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03146_
+ sky130_fd_sc_hd__mux4_1
X_08228_ net509 net184 net685 net424 net2572 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a32o_1
XANTENNA__08642__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__C _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout994_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08159_ net152 net614 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__and2_1
XFILLER_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08711__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ top0.display.delayctr\[19\] _05583_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10052_ net3411 net667 net602 _05535_ _05137_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a221o_1
XFILLER_130_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06231__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05916__B1 _02571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08881__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ clknet_leaf_73_clk _02259_ net1127 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06892__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08094__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12555_ clknet_4_12_0_clk _02194_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06319__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09291__C1 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ clknet_leaf_83_clk net3160 net1110 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06644__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08633__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ net2178 _02125_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[979\]
+ sky130_fd_sc_hd__dfrtp_1
X_11437_ clknet_leaf_60_clk _01085_ net1100 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10319_ net2249 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653__305 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__inv_2
XFILLER_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05860_ top0.CPU.Op\[5\] net629 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__nand2_2
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06255__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05791_ top0.CPU.Op\[5\] _02339_ _02340_ _02372_ vssd1 vssd1 vccd1 vccd1 _02448_
+ sky130_fd_sc_hd__and4_4
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06007__S0 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07530_ _02790_ _03443_ _04155_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__and3b_1
XANTENNA__07480__B _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07461_ _03878_ _03933_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__or2_1
XANTENNA__08872__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09200_ top0.CPU.internalMem.prev_busy_o _04861_ vssd1 vssd1 vccd1 vccd1 _04862_
+ sky130_fd_sc_hd__and2_1
X_07392_ _02716_ net524 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06412_ top0.CPU.register.registers\[28\] top0.CPU.register.registers\[60\] top0.CPU.register.registers\[92\]
+ top0.CPU.register.registers\[124\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03069_
+ sky130_fd_sc_hd__mux4_1
X_09131_ top0.CPU.register.registers\[72\] net570 net217 net684 net557 vssd1 vssd1
+ vccd1 vccd1 _04837_ sky130_fd_sc_hd__o2111a_1
X_06343_ net780 _02995_ _02997_ _02999_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_20_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10428__80 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__inv_2
X_09062_ _04680_ net552 _04814_ net255 net3071 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__a32o_1
XANTENNA__06635__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06316__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06274_ _02929_ _02930_ net724 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__mux2_1
X_08013_ net512 net150 net709 net439 net2343 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_96_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold600 top0.CPU.intMemAddr\[15\] vssd1 vssd1 vccd1 vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold611 top0.CPU.register.registers\[942\] vssd1 vssd1 vccd1 vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 top0.CPU.register.registers\[371\] vssd1 vssd1 vccd1 vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 top0.CPU.register.registers\[42\] vssd1 vssd1 vccd1 vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 top0.CPU.intMemAddr\[18\] vssd1 vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 top0.CPU.register.registers\[84\] vssd1 vssd1 vccd1 vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 top0.CPU.register.registers\[829\] vssd1 vssd1 vccd1 vccd1 net2910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 top0.CPU.register.registers\[764\] vssd1 vssd1 vccd1 vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 top0.CPU.register.registers\[853\] vssd1 vssd1 vccd1 vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1115_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ net235 _05455_ _05456_ _05454_ net645 vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__o311a_1
Xhold699 top0.CPU.register.registers\[891\] vssd1 vssd1 vccd1 vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
X_08915_ _04732_ net949 net710 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__or3b_4
XANTENNA_fanout575_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ _05387_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__xor2_1
X_11230__882 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__inv_2
XFILLER_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06986__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06246__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ net222 net3170 net353 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__mux2_1
XANTENNA__08560__A1 _04498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _04701_ net328 net292 net2525 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05989_ top0.CPU.register.registers\[133\] top0.CPU.register.registers\[165\] top0.CPU.register.registers\[197\]
+ top0.CPU.register.registers\[229\] net849 net814 vssd1 vssd1 vccd1 vccd1 _02646_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout742_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _02944_ net520 net446 _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__o31a_1
XANTENNA__06549__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ _04087_ _04310_ _04315_ _04309_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_105_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09329_ _04601_ _04977_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and2_1
XFILLER_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08706__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12340_ net2032 _01979_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[833\]
+ sky130_fd_sc_hd__dfrtp_1
X_12271_ net1963 _01910_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[764\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08441__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05918__X _02575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ top0.display.delayctr\[16\] _05569_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__or2_1
X_10035_ net589 _04475_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a21o_1
XANTENNA__06237__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10988__640 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__inv_2
XANTENNA__07581__A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ net1678 _01625_ net1053 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08303__A1 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ clknet_leaf_81_clk _02242_ net1112 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08606__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12538_ clknet_leaf_77_clk net3378 net1117 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07814__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06093__A2 _02734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06712__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173__825 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__inv_2
X_12469_ net2161 _02108_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[962\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_4
XANTENNA__07475__B _03637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11214__866 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06961_ _03603_ net522 vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nor2_1
X_09680_ top0.CPU.internalMem.pcOut\[3\] net768 vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__or2_1
X_05912_ top0.CPU.register.registers\[2\] top0.CPU.register.registers\[34\] top0.CPU.register.registers\[66\]
+ top0.CPU.register.registers\[98\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02569_
+ sky130_fd_sc_hd__mux4_1
X_08700_ net210 net3040 net357 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06892_ net760 _03546_ net751 vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21o_1
XANTENNA__06002__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06779__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ _04640_ net311 net301 net2686 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__a22o_1
X_05843_ _02498_ _02499_ net730 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XFILLER_82_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05774_ net942 _02413_ _02424_ _02429_ _02375_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a311o_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09098__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ net2886 _04510_ net333 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__mux2_1
X_07513_ net470 _03356_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__and2_1
X_11108__760 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__inv_2
X_08493_ _04694_ net385 net365 net2743 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__a22o_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout156_A _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07444_ _03999_ _04007_ net347 vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__mux2_1
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781__433 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__inv_2
XANTENNA__06951__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout323_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07375_ _03876_ _03880_ net479 vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__mux2_1
XANTENNA__08058__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ top0.CPU.register.registers\[82\] net574 net558 vssd1 vssd1 vccd1 vccd1 _04830_
+ sky130_fd_sc_hd__o21a_1
X_06326_ net580 _02455_ _02980_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a31o_1
X_10822__474 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__inv_2
X_06257_ top0.CPU.register.registers\[537\] top0.CPU.register.registers\[569\] top0.CPU.register.registers\[601\]
+ top0.CPU.register.registers\[633\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02914_
+ sky130_fd_sc_hd__mux4_1
X_09045_ net157 net3199 net349 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__mux2_1
Xhold452 top0.CPU.register.registers\[685\] vssd1 vssd1 vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold463 top0.CPU.register.registers\[903\] vssd1 vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 top0.CPU.register.registers\[123\] vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 top0.CPU.register.registers\[310\] vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ net781 _02844_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__nor2_1
Xhold485 top0.CPU.register.registers\[933\] vssd1 vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold474 top0.CPU.register.registers\[807\] vssd1 vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06467__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold496 top0.CPU.register.registers\[334\] vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout932 net934 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_4
Xfanout943 top0.CPU.control.funct3\[1\] vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_2
X_09947_ _05437_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__and2_1
XANTENNA__06241__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout921 net925 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
Xfanout910 net919 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_2
Xfanout954 top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
Xfanout976 net1004 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout965 net968 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_2
Xhold1141 top0.MMIO.WBData_i\[16\] vssd1 vssd1 vccd1 vccd1 net3363 sky130_fd_sc_hd__dlygate4sd3_1
X_09878_ _05375_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__nand2b_1
Xfanout998 net1000 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1130 top0.CPU.register.registers\[977\] vssd1 vssd1 vccd1 vccd1 net3352 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout987 net988 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_4
Xhold1185 top0.CPU.intMem_out\[27\] vssd1 vssd1 vccd1 vccd1 net3407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1174 top0.display.delayctr\[7\] vssd1 vssd1 vccd1 vccd1 net3396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1163 top0.display.delayctr\[23\] vssd1 vssd1 vccd1 vccd1 net3385 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06729__B _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1152 top0.display.delayctr\[27\] vssd1 vssd1 vccd1 vccd1 net3374 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ net158 net668 net306 net285 net2490 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__a32o_1
X_11840_ net1532 _01479_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[333\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1196 top0.display.delayctr\[18\] vssd1 vssd1 vccd1 vccd1 net3418 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09105__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ net1463 _01410_ net1011 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[264\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06847__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08436__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08049__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157__809 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12323_ net2015 _01962_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[816\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload19 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_11_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09549__A0 top0.CPU.control.funct7\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ net1946 _01893_ net1007 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08221__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ net1877 _01824_ net1000 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[678\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10018_ top0.CPU.internalMem.pcOut\[29\] net649 vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__or2_1
XFILLER_76_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06630__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10765__417 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__inv_2
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08827__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ net1661 _01608_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07250__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806__458 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__inv_2
X_07160_ net526 net527 net468 vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06111_ top0.CPU.control.funct3\[0\] _02474_ _02472_ vssd1 vssd1 vccd1 vccd1 _02768_
+ sky130_fd_sc_hd__a21o_1
X_07091_ net518 _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__nor2_1
XANTENNA__08055__A3 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06042_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__inv_2
XANTENNA__08460__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10659__311 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__inv_2
XANTENNA__06449__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09801_ net587 _02734_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__nor2_1
Xfanout217 _04603_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__D _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 _04533_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlymetal6s2s_1
X_09732_ top0.CPU.internalMem.pcOut\[7\] net650 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__nor2_1
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
X_07993_ top0.CPU.internalMem.pcOut\[3\] net640 net635 _04621_ vssd1 vssd1 vccd1 vccd1
+ _04622_ sky130_fd_sc_hd__o211a_4
XANTENNA_clkload10_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06944_ _03584_ net523 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08515__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ top0.CPU.register.registers\[137\] top0.CPU.register.registers\[169\] top0.CPU.register.registers\[201\]
+ top0.CPU.register.registers\[233\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03532_
+ sky130_fd_sc_hd__mux4_1
X_09663_ net768 _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout273_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ net723 net191 net327 net332 net2508 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a32o_1
XANTENNA__06621__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05826_ net729 _02482_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__and2_1
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _02614_ _05007_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_120_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ net219 net672 net399 net363 net2298 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a32o_1
XANTENNA__08279__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08818__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__B net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05757_ _02338_ _02375_ _02406_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__nor3_1
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout538_A _03073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_128_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11342__994 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__inv_2
X_08476_ net185 net621 net402 net372 net2305 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a32o_1
X_05688_ net860 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07427_ _03740_ _04082_ _04083_ net443 _04081_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__a221o_1
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout705_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ net451 _04011_ _04013_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_118_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08046__A3 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06309_ top0.CPU.register.registers\[796\] top0.CPU.register.registers\[828\] top0.CPU.register.registers\[860\]
+ top0.CPU.register.registers\[892\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02966_
+ sky130_fd_sc_hd__mux4_1
X_07289_ _03723_ _03734_ net481 vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__mux2_1
XANTENNA__06688__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05909__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ net221 net3052 net350 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__mux2_1
XANTENNA__12324__RESET_B net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold260 top0.CPU.register.registers\[804\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 top0.CPU.register.registers\[113\] vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 top0.CPU.intMemAddr\[14\] vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold293 top0.CPU.register.registers\[482\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout740 _02348_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_113_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout751 net755 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_4
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout773 net775 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
Xfanout784 net787 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06860__S0 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout762 net763 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
XFILLER_1_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06612__S0 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10452__104 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__inv_2
XFILLER_46_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11823_ net1515 _01462_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08809__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06746__Y _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11754_ net1446 _01393_ net965 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08285__A3 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ net1377 _01324_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08690__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__X _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload108 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__clkinv_16
Xclkload119 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__inv_6
XANTENNA__07245__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ net1998 _01945_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[799\]
+ sky130_fd_sc_hd__dfrtp_1
X_12237_ net1929 _01876_ net958 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[730\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10001__B1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06205__C1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ net1860 _01807_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[661\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06851__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_12099_ net1791 _01738_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[592\]
+ sky130_fd_sc_hd__dfrtp_1
X_11285__937 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__inv_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_11326__978 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__inv_2
XANTENNA__06603__S0 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ net858 _03316_ _03309_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__o21ai_4
XFILLER_37_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06591_ _02618_ _02651_ net542 vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08276__A3 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08330_ net3075 net409 net387 _04529_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XANTENNA__08681__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06287__A2 _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179__831 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__inv_2
X_08261_ net2990 net418 _04715_ net501 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XFILLER_20_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07212_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__inv_2
X_08192_ net946 _02399_ net688 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__nand3_4
XANTENNA__07236__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07143_ net465 _03799_ _03798_ net477 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o211a_1
XANTENNA__05729__A top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _03729_ _03730_ net459 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__mux2_1
X_10893__545 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__inv_2
X_06025_ _02678_ _02681_ net735 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout390_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _04106_ net232 net227 vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__and3_1
X_10934__586 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__inv_2
XANTENNA__06842__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09715_ _05222_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__xnor2_1
X_06927_ _02926_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ top0.display.counter\[3\] top0.display.counter\[2\] _05123_ top0.display.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__o31a_1
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05970__A1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06858_ top0.CPU.register.registers\[394\] top0.CPU.register.registers\[426\] top0.CPU.register.registers\[458\]
+ top0.CPU.register.registers\[490\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03515_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05751__X _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06994__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_A top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05809_ top0.CPU.register.registers\[147\] top0.CPU.register.registers\[179\] top0.CPU.register.registers\[211\]
+ top0.CPU.register.registers\[243\] net856 net821 vssd1 vssd1 vccd1 vccd1 _02466_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06070__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09577_ net604 _05121_ net3389 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
X_06789_ _02619_ _02686_ _02731_ net540 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ _04713_ net395 net362 net2761 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a22o_1
XANTENNA__06295__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828__480 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__inv_2
XANTENNA__08672__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _04676_ net388 net369 net2617 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11470_ clknet_leaf_69_clk _01118_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct7\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08714__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__A1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10389__41 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__inv_2
XANTENNA__05789__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ _04938_ _05572_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__or2_1
XFILLER_3_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ net1714 _01661_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[515\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05884__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11013__665 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__inv_2
Xfanout592 net593 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_2
XANTENNA__07950__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_4
XANTENNA__09137__D1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11806_ net1498 _01445_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ net1429 _01376_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08663__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ net1360 _01307_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[161\]
+ sky130_fd_sc_hd__dfrtp_1
X_10580__232 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__inv_2
X_11599_ net1291 _01238_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08415__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10877__529 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__inv_2
XANTENNA__07769__A2 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621__273 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07830_ top0.CPU.intMem_out\[30\] net628 _04485_ _02382_ vssd1 vssd1 vccd1 vccd1
+ _04486_ sky130_fd_sc_hd__a211o_1
XFILLER_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07483__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ _03872_ _04087_ _04414_ _03849_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__o221a_1
X_09500_ top0.MMIO.WBData_i\[7\] net140 vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_88_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06712_ top0.CPU.register.registers\[644\] top0.CPU.register.registers\[676\] top0.CPU.register.registers\[708\]
+ top0.CPU.register.registers\[740\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03369_
+ sky130_fd_sc_hd__mux4_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07692_ _03736_ net245 _04155_ net442 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__o22a_1
X_09431_ net3399 net598 net130 _05031_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__o22a_1
XANTENNA__06052__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06643_ _03296_ _03299_ net749 vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__mux2_1
X_09362_ net2957 _04604_ net610 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
X_06574_ _03229_ _03230_ net871 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__mux2_1
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08313_ net2690 net174 net415 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__mux2_1
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08654__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _02367_ _04853_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout236_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net3038 net419 _04707_ net513 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08406__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08175_ net2966 net426 _04686_ net502 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ net452 _03757_ _03782_ _03753_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__o211a_1
XANTENNA__08709__A1 _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05866__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07057_ _02432_ _03713_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__nor2_1
X_06008_ net741 _02664_ _02659_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout772_A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06815__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06196__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ top0.CPU.intMem_out\[10\] net628 _04588_ _04594_ vssd1 vssd1 vccd1 vccd1
+ _04595_ sky130_fd_sc_hd__a22o_1
XFILLER_56_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06291__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07145__A0 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ net3255 net605 net659 net3094 _05159_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__a221o_1
XFILLER_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ clknet_leaf_66_clk _02275_ net1103 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07448__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06229__S net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11432__Q top0.CPU.intMem_out\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
X_12571_ clknet_leaf_75_clk _00001_ net1124 vssd1 vssd1 vccd1 vccd1 top0.wishbone0.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10564__216 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__inv_2
XANTENNA__08645__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08444__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ net1214 _01161_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07999__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11453_ clknet_leaf_70_clk _01101_ net1120 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_10605__257 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11384_ clknet_leaf_78_clk _01032_ net1107 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09070__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10335_ net2254 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10266_ net3015 net119 net112 _05655_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a22o_1
X_10458__110 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__inv_2
X_12005_ net1697 _01644_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[498\]
+ sky130_fd_sc_hd__dfrtp_1
X_10197_ _04915_ net129 net121 net3097 net115 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a221o_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07384__B1 _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06282__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05934__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07136__A0 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06034__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06139__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ net61 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_41_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08636__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06111__A1 top0.CPU.control.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141__793 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__inv_2
X_06290_ top0.CPU.register.registers\[923\] top0.CPU.register.registers\[955\] top0.CPU.register.registers\[987\]
+ top0.CPU.register.registers\[1019\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02947_
+ sky130_fd_sc_hd__mux4_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08651__A3 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07478__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06382__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold826 top0.CPU.register.registers\[543\] vssd1 vssd1 vccd1 vccd1 net3048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 top0.CPU.register.registers\[1011\] vssd1 vssd1 vccd1 vccd1 net3059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__A3 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold815 top0.CPU.register.registers\[406\] vssd1 vssd1 vccd1 vccd1 net3037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold804 top0.CPU.register.registers\[469\] vssd1 vssd1 vccd1 vccd1 net3026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold859 top0.CPU.register.registers\[171\] vssd1 vssd1 vccd1 vccd1 net3081 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ net589 _02946_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__nor2_1
Xmax_cap578 _02430_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
Xhold848 top0.CPU.register.registers\[661\] vssd1 vssd1 vccd1 vccd1 net3070 sky130_fd_sc_hd__dlygate4sd3_1
X_08931_ top0.CPU.register.registers\[211\] net575 vssd1 vssd1 vccd1 vccd1 _04776_
+ sky130_fd_sc_hd__or2_1
X_08862_ net158 net3271 net353 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__mux2_1
X_07813_ _03701_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__and2b_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_123_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06273__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08793_ net165 net681 net311 net289 net2354 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a32o_1
X_07744_ _03582_ _03620_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__nand2_1
XANTENNA__05742__A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _03223_ _03941_ _03244_ _03198_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o211a_1
XANTENNA__07678__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09414_ net2980 _04949_ _05020_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout353_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06626_ net470 net462 net542 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05784__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09345_ top0.CPU.internalMem.storeCt\[0\] top0.CPU.internalMem.storeCt\[1\] vssd1
+ vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_32_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06557_ top0.CPU.register.registers\[401\] top0.CPU.register.registers\[433\] top0.CPU.register.registers\[465\]
+ top0.CPU.register.registers\[497\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03214_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout520_A _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09276_ _04932_ net577 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__or2_4
X_06488_ _03143_ _03144_ net870 vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__mux2_1
X_10899__551 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__inv_2
XANTENNA__07850__A1 top0.CPU.intMem_out\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08227_ net506 net188 net683 net423 net2274 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10198__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09052__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08158_ net2971 net426 _04679_ net500 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a22o_1
X_10359__11 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__inv_2
X_08089_ net505 net199 net694 net434 net2277 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a32o_1
XANTENNA__07602__A1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ net534 net535 net473 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__mux2_1
XANTENNA__07602__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__C1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ top0.display.delayctr\[19\] _05583_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _05533_ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08158__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_128_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11427__Q top0.CPU.intMem_out\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05916__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084__736 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__inv_2
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08439__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07669__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125__777 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08618__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_65_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12623_ clknet_leaf_98_clk _02258_ net1077 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08094__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ clknet_leaf_62_clk _02193_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ clknet_leaf_84_clk net3294 net1110 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12485_ net2177 _02124_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[978\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11436_ clknet_leaf_67_clk _01084_ net1101 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09043__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ top0.CPU.internalMem.storeCt\[2\] _05674_ _05675_ _05677_ vssd1 vssd1 vccd1
+ vccd1 _02335_ sky130_fd_sc_hd__a22o_1
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11019__671 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__inv_2
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10249_ net22 net653 net592 top0.MMIO.WBData_i\[28\] vssd1 vssd1 vccd1 vccd1 _02295_
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10692__344 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__inv_2
XANTENNA__06255__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05790_ _02340_ _02378_ _02381_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__or3_4
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07109__A0 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733__385 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__inv_2
XANTENNA__06007__S1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07253__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07460_ _04076_ _04116_ net458 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__mux2_1
X_07391_ _02716_ _03556_ net444 _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__o31a_1
X_06411_ top0.CPU.register.registers\[156\] top0.CPU.register.registers\[188\] top0.CPU.register.registers\[220\]
+ top0.CPU.register.registers\[252\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03068_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08609__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ net179 net685 net278 net253 net2428 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a32o_1
XANTENNA__08592__B _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06342_ net732 _02998_ net739 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_14_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_20_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ top0.CPU.register.registers\[119\] net564 vssd1 vssd1 vccd1 vccd1 _04814_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ net946 _02399_ net710 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand3_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06273_ top0.CPU.register.registers\[538\] top0.CPU.register.registers\[570\] top0.CPU.register.registers\[602\]
+ top0.CPU.register.registers\[634\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02930_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09034__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold601 top0.CPU.register.registers\[604\] vssd1 vssd1 vccd1 vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
X_10443__95 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__inv_2
Xhold612 top0.CPU.register.registers\[662\] vssd1 vssd1 vccd1 vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 top0.CPU.register.registers\[588\] vssd1 vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 top0.CPU.register.registers\[773\] vssd1 vssd1 vccd1 vccd1 net2867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 top0.CPU.register.registers\[177\] vssd1 vssd1 vccd1 vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 top0.CPU.register.registers\[798\] vssd1 vssd1 vccd1 vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05737__A top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ top0.CPU.internalMem.pcOut\[24\] _05426_ top0.CPU.internalMem.pcOut\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a21oi_1
Xhold656 top0.CPU.register.registers\[902\] vssd1 vssd1 vccd1 vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 top0.CPU.register.registers\[1016\] vssd1 vssd1 vccd1 vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xhold689 top0.CPU.register.registers\[128\] vssd1 vssd1 vccd1 vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ net717 net156 net273 _04753_ net2383 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1010_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ _05345_ _05391_ _05390_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1108_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07952__A _03989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ _04555_ net3331 net355 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__mux2_1
XANTENNA__06246__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05743__Y _02400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _04700_ net321 net291 net2546 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout568_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05988_ top0.CPU.register.registers\[389\] top0.CPU.register.registers\[421\] top0.CPU.register.registers\[453\]
+ top0.CPU.register.registers\[485\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02645_
+ sky130_fd_sc_hd__mux4_1
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__A1_N _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07727_ _02944_ _03656_ net341 vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_28_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ _03720_ _04219_ _04311_ _04056_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06609_ top0.CPU.register.registers\[645\] top0.CPU.register.registers\[677\] top0.CPU.register.registers\[709\]
+ top0.CPU.register.registers\[741\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03266_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_105_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09231__X _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ _03907_ _03933_ _04244_ _04245_ _04050_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__o221a_1
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
X_09328_ _04016_ _04044_ net232 net227 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__and4_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08615__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06343__A1_N net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ top0.CPU.intMemAddr\[8\] _04601_ net770 vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__mux2_1
XANTENNA__06182__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08722__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12270_ net1962 _01909_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[763\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08379__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676__328 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ _04957_ _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__or2_1
XANTENNA__08958__A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10717__369 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__inv_2
X_10034_ net589 _03686_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__nor2_1
XANTENNA__06237__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05996__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ net1677 _01624_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12606_ clknet_leaf_81_clk _02241_ net1112 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08067__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12537_ clknet_leaf_77_clk net3416 net1117 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12468_ net2160 _02107_ net961 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[961\]
+ sky130_fd_sc_hd__dfrtp_1
X_11419_ clknet_leaf_69_clk _01067_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12399_ net2091 _02038_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08790__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ net746 _03616_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__o2bb2a_2
Xclkbuf_leaf_3_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_06891_ net871 _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__and2_1
X_05911_ top0.CPU.register.registers\[130\] top0.CPU.register.registers\[162\] top0.CPU.register.registers\[194\]
+ top0.CPU.register.registers\[226\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02568_
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05842_ top0.CPU.register.registers\[527\] top0.CPU.register.registers\[559\] top0.CPU.register.registers\[591\]
+ top0.CPU.register.registers\[623\] net851 net816 vssd1 vssd1 vccd1 vccd1 _02499_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08542__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ _04639_ net317 net302 net2749 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__a22o_1
XANTENNA__05987__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05773_ net942 _02413_ _02424_ _02429_ _02375_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a311oi_4
X_08561_ net3013 _04504_ net333 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XANTENNA__06305__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07512_ net487 net531 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__xnor2_1
X_08492_ _04693_ net388 net365 net2934 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__a22o_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07443_ _03816_ _04087_ _04095_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__o211a_1
XANTENNA__08058__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ _04701_ net560 _04829_ net254 net3261 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a32o_1
XANTENNA__08108__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ net449 _04030_ _04022_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o21a_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_33_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06325_ net775 _02978_ _02970_ net584 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09007__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11395__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ net160 net3317 net350 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__mux2_1
X_06256_ top0.CPU.register.registers\[665\] top0.CPU.register.registers\[697\] top0.CPU.register.registers\[729\]
+ top0.CPU.register.registers\[761\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02913_
+ sky130_fd_sc_hd__mux4_1
XFILLER_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold420 top0.CPU.register.registers\[450\] vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05911__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold453 top0.CPU.register.registers\[582\] vssd1 vssd1 vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 top0.CPU.register.registers\[474\] vssd1 vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ _02842_ _02843_ net731 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__mux2_1
Xhold431 top0.CPU.register.registers\[802\] vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net904 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__buf_2
Xhold486 net40 vssd1 vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06467__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold464 top0.CPU.register.registers\[476\] vssd1 vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 top0.CPU.register.registers\[590\] vssd1 vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08781__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_4
Xhold497 top0.CPU.register.registers\[589\] vssd1 vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09946_ top0.CPU.internalMem.pcOut\[24\] _05438_ vssd1 vssd1 vccd1 vccd1 _05440_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06997__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout911 net913 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_4
Xfanout922 net925 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_4
Xfanout955 top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_1
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_2
XFILLER_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout977 net982 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout852_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ net587 _04546_ _05373_ top0.CPU.internalMem.pcOut\[19\] vssd1 vssd1 vccd1
+ vccd1 _05376_ sky130_fd_sc_hd__a211o_1
Xhold1142 net64 vssd1 vssd1 vccd1 vccd1 net3364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold1120 top0.CPU.register.registers\[75\] vssd1 vssd1 vccd1 vccd1 net3342 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
Xhold1131 top0.CPU.register.registers\[230\] vssd1 vssd1 vccd1 vccd1 net3353 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout988 net995 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_2
Xhold1153 top0.CPU.intMem_out\[18\] vssd1 vssd1 vccd1 vccd1 net3375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 top0.CPU.intMem_out\[8\] vssd1 vssd1 vccd1 vccd1 net3397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 top0.CPU.intMem_out\[2\] vssd1 vssd1 vccd1 vccd1 net3386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08828_ net162 net669 net309 net286 net2362 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__a32o_1
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1186 top0.CPU.intMem_out\[10\] vssd1 vssd1 vccd1 vccd1 net3408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1197 top0.display.delayctr\[6\] vssd1 vssd1 vccd1 vccd1 net3419 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ net213 net615 net309 net293 net2456 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__a32o_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09089__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11770_ net1462 _01409_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[263\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08049__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196__848 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11440__Q top0.CPU.intMem_out\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12322_ net2014 _01961_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05807__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08452__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net1945 _01892_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[746\]
+ sky130_fd_sc_hd__dfrtp_1
X_11237__889 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__inv_2
XANTENNA__05902__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10283__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ net1876 _01823_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08772__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ _05504_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XANTENNA__08524__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06630__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11968_ net1660 _01607_ net1035 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[461\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ net1591 _01538_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06394__S0 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10177__B _03020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06147__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10845__497 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__inv_2
XANTENNA__09966__B _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06146__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05986__S net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06110_ _02422_ _02758_ _02766_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__nor3_1
X_07090_ _02428_ net578 _03712_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_93_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06041_ top0.CPU.control.funct7\[4\] _02518_ _02697_ net581 vssd1 vssd1 vccd1 vccd1
+ _02698_ sky130_fd_sc_hd__a22o_2
XANTENNA__06671__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413__65 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__inv_2
X_10698__350 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__inv_2
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06449__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ net631 _04578_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__nor2_1
Xfanout218 _04603_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dlymetal6s2s_1
X_07992_ top0.CPU.intMem_out\[3\] net629 _04588_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_
+ sky130_fd_sc_hd__a22o_1
Xfanout229 _04473_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08763__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 _04522_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
X_10739__391 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__inv_2
X_09731_ net237 _05240_ _05241_ _05238_ _05239_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__o32a_1
XFILLER_86_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06943_ net745 _03599_ _03591_ _03592_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08515__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05734__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06874_ _03527_ _03530_ net751 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
X_09662_ _02558_ _04623_ net590 vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__mux2_1
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06621__S1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ net718 net193 net324 net331 net2464 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a32o_1
X_05825_ top0.CPU.register.registers\[530\] top0.CPU.register.registers\[562\] top0.CPU.register.registers\[594\]
+ top0.CPU.register.registers\[626\] net846 net811 vssd1 vssd1 vccd1 vccd1 _02482_
+ sky130_fd_sc_hd__mux4_1
X_09593_ net2850 net658 _05132_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout266_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ net181 net674 net401 net364 net2309 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a32o_1
XFILLER_82_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05756_ top0.CPU.control.funct7\[1\] top0.CPU.control.funct7\[0\] top0.CPU.control.funct7\[5\]
+ _02410_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__or4_2
XANTENNA__08279__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08818__A3 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05750__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05687_ net864 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__inv_2
XANTENNA__08684__D1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ net187 net619 net398 net371 net2485 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout433_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06385__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06057__S net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ _02666_ _03262_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09779__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ _03742_ _03997_ _04001_ _03992_ net452 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_118_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06308_ _02963_ _02964_ net726 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__mux2_1
XANTENNA__06137__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09027_ _04571_ net3205 net351 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__mux2_1
XANTENNA__06581__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ _03731_ _03767_ net480 vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06239_ net786 _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold261 top0.CPU.register.registers\[1023\] vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__B1 _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 top0.CPU.register.registers\[931\] vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 top0.CPU.register.registers\[296\] vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top0.CPU.register.registers\[420\] vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 top0.CPU.register.registers\[416\] vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout730 _02349_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 net742 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout785 net787 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_2
Xfanout752 net755 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_2
Xfanout774 net775 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08506__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__S1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _05422_ _05423_ net238 vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a21oi_1
Xfanout763 _02344_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_4
X_10491__143 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__inv_2
Xfanout796 net799 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_2
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08020__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06612__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__Q top0.CPU.intMem_out\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_47_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ net1514 _01461_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[315\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08447__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532__184 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06376__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06475__B _03130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ net1445 _01392_ net1070 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[246\]
+ sky130_fd_sc_hd__dfrtp_1
X_11684_ net1376 _01323_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[177\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload109 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__inv_4
XANTENNA__06128__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ net1997 _01944_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08993__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12236_ net1928 _01875_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08745__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ net1859 _01806_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[660\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06300__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06851__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ net1790 _01737_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[591\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06508__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09170__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06603__S1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09458__B1 _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06590_ net477 net471 net462 net542 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__a31o_1
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06367__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _04539_ net671 vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__and2_1
X_08191_ net955 net951 net953 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__or3b_1
X_07211_ _03763_ _03777_ net465 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__mux2_1
X_07142_ net521 net538 net475 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__mux2_1
XANTENNA__07236__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08984__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ net528 net529 net467 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__mux2_1
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06024_ _02679_ _02680_ net725 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XANTENNA__09933__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06842__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ net714 net498 net177 net546 net2463 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a32o_1
X_10475__127 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__inv_2
XFILLER_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09714_ _05189_ _05202_ _05223_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__o31a_1
X_06926_ _02457_ net242 _02908_ net544 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a31o_1
X_06857_ top0.CPU.register.registers\[10\] top0.CPU.register.registers\[42\] top0.CPU.register.registers\[74\]
+ top0.CPU.register.registers\[106\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03514_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09651__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ top0.display.dataforOutput\[14\] net605 net659 net3159 _05170_ vssd1 vssd1
+ vccd1 vccd1 _01145_ sky130_fd_sc_hd__a221o_1
X_05808_ net781 _02460_ _02463_ _02464_ net774 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout648_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06847__Y _03504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10516__168 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__inv_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ top0.display.state\[0\] net666 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__nand2_1
X_06788_ _03429_ net528 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06358__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05739_ net571 net633 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__and2_4
X_08527_ _04712_ net387 net361 net2625 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a22o_1
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ _04675_ net393 net369 net2828 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a22o_1
XANTENNA__06683__B1 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ net488 _04065_ _03841_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__a21o_1
XFILLER_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ _04654_ net405 net379 net2553 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06515__S net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08424__A1 _04492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06530__S0 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10282_ net3065 net121 net113 _05662_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09924__A1 top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08188__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net1713 _01660_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[514\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06738__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _04754_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_4
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_1
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout571 net574 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_2
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_2
XANTENNA__09137__C1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06597__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08360__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11805_ net1497 _01444_ net1024 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[298\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ net1428 _01375_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07871__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ net1359 _01306_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[160\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252__904 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__inv_2
XANTENNA__09612__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08206__A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ net1290 _01237_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10222__B2 top0.MMIO.WBData_i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08966__A2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06521__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08179__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ net1911 _01858_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05836__Y _02493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07760_ net451 _04118_ _04144_ _03752_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_88_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06711_ _03366_ _03367_ net757 vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__mux2_1
XANTENNA__09143__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ top0.MMIO.WBData_i\[11\] net146 _05028_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__o21a_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07691_ _02514_ _03425_ net445 _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__o31a_1
XANTENNA__08351__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06642_ _03297_ _03298_ net757 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__mux2_1
XFILLER_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ net2885 _04608_ net610 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
XFILLER_80_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06573_ top0.CPU.register.registers\[912\] top0.CPU.register.registers\[944\] top0.CPU.register.registers\[976\]
+ top0.CPU.register.registers\[1008\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03230_
+ sky130_fd_sc_hd__mux4_1
XFILLER_52_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ _02367_ _04853_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__nor2_1
X_08312_ net2959 net177 net415 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__mux2_1
XANTENNA__08103__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ net212 net675 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__and2_1
X_10860__512 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__inv_2
XFILLER_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08174_ net221 net617 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_99_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901__553 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__inv_2
XANTENNA__08957__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ net485 _03768_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a21o_1
XANTENNA__06512__S0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1040_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _02423_ _03712_ _02416_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__nand3b_2
X_06007_ _02660_ _02661_ _02662_ _02663_ net725 net776 vssd1 vssd1 vccd1 vccd1 _02664_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11036__688 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__inv_2
XANTENNA__06815__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08185__A3 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ net562 _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__or2_1
XANTENNA__09134__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06579__S0 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ net591 _02851_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nand2_1
XANTENNA__08342__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ _03411_ net529 _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__o21a_1
XFILLER_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07145__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ net141 _05158_ _04955_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ net945 _02408_ _04217_ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a31o_1
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12570_ clknet_leaf_75_clk _00000_ net1124 vssd1 vssd1 vccd1 vccd1 top0.wishbone0.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_26_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08725__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ net1213 _01160_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ clknet_leaf_66_clk _01100_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire246 _02732_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08026__A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ clknet_leaf_79_clk _01031_ net1114 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08948__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10644__296 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__inv_2
X_10334_ net2239 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09556__S _04175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07620__A2 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10265_ net144 _05146_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__nand2_1
XANTENNA__10291__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__A3 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _04920_ net129 net122 net3364 net115 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a221o_1
X_12004_ net1696 _01643_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07384__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10538__190 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__inv_2
XANTENNA__07136__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__B _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10140__B1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload7_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ net61 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_12699_ clknet_leaf_75_clk _02334_ net1124 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.storeCt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08100__A3 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ net1411 _01358_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[212\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08939__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold827 top0.CPU.register.registers\[650\] vssd1 vssd1 vccd1 vccd1 net3049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 top0.CPU.register.registers\[830\] vssd1 vssd1 vccd1 vccd1 net3038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold805 net87 vssd1 vssd1 vccd1 vccd1 net3027 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__A0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold838 top0.CPU.register.registers\[549\] vssd1 vssd1 vccd1 vccd1 net3060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 top0.CPU.register.registers\[119\] vssd1 vssd1 vccd1 vccd1 net3071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _04648_ net272 net263 net2557 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__a22o_1
XFILLER_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ net162 net2988 net353 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__mux2_1
X_07812_ _03785_ _04468_ net519 vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__nor3b_1
XANTENNA__06583__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08792_ net213 net680 net309 net289 net2695 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__a32o_1
XANTENNA__09116__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ _03715_ _04390_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07127__A1 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ net343 _04322_ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a21o_1
XANTENNA__07678__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06335__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ top0.MMIO.WBData_i\[5\] _04933_ _04953_ top0.MISOtoMMIO\[5\] _05014_ vssd1
+ vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__o221a_1
X_06625_ _03280_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nand2b_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587__239 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__inv_2
XANTENNA_fanout346_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05784__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _04950_ _04986_ _04989_ _04992_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.state_n\[0\]
+ sky130_fd_sc_hd__or4_1
X_06556_ top0.CPU.register.registers\[273\] top0.CPU.register.registers\[305\] top0.CPU.register.registers\[337\]
+ top0.CPU.register.registers\[369\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03213_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_23_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ net577 _04930_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__and2b_1
XANTENNA__07835__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06487_ top0.CPU.register.registers\[405\] top0.CPU.register.registers\[437\] top0.CPU.register.registers\[469\]
+ top0.CPU.register.registers\[501\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03144_
+ sky130_fd_sc_hd__mux4_1
X_08226_ net515 net190 net688 net424 net2269 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a32o_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ net207 net617 vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07108_ net533 _03221_ net473 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout882_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ net2815 net435 _04666_ net495 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22o_1
X_07039_ top0.CPU.register.registers\[31\] top0.CPU.register.registers\[63\] top0.CPU.register.registers\[95\]
+ top0.CPU.register.registers\[127\] net852 net816 vssd1 vssd1 vccd1 vccd1 _03696_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10050_ top0.display.delayctr\[0\] top0.display.delayctr\[1\] top0.display.delayctr\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__o21ai_1
X_10374__26 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08012__C net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05916__A2 _02563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09107__A2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05933__A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06748__B _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06972__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12622_ clknet_leaf_81_clk _02257_ net1109 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ clknet_leaf_62_clk _02192_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_11504_ clknet_leaf_84_clk _01143_ net1107 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12484_ net2176 _02123_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[977\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ clknet_leaf_69_clk _01083_ net1100 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ top0.CPU.internalMem.storeCt\[2\] _05676_ vssd1 vssd1 vccd1 vccd1 _05677_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10248_ net21 net653 net592 top0.MMIO.WBData_i\[27\] vssd1 vssd1 vccd1 vccd1 _02294_
+ sky130_fd_sc_hd__o22a_1
Xfanout1130 net1131 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10179_ top0.display.delayctr\[30\] _05630_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07109__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__B1 _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06410_ net750 _03062_ net859 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__o21ai_1
X_07390_ _02716_ net524 net339 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a21o_1
X_11258__910 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__inv_2
XANTENNA__08085__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06341_ top0.CPU.register.registers\[285\] top0.CPU.register.registers\[317\] top0.CPU.register.registers\[349\]
+ top0.CPU.register.registers\[381\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02998_
+ sky130_fd_sc_hd__mux4_1
X_09060_ _04679_ net555 _04813_ net256 net3263 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__a32o_1
X_06272_ top0.CPU.register.registers\[666\] top0.CPU.register.registers\[698\] top0.CPU.register.registers\[730\]
+ top0.CPU.register.registers\[762\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02929_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_20_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07293__A0 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08011_ net954 net950 net952 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__and3b_1
XFILLER_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold602 top0.CPU.register.registers\[315\] vssd1 vssd1 vccd1 vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__A3 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 top0.CPU.register.registers\[522\] vssd1 vssd1 vccd1 vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 top0.CPU.register.registers\[692\] vssd1 vssd1 vccd1 vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 top0.CPU.register.registers\[828\] vssd1 vssd1 vccd1 vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 top0.CPU.register.registers\[691\] vssd1 vssd1 vccd1 vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 top0.display.counter\[1\] vssd1 vssd1 vccd1 vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ top0.CPU.internalMem.pcOut\[25\] top0.CPU.internalMem.pcOut\[24\] _05426_
+ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__and3_1
XANTENNA__07596__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07596__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972__624 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__inv_2
Xhold657 top0.CPU.register.registers\[471\] vssd1 vssd1 vccd1 vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 top0.CPU.register.registers\[913\] vssd1 vssd1 vccd1 vccd1 net2890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ net713 net157 net267 net282 net2442 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout296_A _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _05353_ _05388_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__and2_1
XANTENNA__08545__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _04550_ net3129 net356 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__mux2_1
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05987_ top0.CPU.register.registers\[261\] top0.CPU.register.registers\[293\] top0.CPU.register.registers\[325\]
+ top0.CPU.register.registers\[357\] net849 net814 vssd1 vssd1 vccd1 vccd1 _02644_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09225__A top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05753__A top0.CPU.control.funct7\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08775_ _04699_ net315 net290 net2722 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _03847_ _03992_ _04382_ net453 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o22a_1
XFILLER_27_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_X net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ _02831_ _03241_ net445 _04312_ _04313_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06608_ _02650_ _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__xnor2_1
X_07588_ net337 _04063_ _04224_ net476 _03743_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a221o_1
XFILLER_25_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _04578_ _04583_ _04870_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__or3_1
X_06539_ _03194_ _03195_ net534 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a21oi_1
X_10419__71 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__inv_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09258_ top0.CPU.internalMem.pcOut\[5\] _04919_ net609 vssd1 vssd1 vccd1 vccd1 _04920_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06182__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09189_ _04851_ _04852_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__or2_1
X_08209_ net3158 net421 _04697_ net491 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
XANTENNA__06523__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08379__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05928__A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051__703 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ _02829_ net550 vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nor2_1
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08958__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__Q top0.CPU.intMem_out\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08536__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _05497_ _05512_ _05514_ _05510_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__o31ai_1
XFILLER_68_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05996__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11984_ net1676 _01623_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[477\]
+ sky130_fd_sc_hd__dfrtp_1
X_12605_ clknet_leaf_92_clk _02240_ net1084 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08067__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12536_ clknet_leaf_74_clk net3380 net1123 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10956__608 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__inv_2
XFILLER_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_12467_ net2159 _02106_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[960\]
+ sky130_fd_sc_hd__dfrtp_1
X_11418_ clknet_leaf_69_clk _01066_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07578__A1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12398_ net2090 _02037_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08775__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700__352 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__inv_2
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06250__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08527__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06890_ top0.CPU.register.registers\[904\] top0.CPU.register.registers\[936\] top0.CPU.register.registers\[968\]
+ top0.CPU.register.registers\[1000\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__mux4_1
XFILLER_67_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05910_ net782 _02564_ net776 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__o21a_1
XFILLER_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05841_ top0.CPU.register.registers\[655\] top0.CPU.register.registers\[687\] top0.CPU.register.registers\[719\]
+ top0.CPU.register.registers\[751\] net851 net816 vssd1 vssd1 vccd1 vccd1 _02498_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08542__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06002__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07491__C _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05987__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05772_ net944 _02408_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__nor2_1
X_08560_ net3197 _04498_ net333 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
X_07511_ net478 _03317_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__xnor2_1
X_08491_ _04692_ net392 net365 net2823 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__a22o_1
X_07442_ _02684_ _03403_ net444 _04097_ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__o311a_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06936__S0 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07373_ _04029_ _04028_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__and2b_1
X_09112_ top0.CPU.register.registers\[83\] net576 vssd1 vssd1 vccd1 vccd1 _04829_
+ sky130_fd_sc_hd__or2_1
X_06324_ _02455_ _02980_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09043_ net164 net613 _04807_ net350 net3283 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout211_A _04498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06255_ top0.CPU.register.registers\[793\] top0.CPU.register.registers\[825\] top0.CPU.register.registers\[857\]
+ top0.CPU.register.registers\[889\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02912_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05748__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__A2 _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 top0.CPU.register.registers\[801\] vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
X_06186_ top0.CPU.register.registers\[21\] top0.CPU.register.registers\[53\] top0.CPU.register.registers\[85\]
+ top0.CPU.register.registers\[117\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02843_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05911__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 top0.CPU.register.registers\[684\] vssd1 vssd1 vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 top0.CPU.register.registers\[435\] vssd1 vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6_0_clk_X clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 top0.CPU.register.registers\[196\] vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 top0.CPU.register.registers\[118\] vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09654__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 top0.CPU.intMemAddr\[16\] vssd1 vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 top0.CPU.register.registers\[694\] vssd1 vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06241__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 top0.CPU.register.registers\[577\] vssd1 vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 top0.CPU.register.registers\[621\] vssd1 vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout934 net938 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
Xfanout901 net903 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_4
XFILLER_104_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07963__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _05438_ top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 _05439_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout580_A _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 net925 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_2
Xfanout912 net913 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_4
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ net631 _04546_ _05374_ top0.CPU.internalMem.pcOut\[19\] vssd1 vssd1 vccd1
+ vccd1 _05375_ sky130_fd_sc_hd__o211a_1
Xfanout945 top0.CPU.control.funct3\[0\] vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_1
Xfanout956 net958 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08518__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
Xhold1110 top0.CPU.register.registers\[368\] vssd1 vssd1 vccd1 vccd1 net3332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 top0.display.dataforOutput\[1\] vssd1 vssd1 vccd1 vccd1 net3354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout978 net982 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_4
X_08827_ net165 net669 net311 net285 net2280 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__a32o_1
Xhold1121 top0.CPU.register.registers\[219\] vssd1 vssd1 vccd1 vccd1 net3343 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net992 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_4
Xhold1165 top0.MISOtoMMIO\[3\] vssd1 vssd1 vccd1 vccd1 net3387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 top0.CPU.intMem_out\[20\] vssd1 vssd1 vccd1 vccd1 net3376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 top0.CPU.control.funct3\[2\] vssd1 vssd1 vccd1 vccd1 net3398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 top0.CPU.register.registers\[301\] vssd1 vssd1 vccd1 vccd1 net3365 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1198 top0.CPU.intMem_out\[22\] vssd1 vssd1 vccd1 vccd1 net3420 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net167 net622 net324 net296 net2334 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__a32o_1
Xhold1187 top0.display.delayctr\[20\] vssd1 vssd1 vccd1 vccd1 net3409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07709_ _03621_ _03659_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__nand2_1
X_08689_ net214 net691 net310 net298 net2516 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_49_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09402__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08018__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05807__A1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12321_ net2013 _01960_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12252_ net1944 _01891_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[745\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05902__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08757__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ net1875 _01822_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[676\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08509__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ top0.CPU.internalMem.pcOut\[29\] _05492_ net238 vssd1 vssd1 vccd1 vccd1 _05505_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_49_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__09182__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11967_ net1659 _01606_ net1097 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05840__B _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11898_ net1590 _01537_ net975 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[391\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06394__S1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06428__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11220__872 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__inv_2
XFILLER_32_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05839__Y _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12519_ net2211 _02158_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1012\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08996__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06146__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06040_ _02691_ _02696_ net743 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_93_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08460__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 _04603_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
X_07991_ net562 _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__or2_1
XANTENNA__08763__A3 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 _04516_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ top0.CPU.internalMem.pcOut\[7\] _05228_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__nor2_1
X_06942_ _03595_ _03598_ net862 vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09173__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ _03528_ _03529_ net760 vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
X_09661_ _02360_ _04857_ net662 _05177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__o31ai_1
XANTENNA__08515__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08920__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06082__S0 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ top0.display.state\[1\] top0.display.state\[0\] top0.display.state\[2\] vssd1
+ vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a21o_1
X_05824_ top0.CPU.register.registers\[658\] top0.CPU.register.registers\[690\] top0.CPU.register.registers\[722\]
+ top0.CPU.register.registers\[754\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02481_
+ sky130_fd_sc_hd__mux4_1
X_08612_ net2893 net330 net316 _04577_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a22o_1
X_08543_ net184 net674 net402 net363 net2644 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a32o_1
X_05755_ net944 _02411_ _02375_ _02342_ net943 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_38_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05750__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08474_ net192 net624 net407 net372 net2401 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_102_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08684__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05686_ net871 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__inv_2
XANTENNA__06338__S net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06385__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07425_ _02666_ _03261_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or2_1
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09649__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07958__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06862__A _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ net490 _03746_ _04010_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a31o_1
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08987__B1 _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07287_ _03196_ _03942_ _03176_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__o21ai_1
X_10978__630 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__inv_2
X_06307_ top0.CPU.register.registers\[540\] top0.CPU.register.registers\[572\] top0.CPU.register.registers\[604\]
+ top0.CPU.register.registers\[636\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02964_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06137__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _04566_ net3165 net351 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__mux2_1
X_06238_ top0.CPU.register.registers\[920\] top0.CPU.register.registers\[952\] top0.CPU.register.registers\[984\]
+ top0.CPU.register.registers\[1016\] net840 net805 vssd1 vssd1 vccd1 vccd1 _02895_
+ sky130_fd_sc_hd__mux4_1
X_11357__1009 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__inv_2
XANTENNA_fanout795_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06169_ top0.CPU.register.registers\[272\] top0.CPU.register.registers\[304\] top0.CPU.register.registers\[336\]
+ top0.CPU.register.registers\[368\] net846 net811 vssd1 vssd1 vccd1 vccd1 _02826_
+ sky130_fd_sc_hd__mux4_1
Xhold251 top0.CPU.register.registers\[432\] vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 top0.CPU.register.registers\[331\] vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 top0.CPU.register.registers\[235\] vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08203__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06801__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 top0.CPU.register.registers\[498\] vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06214__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold273 top0.CPU.register.registers\[484\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 top0.CPU.register.registers\[462\] vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07693__A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout720 net721 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_113_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ _05400_ _05411_ _05413_ _05410_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout742 net744 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
XANTENNA_fanout962_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 top0.CPU.control.rs2\[4\] vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
XANTENNA__09164__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_4
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout786 net787 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08506__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ top0.CPU.internalMem.pcOut\[17\] _05348_ net239 vssd1 vssd1 vccd1 vccd1 _05360_
+ sky130_fd_sc_hd__o21ai_1
Xfanout797 net799 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163__815 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__inv_2
XFILLER_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08728__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11821_ net1513 _01460_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05941__A _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06376__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10278__B _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204__856 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__inv_2
XANTENNA__06248__S net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ net1444 _01391_ net1069 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[245\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11451__Q top0.CPU.decoder.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12774__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ net1375 _01322_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[176\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08690__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08978__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06128__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ net1996 _01943_ net1082 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[797\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08993__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12235_ net1927 _01874_ net1072 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[728\]
+ sky130_fd_sc_hd__dfrtp_1
X_12166_ net1858 _01805_ net1128 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[659\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06205__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06711__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__A0 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771__423 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__inv_2
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06300__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09307__B top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09155__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ net1789 _01736_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[590\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08902__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06064__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10812__464 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__inv_2
XANTENNA__05811__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06367__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09042__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08681__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ net954 net950 net952 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__nor3b_1
XANTENNA__05997__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07210_ net466 _03779_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__or2_1
X_07141_ net475 net539 _03797_ net457 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__a211o_1
XANTENNA__08969__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ net527 _03482_ net468 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__mux2_1
X_06023_ top0.CPU.register.registers\[6\] top0.CPU.register.registers\[38\] top0.CPU.register.registers\[70\]
+ top0.CPU.register.registers\[102\] net831 net795 vssd1 vssd1 vccd1 vccd1 _02680_
+ sky130_fd_sc_hd__mux4_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08197__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ top0.CPU.internalMem.pcOut\[7\] net641 net636 _04606_ vssd1 vssd1 vccd1 vccd1
+ _04607_ sky130_fd_sc_hd__o211a_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07018__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ top0.CPU.internalMem.pcOut\[5\] _05211_ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_
+ sky130_fd_sc_hd__a21oi_1
X_06925_ _03577_ _03578_ _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__and3_1
X_06856_ top0.CPU.register.registers\[138\] top0.CPU.register.registers\[170\] top0.CPU.register.registers\[202\]
+ top0.CPU.register.registers\[234\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03513_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08548__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06055__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ net142 _05169_ net660 vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05807_ net734 _02461_ net739 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a21o_1
XANTENNA__05802__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05761__A top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07452__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09449__A1 top0.MMIO.WBData_i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ top0.display.state\[0\] net666 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__and2_1
X_06787_ _03429_ net528 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08121__A1 _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05738_ top0.CPU.decoder.instruction\[11\] _02393_ vssd1 vssd1 vccd1 vccd1 _02395_
+ sky130_fd_sc_hd__or2_1
XFILLER_51_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08526_ _04711_ net385 net361 net2691 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09520__X _05100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06358__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ _04674_ net397 net370 net2944 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a22o_1
XFILLER_136_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ _04063_ _04064_ net345 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__mux2_1
X_08388_ _04482_ net697 net405 net379 net2576 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a32o_1
X_07339_ _03994_ _03995_ net345 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__mux2_1
X_10350_ net2242 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06530__S1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ _04937_ _05169_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__nand2_1
X_09009_ top0.CPU.register.registers\[156\] net566 vssd1 vssd1 vccd1 vccd1 _04799_
+ sky130_fd_sc_hd__or2_1
XANTENNA__06531__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08188__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ net1712 _01659_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[513\]
+ sky130_fd_sc_hd__dfrtp_1
X_10755__407 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__inv_2
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07935__A1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 net551 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06294__S0 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09137__B1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__Q top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout572 net574 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_4
Xfanout594 _05648_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06046__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06597__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06910__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ net1496 _01443_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[297\]
+ sky130_fd_sc_hd__dfrtp_1
X_10649__301 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__inv_2
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11735_ net1427 _01374_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08663__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ net1358 _01305_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[159\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_14_0_clk_X clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291__943 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__inv_2
XANTENNA__09612__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08206__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11597_ net1289 _01236_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07885__X _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06521__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ net1910 _01857_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[711\]
+ sky130_fd_sc_hd__dfrtp_1
X_11332__984 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__inv_2
XANTENNA__07926__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09037__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net1841 _01788_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09128__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06037__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06710_ top0.CPU.register.registers\[772\] top0.CPU.register.registers\[804\] top0.CPU.register.registers\[836\]
+ top0.CPU.register.registers\[868\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03367_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08876__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _02514_ _03425_ net340 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__a21o_1
X_10354__6 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__inv_2
XFILLER_37_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08351__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06641_ top0.CPU.register.registers\[3\] top0.CPU.register.registers\[35\] top0.CPU.register.registers\[67\]
+ top0.CPU.register.registers\[99\] net916 net882 vssd1 vssd1 vccd1 vccd1 _03298_
+ sky130_fd_sc_hd__mux4_1
X_11356__1008 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__inv_2
X_09360_ net3190 _04612_ net609 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
X_06572_ top0.CPU.register.registers\[784\] top0.CPU.register.registers\[816\] top0.CPU.register.registers\[848\]
+ top0.CPU.register.registers\[880\] net929 net895 vssd1 vssd1 vccd1 vccd1 _03229_
+ sky130_fd_sc_hd__mux4_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08103__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09291_ _02362_ _04946_ _04947_ _04944_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.loadCt_n\[2\]
+ sky130_fd_sc_hd__o211a_1
X_08311_ net2813 net220 net415 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ net512 net150 net675 net420 net2538 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a32o_1
X_08173_ net512 net197 net623 net427 net2550 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_115_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08406__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10940__592 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__inv_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08957__A3 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ net337 _03780_ _03773_ net244 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a211o_1
X_07055_ _02375_ _03710_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__or2_2
XANTENNA__05756__A top0.CPU.control.funct7\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06006_ top0.CPU.register.registers\[263\] top0.CPU.register.registers\[295\] top0.CPU.register.registers\[327\]
+ top0.CPU.register.registers\[359\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02663_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12650__Q top0.MMIO.WBData_i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout493_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06276__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _04016_ net232 net227 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__and3_1
XANTENNA__07971__A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06050__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _03411_ net529 _03429_ _03443_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_52_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06579__S1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _04421_ net234 net229 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__and3_1
XANTENNA__08342__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ _05150_ _02729_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__nand2b_1
X_06839_ net871 _03495_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ net945 _02409_ _04217_ _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__o31ai_1
XFILLER_71_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08509_ net184 net685 net402 net368 net2527 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a32o_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ _02357_ net137 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__nor2_1
X_11520_ net1212 _01159_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08645__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06526__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275__927 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__inv_2
XANTENNA__07853__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ clknet_leaf_67_clk _01099_ net1120 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10204__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ clknet_leaf_79_clk _01030_ net1111 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08026__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316__968 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__inv_2
X_10333_ net2233 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09070__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ net3111 net119 net112 _05654_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XANTENNA__06261__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169__821 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__inv_2
X_10195_ net2803 net121 _05644_ _04903_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
X_12003_ net1695 _01642_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[496\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12560__Q top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout380 _04724_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_4
XANTENNA__06768__Y _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__A1 _02446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10883__535 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__inv_2
XANTENNA__08097__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ net767 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06944__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08636__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ net1410 _01357_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[211\]
+ sky130_fd_sc_hd__dfrtp_1
X_10924__576 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__inv_2
X_12698_ clknet_leaf_75_clk _02333_ net1124 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.storeCt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07844__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
X_11649_ net1341 _01288_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[142\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06008__Y _02665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07072__A1 _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold817 top0.CPU.register.registers\[155\] vssd1 vssd1 vccd1 vccd1 net3039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 top0.CPU.register.registers\[794\] vssd1 vssd1 vccd1 vccd1 net3050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold806 top0.CPU.register.registers\[535\] vssd1 vssd1 vccd1 vccd1 net3028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold839 top0.CPU.register.registers\[509\] vssd1 vssd1 vccd1 vccd1 net3061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06171__S net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08860_ net165 net3008 net353 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__mux2_1
XANTENNA__06258__S0 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08572__A1 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07811_ _04459_ _04460_ _04462_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__and4_1
X_10818__470 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__inv_2
X_08791_ net168 net686 net324 net292 net2512 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a32o_1
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07742_ _04396_ _04397_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and3_1
XANTENNA__07127__A2 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ _04327_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or2_1
XANTENNA__08875__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ net3438 _04949_ _05014_ _05019_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__a22o_1
X_06624_ _03265_ net532 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__nand2_1
XANTENNA__06430__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ top0.CPU.internalMem.state\[3\] top0.CPU.addrControl _04863_ _04987_ _04991_
+ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__a221o_1
XFILLER_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06555_ net749 _03211_ net858 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o21ai_2
X_09274_ _04851_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06486_ top0.CPU.register.registers\[277\] top0.CPU.register.registers\[309\] top0.CPU.register.registers\[341\]
+ top0.CPU.register.registers\[373\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03143_
+ sky130_fd_sc_hd__mux4_1
X_08225_ net510 net194 net686 net423 net2457 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a32o_1
X_11003__655 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__inv_2
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08561__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ net2935 net425 _04678_ net492 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a22o_1
XANTENNA__09052__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _03761_ _03762_ net465 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ net222 net692 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__and2_1
X_07038_ top0.CPU.register.registers\[159\] top0.CPU.register.registers\[191\] top0.CPU.register.registers\[223\]
+ top0.CPU.register.registers\[255\] net851 net816 vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__B1 _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08989_ top0.CPU.register.registers\[171\] net570 net557 vssd1 vssd1 vccd1 vccd1
+ _04794_ sky130_fd_sc_hd__o21a_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10570__222 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10867__519 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__inv_2
XANTENNA__06110__A _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ clknet_leaf_74_clk _02256_ net1127 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
X_10611__263 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__inv_2
XANTENNA__06972__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06109__X _02766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08094__A3 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ clknet_leaf_62_clk _02191_ net1094 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_11503_ clknet_leaf_83_clk _01142_ net1110 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12483_ net2175 _02122_ net1013 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[976\]
+ sky130_fd_sc_hd__dfrtp_1
X_11434_ clknet_leaf_68_clk _01082_ net1101 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09043__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_100_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10316_ _04993_ _05675_ _05676_ _05674_ net3366 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a32o_1
X_11355__1007 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__inv_2
X_10247_ net20 net656 net595 top0.MMIO.WBData_i\[26\] vssd1 vssd1 vccd1 vccd1 _02293_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08003__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1120 net1131 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07357__A2 _03997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ net141 _05633_ net660 vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08306__A1 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06412__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08609__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__A2 _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06340_ net786 _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__nand2_1
XANTENNA__05828__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06271_ top0.CPU.control.funct7\[1\] net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02928_
+ sky130_fd_sc_hd__a21oi_2
XANTENNA__07293__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08490__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08010_ net717 net502 net154 net549 net2337 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a32o_1
XANTENNA__09034__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold603 top0.CPU.register.registers\[445\] vssd1 vssd1 vccd1 vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06690__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338__990 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__inv_2
XANTENNA__08242__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold614 net39 vssd1 vssd1 vccd1 vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 top0.CPU.register.registers\[956\] vssd1 vssd1 vccd1 vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 top0.CPU.register.registers\[187\] vssd1 vssd1 vccd1 vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06479__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ net238 _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__or2_1
Xhold647 net72 vssd1 vssd1 vccd1 vccd1 net2869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 top0.CPU.register.registers\[656\] vssd1 vssd1 vccd1 vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 top0.CPU.register.registers\[955\] vssd1 vssd1 vccd1 vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ net713 net160 _04771_ net282 net3298 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__a32o_1
X_09892_ _05364_ _05388_ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a21o_1
X_10554__206 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__inv_2
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08843_ _04544_ net3091 net355 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__mux2_1
X_05986_ _02639_ _02642_ net737 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
XFILLER_85_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05753__B top0.CPU.control.funct7\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ net682 _04739_ net290 net2724 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__a22o_1
XANTENNA__06651__S0 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07725_ net486 _04333_ _04381_ _04011_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout456_A _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06403__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_clk_X clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _02831_ _03241_ net340 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06607_ net476 net471 net463 net449 net542 vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a41o_1
X_07587_ net482 _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and2_1
X_09326_ _04879_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nor2_1
X_06538_ net543 _02833_ _02496_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o21ai_1
X_10448__100 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__inv_2
XFILLER_138_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ top0.CPU.intMemAddr\[5\] _04612_ net769 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__mux2_1
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09387__S top0.CPU.control.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06469_ top0.CPU.register.registers\[276\] top0.CPU.register.registers\[308\] top0.CPU.register.registers\[340\]
+ top0.CPU.register.registers\[372\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03126_
+ sky130_fd_sc_hd__mux4_1
X_08208_ net152 net679 vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__and2_1
XFILLER_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06804__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09188_ top0.CPU.internalMem.state\[3\] top0.CPU.internalMem.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _04853_ sky130_fd_sc_hd__nand2b_1
X_10434__86 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__inv_2
XANTENNA__08291__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout992_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ net2620 _04630_ net429 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
X_11090__742 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__inv_2
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ net3291 net665 _05170_ _05571_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06890__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11131__783 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__inv_2
XFILLER_103_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10032_ top0.CPU.internalMem.pcOut\[30\] _05519_ net646 vssd1 vssd1 vccd1 vccd1 _02207_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05755__D1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11454__Q top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08974__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ net1675 _01622_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[476\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_80_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06494__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ clknet_leaf_92_clk _02239_ net1084 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12535_ clknet_leaf_76_clk _02174_ net1123 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07275__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08472__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995__647 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__inv_2
X_12466_ net2158 _02105_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[959\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06714__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09016__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11417_ clknet_leaf_69_clk _01065_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12397_ net2089 _02036_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[890\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08214__B net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05854__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06538__B1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_05840_ _02477_ _02496_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nand2_1
XFILLER_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06633__S0 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07750__A2 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889__541 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__inv_2
XANTENNA__05860__Y _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05771_ _02423_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__nor2_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _04083_ _04096_ _04124_ _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or4_1
XANTENNA__08884__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ _04691_ net397 net366 net2728 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a22o_1
X_07441_ _02684_ _03403_ net339 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a21o_1
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06936__S1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07372_ net490 _03746_ _04025_ _04012_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a31o_1
X_06323_ top0.CPU.control.funct7\[3\] net644 vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__nand2_1
X_09111_ _04700_ net279 net253 net2899 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a22o_1
XANTENNA__08058__A3 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08463__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ top0.CPU.register.registers\[131\] net565 vssd1 vssd1 vccd1 vccd1 _04807_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_13_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06254_ top0.CPU.register.registers\[921\] top0.CPU.register.registers\[953\] top0.CPU.register.registers\[985\]
+ top0.CPU.register.registers\[1017\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02911_
+ sky130_fd_sc_hd__mux4_1
XFILLER_135_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold400 top0.CPU.intMemAddr\[17\] vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 top0.CPU.register.registers\[295\] vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
X_11074__726 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__inv_2
X_06185_ top0.CPU.register.registers\[149\] top0.CPU.register.registers\[181\] top0.CPU.register.registers\[213\]
+ top0.CPU.register.registers\[245\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02842_
+ sky130_fd_sc_hd__mux4_1
Xhold422 top0.CPU.register.registers\[554\] vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold444 top0.CPU.register.registers\[382\] vssd1 vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 top0.CPU.register.registers\[601\] vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 top0.CPU.register.registers\[677\] vssd1 vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__A3 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold477 top0.CPU.register.registers\[530\] vssd1 vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 top0.CPU.register.registers\[309\] vssd1 vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06872__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold488 top0.CPU.register.registers\[41\] vssd1 vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ _02907_ _04519_ net585 vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__mux2_1
Xhold499 top0.CPU.intMemAddr\[25\] vssd1 vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
X_11115__767 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__inv_2
Xfanout924 net925 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_4
Xfanout913 net919 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_4
Xhold1100 top0.MMIO.WBData_i\[4\] vssd1 vssd1 vccd1 vccd1 net3322 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_4
X_09875_ net631 _02475_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__nand2_1
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
Xfanout968 net1004 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_2
Xhold1111 top0.CPU.register.registers\[233\] vssd1 vssd1 vccd1 vccd1 net3333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net982 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
Xhold1133 top0.display.dataforOutput\[5\] vssd1 vssd1 vccd1 vccd1 net3355 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net213 net669 net309 net285 net2281 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__a32o_1
Xhold1122 top0.CPU.register.registers\[152\] vssd1 vssd1 vccd1 vccd1 net3344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _02173_ vssd1 vssd1 vccd1 vccd1 net3388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 top0.MISOtoMMIO\[7\] vssd1 vssd1 vccd1 vccd1 net3377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 top0.CPU.internalMem.storeCt\[1\] vssd1 vssd1 vccd1 vccd1 net3366 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07741__A2 _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1177 top0.CPU.intMem_out\[11\] vssd1 vssd1 vccd1 vccd1 net3399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 top0.CPU.intMem_out\[28\] vssd1 vssd1 vccd1 vccd1 net3421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1188 top0.display.delayctr\[19\] vssd1 vssd1 vccd1 vccd1 net3410 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net172 net616 net312 net293 net3019 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__a32o_1
X_05969_ net725 _02625_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ net168 net696 net322 net299 net2964 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a32o_1
X_07708_ _03913_ _03940_ _04344_ _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_49_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11009__661 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__inv_2
XANTENNA__07043__X _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354__1006 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__inv_2
X_07639_ _03385_ _03407_ _03409_ _03560_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__or4_1
XFILLER_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10682__334 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__inv_2
XANTENNA__08049__A3 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _04951_ _04953_ _04961_ vssd1 vssd1 vccd1 vccd1 top0.display.next_state\[1\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ net2012 _01959_ net1044 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06534__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net1943 _01890_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[744\]
+ sky130_fd_sc_hd__dfrtp_1
X_10723__375 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__inv_2
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__B1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08034__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__Q top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__A3 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net1874 _01821_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[675\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__B net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10015_ top0.CPU.internalMem.pcOut\[29\] _05492_ vssd1 vssd1 vccd1 vccd1 _05504_
+ sky130_fd_sc_hd__and2_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05680__Y _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ net1658 _01605_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[459\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07040__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08693__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ net1589 _01536_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12518_ net2210 _02157_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1011\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12449_ net2141 _02088_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[942\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06854__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07990_ _04260_ net231 net226 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__and3_2
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout209 _04510_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
X_06941_ _03596_ _03597_ net756 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__mux2_1
X_09660_ _04955_ _04959_ _05176_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__or3b_1
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ net721 net198 net325 net331 net2405 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a32o_1
X_06872_ top0.CPU.register.registers\[521\] top0.CPU.register.registers\[553\] top0.CPU.register.registers\[585\]
+ top0.CPU.register.registers\[617\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03529_
+ sky130_fd_sc_hd__mux4_1
XFILLER_95_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06082__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07870__A1_N _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05823_ _02478_ _02479_ net729 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
X_09591_ _04957_ _05131_ net661 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__o21a_1
X_08542_ net188 net672 net398 net363 net2536 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__a32o_1
X_05754_ top0.CPU.control.funct7\[1\] top0.CPU.control.funct7\[0\] _02410_ vssd1 vssd1
+ vccd1 vccd1 _02411_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_38_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07031__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ net194 net622 net403 net372 net2720 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a32o_1
XANTENNA__08279__A3 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05685_ net944 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__inv_2
X_07424_ _02666_ _03261_ _03738_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__and3_1
X_10666__318 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__inv_2
XANTENNA_fanout154_A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08834__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout321_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ _03747_ _03835_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1063_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707__359 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__inv_2
XANTENNA_fanout419_A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07286_ _03176_ _03196_ _03942_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__or3_1
X_06306_ top0.CPU.register.registers\[668\] top0.CPU.register.registers\[700\] top0.CPU.register.registers\[732\]
+ top0.CPU.register.registers\[764\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02963_
+ sky130_fd_sc_hd__mux4_1
X_06237_ top0.CPU.register.registers\[792\] top0.CPU.register.registers\[824\] top0.CPU.register.registers\[856\]
+ top0.CPU.register.registers\[888\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02894_
+ sky130_fd_sc_hd__mux4_1
X_09025_ net222 net3198 net349 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__mux2_1
XANTENNA__08739__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404__56 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__inv_2
XANTENNA_fanout207_X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 top0.CPU.register.registers\[204\] vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07947__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06168_ top0.CPU.register.registers\[400\] top0.CPU.register.registers\[432\] top0.CPU.register.registers\[464\]
+ top0.CPU.register.registers\[496\] net846 net811 vssd1 vssd1 vccd1 vccd1 _02825_
+ sky130_fd_sc_hd__mux4_1
Xhold241 top0.CPU.register.registers\[999\] vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 top0.CPU.register.registers\[67\] vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 top0.CPU.register.registers\[716\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08141__Y _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06099_ _02754_ _02755_ net786 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
Xhold296 top0.CPU.register.registers\[201\] vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06845__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 top0.CPU.register.registers\[619\] vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05765__Y _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold285 top0.CPU.register.registers\[110\] vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_4
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_113_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09927_ top0.CPU.internalMem.pcOut\[23\] _05421_ vssd1 vssd1 vccd1 vccd1 _05422_
+ sky130_fd_sc_hd__xor2_1
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_2
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_8
Xfanout743 net744 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_6
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout776 net779 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_4
Xfanout787 top0.CPU.control.rs2\[2\] vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_8
X_09858_ top0.CPU.internalMem.pcOut\[17\] _05348_ vssd1 vssd1 vccd1 vccd1 _05359_
+ sky130_fd_sc_hd__and2_1
XFILLER_73_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_2
X_09789_ _05273_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ _04716_ net321 net287 net2747 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a22o_1
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11820_ net1512 _01459_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05941__B _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ net1443 _01390_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
X_11243__895 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__inv_2
XFILLER_14_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08675__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11682_ net1374 _01321_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[175\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12303_ net1995 _01942_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[796\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07650__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12234_ net1926 _01873_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[727\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ net1857 _01804_ net1038 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[658\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07402__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12096_ net1788 _01735_ net1044 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[589\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_10_0_clk_X clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06064__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09604__A _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09323__B top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07469__A1 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_71_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08666__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ net1641 _01588_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08681__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08418__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10225__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ net474 _03054_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nor2_1
XFILLER_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09091__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07071_ _03723_ _03727_ net348 vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__mux2_1
X_06022_ top0.CPU.register.registers\[134\] top0.CPU.register.registers\[166\] top0.CPU.register.registers\[198\]
+ top0.CPU.register.registers\[230\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02679_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08197__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353__1005 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__inv_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ top0.CPU.internalMem.pcOut\[5\] _05211_ _05199_ vssd1 vssd1 vccd1 vccd1 _05224_
+ sky130_fd_sc_hd__o21a_1
X_07973_ top0.CPU.intMem_out\[7\] net629 _04588_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06203__A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06924_ _03094_ _03115_ _03579_ _03580_ _03093_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__o32a_1
X_11186__838 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__inv_2
XANTENNA__05959__B1_N _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06855_ _03508_ _03509_ _03510_ _03511_ net761 net751 vssd1 vssd1 vccd1 vccd1 _03512_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06055__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _02505_ _02511_ _05150_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__o21bai_4
XANTENNA_fanout271_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05806_ net786 _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__and2_1
X_09574_ top0.CPU.internalMem.pcOut\[1\] _05120_ _05110_ vssd1 vssd1 vccd1 vccd1 _01124_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout369_A _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227__879 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__inv_2
XFILLER_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08525_ _04710_ net388 net361 net3185 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a22o_1
X_06786_ net859 _03434_ _03438_ _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
X_05737_ top0.CPU.decoder.instruction\[11\] _02393_ vssd1 vssd1 vccd1 vccd1 _02394_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08657__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ _04673_ net405 net371 net2669 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
XANTENNA__08564__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ net948 net545 net700 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__or3b_1
XANTENNA__08409__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07407_ net529 net528 _03482_ net527 net468 net460 vssd1 vssd1 vccd1 vccd1 _04064_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07338_ _03221_ net533 net529 net528 net467 net459 vssd1 vssd1 vccd1 vccd1 _03995_
+ sky130_fd_sc_hd__mux4_1
XFILLER_129_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09082__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ net486 net481 vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__nand2_4
XFILLER_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10280_ net3247 net119 net112 _05168_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a22o_1
X_09008_ net224 net3107 net350 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_105_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06818__S0 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10794__446 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__inv_2
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout551 _04958_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06113__A _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _02434_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
XANTENNA__06294__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835__487 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__inv_2
Xfanout573 net574 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_4
Xfanout562 _04477_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_2
Xfanout584 _02421_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
XANTENNA__08896__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06046__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10688__340 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__inv_2
XANTENNA__11462__Q top0.CPU.decoder.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11803_ net1495 _01442_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[296\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_53_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08648__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11734_ net1426 _01373_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07320__A0 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ net1357 _01304_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[158\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07871__A1 top0.CPU.intMem_out\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10729__381 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__inv_2
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10207__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09073__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ net1288 _01235_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08820__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12217_ net1909 _01856_ net980 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10395__47 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__inv_2
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12148_ net1840 _01787_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07119__A _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12079_ net1771 _01718_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[572\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06037__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08887__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ top0.CPU.register.registers\[131\] top0.CPU.register.registers\[163\] top0.CPU.register.registers\[195\]
+ top0.CPU.register.registers\[227\] net916 net882 vssd1 vssd1 vccd1 vccd1 _03297_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09053__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_06571_ _03226_ _03227_ net762 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__mux2_1
XANTENNA__08639__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09290_ _02362_ _04946_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__nand2_1
X_08310_ net3163 net181 net416 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__mux2_1
XANTENNA__08103__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ net946 _02399_ net677 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__nand3_4
XANTENNA_14 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08406__A3 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ net507 net199 net619 net427 net2375 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a32o_1
XANTENNA__09603__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__X _03637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09064__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08811__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481__133 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__inv_2
XANTENNA__07614__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__B2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07123_ _03778_ _03779_ net465 vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__mux2_1
X_07054_ net944 _02408_ _02411_ _03709_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout117_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_06005_ top0.CPU.register.registers\[391\] top0.CPU.register.registers\[423\] top0.CPU.register.registers\[455\]
+ top0.CPU.register.registers\[487\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02662_
+ sky130_fd_sc_hd__mux4_1
X_10522__174 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__inv_2
XANTENNA__05756__B top0.CPU.control.funct7\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06276__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07956_ net718 net504 net188 net547 net2333 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a32o_1
XANTENNA__08559__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ _03426_ _03445_ _03484_ _03563_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_52_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ net2782 net549 net500 _04534_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XANTENNA__08878__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06838_ top0.CPU.register.registers\[907\] top0.CPU.register.registers\[939\] top0.CPU.register.registers\[971\]
+ top0.CPU.register.registers\[1003\] net929 net895 vssd1 vssd1 vccd1 vccd1 _03495_
+ sky130_fd_sc_hd__mux4_1
X_09626_ net3330 net605 net658 net3255 _05157_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__a221o_1
XANTENNA__05787__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout820_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ _05102_ _05103_ _05104_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__and3_1
X_06769_ _03411_ net529 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_35_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
X_09488_ top0.MMIO.WBData_i\[20\] net149 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__and2_1
X_08508_ net186 net683 net398 net367 net2292 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ net3099 net221 net374 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11947__RESET_B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ clknet_leaf_67_clk _01098_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09055__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ clknet_leaf_79_clk _01029_ net1111 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08802__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ net2229 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09358__A1 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ net1694 _01641_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[495\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10263_ _04932_ net577 _05144_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__or3b_1
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ _05639_ _05642_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__nor2_1
XANTENNA__06041__B1 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05682__A top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_8
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06019__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout370 _04727_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06130__X _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10140__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05778__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_45_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11352__1004 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__inv_2
X_12766_ net58 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11717_ net1409 _01356_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[210\]
+ sky130_fd_sc_hd__dfrtp_1
X_12697_ clknet_leaf_93_clk _02332_ net1082 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_10465__117 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__inv_2
X_11648_ net1340 _01287_ net1035 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[141\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05950__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
X_11579_ net1271 _01218_ net1009 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506__158 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__inv_2
Xhold818 top0.CPU.register.registers\[411\] vssd1 vssd1 vccd1 vccd1 net3040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold807 top0.CPU.register.registers\[750\] vssd1 vssd1 vccd1 vccd1 net3029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09349__A1 _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold829 top0.CPU.register.registers\[390\] vssd1 vssd1 vccd1 vccd1 net3051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08520__X _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08021__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06258__S1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ net172 net681 net312 net289 net2513 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a32o_1
X_07810_ _04463_ _04464_ _04465_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__and4_1
XANTENNA__06583__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _02925_ _03600_ net446 _04391_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__o31a_1
XANTENNA__06040__X _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07532__B1 _03540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06335__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ net244 _03825_ _04328_ net452 vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09411_ _02355_ net147 net143 _02363_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__o22ai_1
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06623_ _03265_ net532 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nor2_1
XANTENNA__06430__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _02365_ _04864_ _04944_ _04990_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06554_ _03209_ _03210_ net869 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08088__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ _04852_ _04864_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__and2_1
XANTENNA__07835__A1 top0.CPU.intMem_out\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06485_ net866 _03141_ _03138_ net859 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__o211a_1
XANTENNA__05750__D_N top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042__694 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__inv_2
X_08224_ net3119 net422 _04703_ net502 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a22o_1
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08842__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08155_ net208 net614 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and2_1
X_07106_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__inv_2
X_08086_ net508 net203 net695 net434 net2262 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a32o_1
XFILLER_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07037_ net779 _03689_ net773 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_54_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08797__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08988_ _04587_ net699 _04793_ net262 net3281 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__a32o_1
XANTENNA__08289__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ _04452_ net234 net229 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06110__B _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06326__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07523__B1 _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09609_ net141 _05144_ net660 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ clknet_leaf_98_clk _02255_ net1076 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10947__599 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__inv_2
XANTENNA__07826__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ clknet_leaf_61_clk _02190_ net1094 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06185__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12482_ net2174 _02121_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[975\]
+ sky130_fd_sc_hd__dfrtp_1
X_11502_ clknet_leaf_81_clk net3095 net1109 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ clknet_leaf_70_clk _01081_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05932__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__A2 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10315_ top0.CPU.internalMem.storeCt\[0\] top0.CPU.internalMem.storeCt\[1\] vssd1
+ vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__nand2_1
XFILLER_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10246_ net19 net653 net592 net3392 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__o22a_1
X_10365__17 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__inv_2
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1121 net1131 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_4
Xfanout1132 top0.CPU.internalMem.nrst vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_8
XFILLER_105_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1110 net1115 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_4
X_10850__502 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__inv_2
X_10177_ net550 _03020_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nand2b_1
XANTENNA__05999__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06565__A1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__10113__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06412__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026__678 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__inv_2
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06270_ _02457_ net242 _02908_ _02925_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__and4_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05923__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07278__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold626 top0.CPU.register.registers\[915\] vssd1 vssd1 vccd1 vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 top0.CPU.register.registers\[446\] vssd1 vssd1 vccd1 vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06479__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 top0.CPU.register.registers\[899\] vssd1 vssd1 vccd1 vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09960_ _05451_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__xor2_1
Xhold659 top0.CPU.register.registers\[508\] vssd1 vssd1 vccd1 vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
Xhold637 top0.CPU.register.registers\[215\] vssd1 vssd1 vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 top0.CPU.register.registers\[696\] vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08911_ top0.CPU.register.registers\[226\] net565 net553 vssd1 vssd1 vccd1 vccd1
+ _04771_ sky130_fd_sc_hd__o21a_1
X_09891_ top0.CPU.internalMem.pcOut\[18\] _05362_ _05376_ _05375_ vssd1 vssd1 vccd1
+ vccd1 _05389_ sky130_fd_sc_hd__a31o_1
XANTENNA__08545__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10593__245 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__inv_2
X_08842_ net204 net3012 net354 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__mux2_1
X_05985_ _02640_ _02641_ net728 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
XANTENNA__05753__C top0.CPU.control.funct7\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ _04697_ net307 net289 net2764 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__a22o_1
XANTENNA__06651__S1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_A _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06172__A1_N net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ _03719_ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08837__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07655_ net443 _04150_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__nand2_1
X_10634__286 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__inv_2
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1093_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _03250_ _03261_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout449_A _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06403__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _04059_ _04064_ net478 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
XANTENNA__12656__Q top0.MMIO.WBData_i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ _04524_ _04868_ _04869_ _04872_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__or4_1
X_06537_ net543 _02496_ _02833_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__or3_1
XANTENNA__07977__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _04901_ _04905_ _04909_ _04917_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ top0.CPU.register.registers\[404\] top0.CPU.register.registers\[436\] top0.CPU.register.registers\[468\]
+ top0.CPU.register.registers\[500\] net918 net884 vssd1 vssd1 vccd1 vccd1 _03125_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout616_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08207_ net3056 net422 _04696_ net500 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
X_09187_ top0.CPU.internalMem.state\[3\] top0.CPU.internalMem.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _04852_ sky130_fd_sc_hd__and2b_1
X_10528__180 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__inv_2
X_06399_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__inv_2
X_08138_ net2954 net161 net429 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout985_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ net2891 net433 _04657_ net494 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a22o_1
X_10100_ _05569_ _05570_ net601 vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351__1003 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__inv_2
XANTENNA__09733__A1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net235 _05515_ _05516_ _05517_ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a32o_1
XANTENNA__06890__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06547__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11982_ net1674 _01621_ net992 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[475\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__11470__Q top0.CPU.control.funct7\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ clknet_leaf_92_clk _02238_ net1080 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12534_ clknet_leaf_77_clk net3388 net1123 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06158__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05905__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ net2157 _02104_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[958\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07680__C1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11416_ clknet_leaf_77_clk _01064_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08224__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12396_ net2088 _02035_ net984 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10031__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10577__229 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10229_ net32 net656 net595 top0.MMIO.WBData_i\[8\] vssd1 vssd1 vccd1 vccd1 _02275_
+ sky130_fd_sc_hd__a22o_1
Xhold1 top0.CPU.register.registers\[30\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05770_ _02411_ _02415_ _02426_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__o21bai_2
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07561__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ net443 _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__nand2_1
XFILLER_50_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11632__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09061__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07371_ _03850_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__or2_1
X_06322_ net771 _02978_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__or2_1
XANTENNA__06149__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ _04699_ net555 _04828_ net252 net3103 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_33_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09041_ net214 net3214 net349 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__mux2_1
X_06253_ top0.CPU.control.funct7\[0\] net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02910_
+ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_13_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08215__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 top0.CPU.register.registers\[834\] vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
X_06184_ _02837_ _02840_ net780 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
Xhold423 top0.CPU.register.registers\[714\] vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold412 top0.CPU.intMemAddr\[11\] vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__A1 top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold434 top0.CPU.register.registers\[848\] vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__C1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 top0.CPU.register.registers\[576\] vssd1 vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07974__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 top0.CPU.register.registers\[454\] vssd1 vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 top0.CPU.register.registers\[380\] vssd1 vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 top0.CPU.register.registers\[433\] vssd1 vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 top0.CPU.register.registers\[575\] vssd1 vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06872__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08421__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09943_ _05345_ _05391_ _05431_ _05433_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a311o_1
Xfanout914 net916 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_4
Xfanout947 net949 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_2
X_09874_ net587 _02475_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout958 net962 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
XANTENNA__08518__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1106_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ net167 net674 net324 net288 net2376 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a32o_1
Xhold1101 top0.CPU.register.registers\[990\] vssd1 vssd1 vccd1 vccd1 net3323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 top0.display.dataforOutput\[11\] vssd1 vssd1 vccd1 vccd1 net3334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 top0.CPU.register.registers\[388\] vssd1 vssd1 vccd1 vccd1 net3345 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 net976 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
Xhold1156 _02177_ vssd1 vssd1 vccd1 vccd1 net3378 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 top0.CPU.register.registers\[562\] vssd1 vssd1 vccd1 vccd1 net3367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1167 top0.display.counter\[0\] vssd1 vssd1 vccd1 vccd1 net3389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1134 _01135_ vssd1 vssd1 vccd1 vccd1 net3356 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A3 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1178 top0.display.delayctr\[9\] vssd1 vssd1 vccd1 vccd1 net3400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08756_ net176 net615 net318 net295 net2498 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__a32o_1
Xhold1189 top0.display.delayctr\[2\] vssd1 vssd1 vccd1 vccd1 net3411 sky130_fd_sc_hd__dlygate4sd3_1
X_05968_ top0.CPU.register.registers\[900\] top0.CPU.register.registers\[932\] top0.CPU.register.registers\[964\]
+ top0.CPU.register.registers\[996\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02625_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08567__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05899_ top0.CPU.decoder.instruction\[9\] _02448_ vssd1 vssd1 vccd1 vccd1 _02556_
+ sky130_fd_sc_hd__nand2_1
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07707_ _04354_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__or2_1
X_08687_ net172 net692 net312 net298 net2282 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06388__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout733_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ _04069_ _04088_ _04232_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__or4bb_1
XFILLER_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout900_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07569_ net462 _03812_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ net660 _04959_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ top0.CPU.internalMem.pcOut\[0\] top0.CPU.addrControl _04899_ _04900_ vssd1
+ vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a22o_1
X_12250_ net1942 _01889_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[743\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06560__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ net1873 _01820_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06768__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05955__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold990 top0.CPU.register.registers\[986\] vssd1 vssd1 vccd1 vccd1 net3212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06550__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08509__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_73_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248__900 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__inv_2
XANTENNA__09861__S net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _05499_ _05501_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09182__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05690__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ net1657 _01604_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[458\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06379__S0 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07040__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10962__614 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__inv_2
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11896_ net1588 _01535_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[389\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11097__749 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__inv_2
X_12517_ net2209 _02156_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1010\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08996__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12448_ net2140 _02087_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[941\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08748__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ net2071 _02018_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[872\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05865__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06854__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ top0.CPU.register.registers\[281\] top0.CPU.register.registers\[313\] top0.CPU.register.registers\[345\]
+ top0.CPU.register.registers\[377\] net910 net876 vssd1 vssd1 vccd1 vccd1 _03597_
+ sky130_fd_sc_hd__mux4_1
X_06871_ top0.CPU.register.registers\[649\] top0.CPU.register.registers\[681\] top0.CPU.register.registers\[713\]
+ top0.CPU.register.registers\[745\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03528_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09173__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08381__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ net719 net200 net319 net331 net2311 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a32o_1
X_05822_ top0.CPU.register.registers\[786\] top0.CPU.register.registers\[818\] top0.CPU.register.registers\[850\]
+ top0.CPU.register.registers\[882\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02479_
+ sky130_fd_sc_hd__mux4_1
XFILLER_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08920__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09590_ _02596_ _05007_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08541_ net192 net677 net407 net364 net2791 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a32o_1
X_05753_ top0.CPU.control.funct7\[3\] top0.CPU.control.funct7\[2\] top0.CPU.control.funct7\[4\]
+ top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__or4_1
X_05684_ net942 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__inv_2
XFILLER_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08472_ _04686_ net394 net370 net2693 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07423_ _03934_ _04078_ _04079_ net482 net454 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_18_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11350__1002 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__inv_2
XFILLER_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07354_ _03850_ _04009_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nor2_1
XANTENNA__08436__A1 _04561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10746__398 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__inv_2
XANTENNA__08987__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ _03243_ _03941_ _03198_ _03223_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a211oi_1
X_06305_ net580 _02946_ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a21o_1
XANTENNA__09011__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06447__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07644__C1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ _04555_ net2994 net351 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1056_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06236_ _02891_ _02892_ net731 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold220 top0.CPU.register.registers\[225\] vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 top0.CPU.register.registers\[493\] vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ _02822_ _02823_ net728 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
Xhold231 top0.CPU.register.registers\[198\] vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 top0.CPU.register.registers\[227\] vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
X_10599__251 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__inv_2
Xhold286 top0.CPU.register.registers\[492\] vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _04652_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
X_06098_ top0.CPU.register.registers\[908\] top0.CPU.register.registers\[940\] top0.CPU.register.registers\[972\]
+ top0.CPU.register.registers\[1004\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02755_
+ sky130_fd_sc_hd__mux4_1
Xhold264 top0.CPU.register.registers\[745\] vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05958__C1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06845__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 top0.CPU.register.registers\[742\] vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout722 net723 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_113_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09926_ net585 _04524_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__a21o_1
Xhold297 top0.CPU.register.registers\[740\] vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout733 net734 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_4
Xfanout766 _02344_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
Xfanout755 _02345_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_4
XANTENNA__09164__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout744 _02347_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_4
XANTENNA__07990__A _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout850_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _05353_ _05354_ _05356_ net239 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a31o_1
Xfanout777 net779 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_4
Xfanout799 top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_2
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08372__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 net790 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_4
X_09788_ top0.CPU.internalMem.pcOut\[12\] _05293_ vssd1 vssd1 vccd1 vccd1 _05294_
+ sky130_fd_sc_hd__xor2_2
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08297__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _04715_ net315 net286 net2677 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a22o_1
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08739_ net617 _04739_ net294 net2595 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a22o_1
X_11750_ net1442 _01389_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ net1373 _01320_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[174\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08427__A1 _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08978__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06533__S0 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12302_ net1994 _01941_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[795\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12233_ net1925 _01872_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[726\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07938__B1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ net1856 _01803_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07402__A2 _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12095_ net1787 _01734_ net1097 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[588\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_110_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09155__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05691__Y _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08902__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07013__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ net1640 _01587_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[441\]
+ sky130_fd_sc_hd__dfrtp_1
X_11879_ net1571 _01518_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08969__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06429__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06524__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ _03724_ _03726_ net455 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__mux2_1
XANTENNA__12083__RESET_B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06021_ _02676_ _02677_ net782 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
XANTENNA__12012__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09146__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _05201_ _05212_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__nand2_1
X_07972_ net562 _04604_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__or2_1
X_06923_ _03078_ net537 _03096_ net536 vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__o22a_1
X_06854_ top0.CPU.register.registers\[522\] top0.CPU.register.registers\[554\] top0.CPU.register.registers\[586\]
+ top0.CPU.register.registers\[618\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__mux4_1
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09642_ net3293 net604 net659 top0.display.dataforOutput\[14\] _05167_ vssd1 vssd1
+ vccd1 vccd1 _01144_ sky130_fd_sc_hd__a221o_1
XANTENNA__09006__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05805_ top0.CPU.register.registers\[915\] top0.CPU.register.registers\[947\] top0.CPU.register.registers\[979\]
+ top0.CPU.register.registers\[1011\] net856 net821 vssd1 vssd1 vccd1 vccd1 _02462_
+ sky130_fd_sc_hd__mux4_1
X_09573_ _05114_ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06785_ net753 _03441_ net746 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__o21ai_1
X_05736_ net954 net947 net950 net952 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__or4_2
XANTENNA__11482__D top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ _04709_ net392 net361 net2591 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout264_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08106__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08845__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ net151 net622 net404 net371 net2347 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout431_A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout529_A _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07406_ _03993_ _04062_ net461 vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__mux2_1
X_08386_ net153 net705 net394 net382 net2454 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a32o_1
XFILLER_137_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ _03482_ net526 net527 _03519_ net458 net468 vssd1 vssd1 vccd1 vccd1 _03994_
+ sky130_fd_sc_hd__mux4_1
XFILLER_137_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ net489 _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__nand2_1
X_09007_ net212 net3053 net351 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
XANTENNA__09909__A1 top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06840__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ _03005_ _03053_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__or2_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06219_ top0.CPU.register.registers\[918\] top0.CPU.register.registers\[950\] top0.CPU.register.registers\[982\]
+ top0.CPU.register.registers\[1014\] net838 net803 vssd1 vssd1 vccd1 vccd1 _02876_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06818__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_3_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08188__A3 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout541 _02434_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_2
Xfanout530 _03379_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_2
XANTENNA__09137__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ top0.CPU.internalMem.pcOut\[21\] _05394_ _05405_ vssd1 vssd1 vccd1 vccd1
+ _05406_ sky130_fd_sc_hd__a21o_1
XANTENNA__08345__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net576 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_2
Xfanout563 _04477_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_70_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11210__862 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__inv_2
Xfanout552 net554 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_4
Xfanout596 _05647_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_2
Xfanout585 net588 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_2
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11802_ net1494 _01441_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[295\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12594__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net1425 _01372_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07320__A1 _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11664_ net1356 _01303_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[157\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10207__A1 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11595_ net1287 _01234_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05686__Y _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ net1908 _01855_ net1029 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08179__A3 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06304__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ net1839 _01786_ net1059 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[640\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07119__B _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09128__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11405__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ net1770 _01717_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[571\]
+ sky130_fd_sc_hd__dfrtp_1
X_10968__620 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06347__C1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08351__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06993__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06570_ top0.CPU.register.registers\[528\] top0.CPU.register.registers\[560\] top0.CPU.register.registers\[592\]
+ top0.CPU.register.registers\[624\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03227_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08103__A3 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08240_ net951 net953 net955 vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or3b_1
X_08171_ net3140 net425 _04685_ net494 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XANTENNA__07075__A0 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ net520 net521 net473 vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
X_07053_ net944 _02408_ _02411_ _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a31oi_2
X_11153__805 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06004_ top0.CPU.register.registers\[7\] top0.CPU.register.registers\[39\] top0.CPU.register.registers\[71\]
+ top0.CPU.register.registers\[103\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02661_
+ sky130_fd_sc_hd__mux4_1
XFILLER_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05756__C top0.CPU.control.funct7\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ top0.CPU.internalMem.pcOut\[11\] net639 net636 _04591_ vssd1 vssd1 vccd1
+ vccd1 _04592_ sky130_fd_sc_hd__o211a_2
XANTENNA__06050__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05772__B _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ _03464_ _03485_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__nor2_1
XFILLER_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout479_A _02575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08342__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ net141 _05156_ net660 vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a21oi_1
X_07886_ net717 net205 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout646_A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ top0.CPU.register.registers\[779\] top0.CPU.register.registers\[811\] top0.CPU.register.registers\[843\]
+ top0.CPU.register.registers\[875\] net929 net895 vssd1 vssd1 vccd1 vccd1 _03494_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06984__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05787__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06768_ net747 _03424_ _03419_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08575__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09556_ _02406_ _05002_ _04175_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ net192 net688 net407 net368 net2856 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a32o_1
X_09487_ _02352_ net148 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05719_ top0.CPU.Op\[5\] _02371_ _02373_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__or3_4
X_06699_ net746 _03355_ _03347_ _03348_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__o2bb2a_2
X_08438_ net2983 net198 net375 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
XFILLER_62_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06416__A1_N net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761__413 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__inv_2
XANTENNA__07853__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ _04650_ net389 net381 net3239 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a22o_1
XANTENNA__06823__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ clknet_leaf_85_clk _01028_ net1111 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10331_ net2245 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10802__454 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__inv_2
X_10262_ net3084 net119 net112 _05142_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
XANTENNA__11916__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ net1693 _01640_ net1059 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[494\]
+ sky130_fd_sc_hd__dfrtp_1
X_10193_ _04907_ net129 net121 net3231 net115 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a221o_1
XANTENNA__06041__A1 top0.CPU.control.funct7\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout360 _04744_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_4
Xfanout393 net408 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_2
Xfanout382 net384 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11473__Q top0.CPU.control.funct7\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05778__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__C1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11716_ net1408 _01355_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[209\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ clknet_leaf_80_clk _02331_ net1113 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
X_11647_ net1339 _01286_ net1101 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[140\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 gpio_in[2] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06733__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11578_ net1270 _01217_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05950__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold819 top0.CPU.register.registers\[414\] vssd1 vssd1 vccd1 vccd1 net3041 sky130_fd_sc_hd__dlygate4sd3_1
X_10545__197 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__inv_2
Xhold808 top0.CPU.register.registers\[218\] vssd1 vssd1 vccd1 vccd1 net3030 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11657__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09048__C _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08021__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06321__X _02978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ net442 _04135_ _04394_ _04395_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ net477 _03758_ _03788_ _04323_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_125_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09410_ net3434 _04949_ _05018_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__a21o_1
X_06622_ net747 _03278_ _03273_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a21oi_4
X_09341_ top0.CPU.internalMem.loadCt\[0\] top0.CPU.internalMem.loadCt\[2\] top0.CPU.internalMem.loadCt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or3b_1
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08088__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06553_ top0.CPU.register.registers\[913\] top0.CPU.register.registers\[945\] top0.CPU.register.registers\[977\]
+ top0.CPU.register.registers\[1009\] net913 net879 vssd1 vssd1 vccd1 vccd1 _03210_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _02364_ _04863_ _04929_ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__nand4_2
X_06484_ _03139_ _03140_ net764 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__mux2_1
X_08223_ net221 net682 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06643__S net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ net3191 net425 _04677_ net491 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a22o_1
X_08085_ net2909 net436 _04665_ net515 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a22o_1
XANTENNA__08796__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ net536 net537 net473 vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__mux2_1
X_07036_ net738 _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__nor2_1
XANTENNA__11398__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06271__A1 top0.CPU.control.funct7\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05783__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ top0.CPU.register.registers\[172\] net575 _04754_ vssd1 vssd1 vccd1 vccd1
+ _04793_ sky130_fd_sc_hd__o21a_1
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout763_A _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ net3181 net549 net502 _04577_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a22o_1
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout930_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11281__933 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__inv_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06110__C _02766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ net550 _05006_ _02649_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06957__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ net873 _05069_ net125 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XANTENNA__07062__X _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322__974 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06709__S0 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08079__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ clknet_leaf_61_clk _02189_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06185__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11501_ clknet_leaf_82_clk _01140_ net1109 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12481_ net2173 _02120_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[974\]
+ sky130_fd_sc_hd__dfrtp_1
X_11432_ clknet_leaf_70_clk _01080_ net1120 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05932__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11468__Q top0.CPU.control.funct7\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10314_ _05675_ _05674_ net3436 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08539__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net18 net657 net596 top0.MMIO.WBData_i\[24\] vssd1 vssd1 vccd1 vccd1 _02291_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08003__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout1122 net1131 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_2
Xfanout1100 net1105 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_2
Xfanout1111 net1114 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_4
X_10176_ net3440 net664 _05141_ _05629_ _05632_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a221o_1
XFILLER_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05999__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _04587_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
XFILLER_94_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930__582 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__inv_2
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload5_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06029__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ clknet_leaf_81_clk _02314_ net1112 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05828__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05923__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08778__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold627 top0.CPU.register.registers\[580\] vssd1 vssd1 vccd1 vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 top0.CPU.register.registers\[516\] vssd1 vssd1 vccd1 vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09059__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold605 top0.CPU.register.registers\[693\] vssd1 vssd1 vccd1 vccd1 net2827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 top0.CPU.intMem_out\[0\] vssd1 vssd1 vccd1 vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06253__A1 top0.CPU.control.funct7\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold649 top0.CPU.register.registers\[666\] vssd1 vssd1 vccd1 vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ _05377_ _05354_ _05363_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__and3b_1
X_08910_ net715 net164 net270 net282 net2475 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__a32o_1
XANTENNA__08545__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ net205 net3202 net354 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__mux2_1
XANTENNA__07202__A0 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11265__917 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__inv_2
XFILLER_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08950__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05984_ top0.CPU.register.registers\[517\] top0.CPU.register.registers\[549\] top0.CPU.register.registers\[581\]
+ top0.CPU.register.registers\[613\] net849 net814 vssd1 vssd1 vccd1 vccd1 _02641_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05753__D top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ _04696_ net314 net290 net2679 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__a22o_1
X_07723_ net338 _03792_ _03803_ _02577_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ net487 net245 vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__or2_1
XANTENNA__06939__S0 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306__958 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__inv_2
X_06605_ _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__inv_2
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout1086_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07585_ _03907_ _03933_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__or2_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ top0.CPU.internalMem.state\[1\] top0.CPU.internalMem.state\[0\] _02365_ vssd1
+ vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__and3_1
XANTENNA__08853__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06536_ net747 _03192_ _03184_ _03185_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout511_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159__811 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__inv_2
X_09255_ _04903_ _04907_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__or3_1
X_06467_ top0.CPU.register.registers\[20\] top0.CPU.register.registers\[52\] top0.CPU.register.registers\[84\]
+ top0.CPU.register.registers\[116\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03124_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06373__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ net207 net682 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__and2_1
X_09186_ top0.CPU.internalMem.state\[1\] top0.CPU.internalMem.state\[2\] top0.CPU.internalMem.state\[3\]
+ top0.CPU.internalMem.state\[0\] vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__and4bb_1
X_06398_ _03041_ _03053_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__or2_1
XANTENNA__08769__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ net2826 net165 net429 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
XANTENNA__08784__A3 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout880_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ net210 net692 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__and2_1
X_07019_ net763 _03673_ net751 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__a21o_1
XANTENNA__07992__A1 top0.CPU.intMem_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873__525 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__inv_2
XANTENNA_fanout978_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ top0.CPU.internalMem.pcOut\[30\] _05504_ net238 vssd1 vssd1 vccd1 vccd1 _05518_
+ sky130_fd_sc_hd__o21a_1
XFILLER_130_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__C net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10914__566 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__inv_2
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05850__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ net1673 _01620_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12602_ clknet_leaf_92_clk _02237_ net1086 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10808__460 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__inv_2
X_12533_ clknet_leaf_77_clk net3384 net1117 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06158__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05688__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08472__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05905__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ net2156 _02103_ net1081 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[957\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08064__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11415_ clknet_leaf_76_clk _01063_ net1123 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09421__A1 top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10425__77 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08224__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ net2087 _02034_ net1072 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[888\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10228_ net31 net654 net593 net3413 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__o22a_1
XANTENNA__06094__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10159_ _05617_ _05618_ net600 vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a21oi_1
Xhold2 top0.CPU.register.registers\[23\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05841__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07499__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08160__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06982__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07370_ _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__nand2_1
XANTENNA__08999__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06321_ net777 _02973_ _02975_ _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__06149__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ net168 net3228 net352 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__mux2_1
X_06252_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__inv_2
XANTENNA__07289__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10560__212 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__inv_2
Xhold402 top0.CPU.intMemAddr\[24\] vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08215__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857__509 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__inv_2
X_06183_ _02838_ _02839_ net786 vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
Xhold424 top0.CPU.register.registers\[327\] vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 top0.CPU.register.registers\[369\] vssd1 vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 top0.CPU.register.registers\[217\] vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09942_ _05434_ _05435_ _05429_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__a21oi_1
Xhold446 top0.CPU.register.registers\[372\] vssd1 vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 top0.CPU.register.registers\[774\] vssd1 vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 top0.CPU.register.registers\[344\] vssd1 vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 net907 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_2
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_4
XANTENNA__09176__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10601__253 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__inv_2
Xhold479 top0.CPU.register.registers\[65\] vssd1 vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_2
Xfanout937 net938 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_4
X_09873_ top0.CPU.internalMem.pcOut\[18\] net647 _05372_ vssd1 vssd1 vccd1 vccd1 _02195_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05764__C net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_A _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout926 net941 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08518__A3 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1113 net68 vssd1 vssd1 vccd1 vccd1 net3335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1102 top0.CPU.register.registers\[208\] vssd1 vssd1 vccd1 vccd1 net3324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 top0.CPU.register.registers\[199\] vssd1 vssd1 vccd1 vccd1 net3346 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ net172 net670 net312 net285 net2784 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1001_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net962 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
Xhold1157 top0.MISOtoMMIO\[4\] vssd1 vssd1 vccd1 vccd1 net3379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 top0.CPU.intMem_out\[6\] vssd1 vssd1 vccd1 vccd1 net3368 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net217 net619 net318 net295 net2436 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a32o_1
Xhold1135 top0.CPU.register.registers\[439\] vssd1 vssd1 vccd1 vccd1 net3357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 top0.MMIO.WBData_i\[13\] vssd1 vssd1 vccd1 vccd1 net3401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1168 top0.display.reading_flag vssd1 vssd1 vccd1 vccd1 net3390 sky130_fd_sc_hd__dlygate4sd3_1
X_07706_ net343 _03915_ _04355_ _04362_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__a31o_1
X_05967_ top0.CPU.register.registers\[772\] top0.CPU.register.registers\[804\] top0.CPU.register.registers\[836\]
+ top0.CPU.register.registers\[868\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02624_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout461_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ net175 net691 net310 net298 net2995 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a32o_1
X_05898_ _02552_ _02553_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_49_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06388__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07637_ _04106_ _04127_ _04293_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ net531 _03317_ net470 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__mux2_1
X_09307_ top0.display.counter\[4\] top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 _04960_
+ sky130_fd_sc_hd__nor2_1
X_06519_ _03174_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09100__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ _02788_ _02789_ net528 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__a21oi_1
X_09238_ net769 top0.CPU.intMemAddr\[0\] net611 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o21a_1
XANTENNA__09403__A1 top0.MMIO.WBData_i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ net194 net674 _04847_ net249 net3258 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a32o_1
XANTENNA__06560__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net1872 _01819_ net961 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[673\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09167__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold980 top0.CPU.register.registers\[278\] vssd1 vssd1 vccd1 vccd1 net3202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 top0.CPU.register.registers\[385\] vssd1 vssd1 vccd1 vccd1 net3213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07717__A1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ _05487_ _05490_ _05500_ net240 vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a31o_1
XANTENNA__08914__B1 _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328__980 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__inv_2
X_11964_ net1656 _01603_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09162__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06379__S1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11895_ net1587 _01534_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[388\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08693__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05900__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ net2208 _02155_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1009\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12447_ net2139 _02086_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[940\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09618__A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06741__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__A0 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ net2070 _02017_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06313__Y _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09158__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ _03525_ _03526_ net761 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
XANTENNA__06067__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05821_ top0.CPU.register.registers\[914\] top0.CPU.register.registers\[946\] top0.CPU.register.registers\[978\]
+ top0.CPU.register.registers\[1010\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02478_
+ sky130_fd_sc_hd__mux4_1
X_08540_ net194 net675 net401 net364 net2489 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a32o_1
X_05752_ _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__inv_2
X_08471_ net197 net622 net404 net371 net2412 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a32o_1
X_05683_ top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__inv_2
XANTENNA__06144__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080__732 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07422_ _03952_ _03982_ net478 vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__mux2_1
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05820__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__A1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07353_ net481 _03788_ _03832_ _04008_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o31a_1
X_11121__773 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10243__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07284_ _03562_ _03571_ _03573_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a21o_1
X_06304_ net580 _02952_ _02960_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__nor3_1
XANTENNA__06447__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09023_ _04548_ net613 _04803_ net352 net3296 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__a32o_1
X_06235_ top0.CPU.register.registers\[536\] top0.CPU.register.registers\[568\] top0.CPU.register.registers\[600\]
+ top0.CPU.register.registers\[632\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02892_
+ sky130_fd_sc_hd__mux4_1
Xhold210 top0.CPU.register.registers\[417\] vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout307_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07947__B2 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06166_ top0.CPU.register.registers\[16\] top0.CPU.register.registers\[48\] top0.CPU.register.registers\[80\]
+ top0.CPU.register.registers\[112\] net844 net809 vssd1 vssd1 vccd1 vccd1 _02823_
+ sky130_fd_sc_hd__mux4_1
Xhold243 top0.CPU.register.registers\[99\] vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 top0.CPU.register.registers\[704\] vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 top0.CPU.register.registers\[320\] vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_06097_ top0.CPU.register.registers\[780\] top0.CPU.register.registers\[812\] top0.CPU.register.registers\[844\]
+ top0.CPU.register.registers\[876\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02754_
+ sky130_fd_sc_hd__mux4_1
XFILLER_116_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold254 top0.CPU.register.registers\[939\] vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 top0.CPU.register.registers\[359\] vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 top0.CPU.register.registers\[103\] vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08151__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 top0.CPU.register.registers\[698\] vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 _04636_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
Xfanout723 _02390_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_113_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09925_ net585 _02456_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nor2_1
XANTENNA__09149__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 net704 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
Xhold298 top0.CPU.register.registers\[288\] vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout676_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 _02349_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_8
Xfanout767 net3435 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_2
X_09856_ _05353_ _05354_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout745 net746 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net759 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
XANTENNA__05805__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08578__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05791__A top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08807_ net671 _04739_ net286 net2663 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__a22o_1
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout843_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ _02768_ _04583_ net587 vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__mux2_1
XFILLER_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06999_ net745 _03655_ _03644_ _03648_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08124__A1 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985__637 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__inv_2
X_08738_ _04680_ net307 net293 net2552 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a22o_1
XFILLER_54_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _04661_ net307 net297 net3357 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ net1372 _01319_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[173\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07883__B1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07511__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06533__S1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12301_ net1993 _01940_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879__531 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__inv_2
X_12232_ net1924 _01871_ net1077 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[725\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net1855 _01802_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[656\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06297__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__A3 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ net1786 _01733_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09560__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06374__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11064__716 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__inv_2
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ net1639 _01586_ net1070 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[440\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08666__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105__757 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__inv_2
X_11878_ net1570 _01517_ net1129 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[371\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08418__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10225__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06429__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06524__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09091__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06020_ top0.CPU.register.registers\[390\] top0.CPU.register.registers\[422\] top0.CPU.register.registers\[454\]
+ top0.CPU.register.registers\[486\] net832 net798 vssd1 vssd1 vccd1 vccd1 _02677_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_130_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07929__B2 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08051__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ _04088_ net232 net227 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__and3_1
X_09710_ _05220_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__nand2_1
X_06922_ _03131_ _03151_ _03152_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__o21a_1
XANTENNA__09551__A0 top0.CPU.control.funct7\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672__324 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__inv_2
X_06853_ top0.CPU.register.registers\[650\] top0.CPU.register.registers\[682\] top0.CPU.register.registers\[714\]
+ top0.CPU.register.registers\[746\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03510_
+ sky130_fd_sc_hd__mux4_1
X_09641_ _02787_ _05154_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__nor2_1
XANTENNA__10161__A1 _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05804_ top0.CPU.register.registers\[787\] top0.CPU.register.registers\[819\] top0.CPU.register.registers\[851\]
+ top0.CPU.register.registers\[883\] net856 net821 vssd1 vssd1 vccd1 vccd1 _02461_
+ sky130_fd_sc_hd__mux4_1
X_10713__365 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__inv_2
X_09572_ _05117_ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__nand2b_1
X_06784_ _03439_ _03440_ net765 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__mux2_1
X_05735_ top0.CPU.decoder.instruction\[11\] net946 net575 net722 vssd1 vssd1 vccd1
+ vccd1 _02392_ sky130_fd_sc_hd__nand4_1
X_08523_ _04708_ net397 net362 net3031 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a22o_1
XANTENNA__08106__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07314__C1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08657__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net948 net545 _04671_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__or3_4
XANTENNA__07865__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout424_A _04689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08409__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07405_ net525 net524 net469 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__mux2_1
X_08385_ net157 net701 net386 net381 net2715 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a32o_1
XANTENNA__10216__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08861__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ net526 _03519_ net469 vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__mux2_1
XANTENNA__09082__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09006_ _04481_ net3192 net352 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ net480 _03923_ _03921_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06840__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ net343 _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__nand2_1
X_06218_ top0.CPU.register.registers\[790\] top0.CPU.register.registers\[822\] top0.CPU.register.registers\[854\]
+ top0.CPU.register.registers\[886\] net838 net803 vssd1 vssd1 vccd1 vccd1 _02875_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout793_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06149_ top0.CPU.register.registers\[273\] top0.CPU.register.registers\[305\] top0.CPU.register.registers\[337\]
+ top0.CPU.register.registers\[369\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02806_
+ sky130_fd_sc_hd__mux4_1
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_132_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout542 net544 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
Xfanout531 _03301_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_2
Xfanout520 _03656_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09542__A0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ top0.CPU.internalMem.pcOut\[21\] _05394_ net239 vssd1 vssd1 vccd1 vccd1 _05405_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__08345__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 net567 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
Xfanout597 net599 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_2
X_09839_ _05320_ _05330_ _05340_ _05339_ _05329_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a32oi_4
XANTENNA__08896__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 net588 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09721__A top0.CPU.control.funct7\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11801_ net1493 _01440_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06108__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08648__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11732_ net1424 _01371_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[225\]
+ sky130_fd_sc_hd__dfrtp_1
X_11663_ net1355 _01302_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09073__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11594_ net1286 _01233_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08281__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05696__A top0.MMIO.WBData_i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08072__A _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net1907 _01854_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[708\]
+ sky130_fd_sc_hd__dfrtp_1
X_12146_ net1838 _01785_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[639\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656__308 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__inv_2
XANTENNA__06304__B _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07119__C net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09533__A0 top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ net1769 _01716_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[570\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08887__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06993__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08170_ net222 net614 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__and2_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07075__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09064__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__inv_2
X_11192__844 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08811__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_121_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09521__A_N _05100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07052_ _02342_ net943 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__and2_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__09221__C1 top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06003_ top0.CPU.register.registers\[135\] top0.CPU.register.registers\[167\] top0.CPU.register.registers\[199\]
+ top0.CPU.register.registers\[231\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02660_
+ sky130_fd_sc_hd__mux4_1
X_11233__885 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__inv_2
XANTENNA__08575__A1 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05893__X _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10386__38 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__inv_2
XANTENNA__09119__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07954_ top0.CPU.intMem_out\[11\] net628 _04588_ _04590_ vssd1 vssd1 vccd1 vccd1
+ _04591_ sky130_fd_sc_hd__a22o_1
X_07885_ top0.CPU.internalMem.pcOut\[22\] net641 net635 _04532_ vssd1 vssd1 vccd1
+ vccd1 _04533_ sky130_fd_sc_hd__o211a_2
X_06905_ _03385_ _03407_ _03409_ _03561_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_52_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06836_ _03491_ _03492_ net760 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__mux2_1
X_09624_ _05150_ _02697_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout374_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06433__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06984__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06767_ _03420_ _03421_ _03423_ _03422_ net872 net752 vssd1 vssd1 vccd1 vccd1 _03424_
+ sky130_fd_sc_hd__mux4_2
X_09555_ net942 net943 net945 _04216_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__nand4_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06884__B net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _02353_ net148 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__nand2_1
X_08506_ net194 net686 net401 net368 net2719 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a32o_1
X_05718_ _02372_ _02374_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__nand2_2
XANTENNA__07332__Y _03989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08157__A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06698_ _03351_ _03354_ net866 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__mux2_1
XFILLER_24_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ net2880 _04566_ net375 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__mux2_1
XANTENNA__07302__A2 _03173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A top0.CPU.control.rs2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ net203 net707 net400 net383 net2615 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a32o_1
XANTENNA__09055__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ net3022 _04544_ net415 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
X_07319_ _03850_ _03949_ _03975_ _03747_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__o22a_1
XANTENNA__08802__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10841__493 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__inv_2
X_10330_ net2228 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ net3152 net117 net111 _05653_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a22o_1
XFILLER_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12000_ net1692 _01639_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[493\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ _04909_ net129 net122 net3167 net115 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a221o_1
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06041__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 _04798_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_6
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_4
Xfanout372 _04727_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_4
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout361 _04729_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06140__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08869__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout394 net397 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_2
XFILLER_62_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06975__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08097__A3 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ net1407 _01354_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[208\]
+ sky130_fd_sc_hd__dfrtp_1
X_12695_ clknet_leaf_91_clk _02330_ net1085 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ net1338 _01285_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[139\]
+ sky130_fd_sc_hd__dfrtp_1
X_11176__828 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__inv_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 nrst vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05697__Y _02355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ net1269 _01216_ net980 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[70\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_103_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_114_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap517 _03746_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_2
Xhold809 top0.CPU.register.registers\[573\] vssd1 vssd1 vccd1 vccd1 net3031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11217__869 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__inv_2
XANTENNA__08557__A1 _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12129_ net1821 _01768_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06415__S0 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07532__A2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ _03738_ _04156_ _04158_ _04326_ _04325_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__a221o_1
XANTENNA__07580__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06621_ _03274_ _03275_ _03277_ _03276_ net872 net751 vssd1 vssd1 vccd1 vccd1 _03278_
+ sky130_fd_sc_hd__mux4_2
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ _02338_ net630 _04973_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__and3_1
X_10784__436 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__inv_2
X_06552_ top0.CPU.register.registers\[785\] top0.CPU.register.registers\[817\] top0.CPU.register.registers\[849\]
+ top0.CPU.register.registers\[881\] net912 net878 vssd1 vssd1 vccd1 vccd1 _03209_
+ sky130_fd_sc_hd__mux4_1
X_09271_ _04865_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__or2_4
XFILLER_61_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06718__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08222_ net512 net197 net686 net423 net2394 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a32o_1
XANTENNA__08493__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06483_ top0.CPU.register.registers\[533\] top0.CPU.register.registers\[565\] top0.CPU.register.registers\[597\]
+ top0.CPU.register.registers\[629\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03140_
+ sky130_fd_sc_hd__mux4_1
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10825__477 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__inv_2
XANTENNA_fanout122_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ net209 net614 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__and2_1
X_08084_ net637 _04548_ net699 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and3_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07104_ _03129_ net447 net473 vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__mux2_1
X_07035_ _03690_ _03691_ net785 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__mux2_1
XANTENNA__08143__C net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678__330 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1031_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout491_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08986_ net193 net695 _04792_ net261 net3225 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__a32o_1
XANTENNA__06654__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ net717 _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__and2_1
X_10719__371 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__inv_2
XFILLER_84_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout756_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A3 top0.MMIO.WBData_i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07868_ _04411_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__and3_1
XANTENNA__06406__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08586__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06819_ _03474_ _03475_ net761 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ _03852_ _03886_ _04365_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or4_1
X_09607_ _05140_ _05143_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout923_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ net905 _05088_ net125 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06709__S1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ top0.MMIO.WBData_i\[28\] net145 net135 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ clknet_leaf_82_clk _01139_ net1108 vssd1 vssd1 vccd1 vccd1 top0.display.dataforOutput\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08484__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ net2172 _02119_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[973\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07883__A1_N _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ clknet_leaf_61_clk _01079_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08236__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__B1 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06798__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ _04851_ _04862_ _04935_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__and3b_1
XANTENNA__06135__A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net17 net654 net593 net3422 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__o22a_1
XFILLER_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1101 net1105 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_4
Xfanout1112 net1114 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
X_10175_ _05630_ _05631_ net600 vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a21oi_1
Xfanout1123 net1130 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout191 _04587_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
Xfanout180 _04600_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05773__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471__123 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__inv_2
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05913__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512__164 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__inv_2
XANTENNA__08475__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12678_ clknet_leaf_91_clk _02313_ net1084 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06744__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08227__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11629_ net1321 _01268_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08242__A3 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 top0.CPU.register.registers\[521\] vssd1 vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06789__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold606 top0.CPU.register.registers\[636\] vssd1 vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 top0.CPU.register.registers\[518\] vssd1 vssd1 vccd1 vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 top0.display.dataforOutput\[0\] vssd1 vssd1 vccd1 vccd1 net2850 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08260__A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ net152 net3042 net353 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__mux2_1
XANTENNA__07202__A1 _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05983_ top0.CPU.register.registers\[645\] top0.CPU.register.registers\[677\] top0.CPU.register.registers\[709\]
+ top0.CPU.register.registers\[741\] net849 net813 vssd1 vssd1 vccd1 vccd1 _02640_
+ sky130_fd_sc_hd__mux4_1
X_08771_ _04695_ net305 net289 net2751 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _03664_ _04366_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__nor2_1
XFILLER_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05823__S net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07653_ _03889_ _03908_ net346 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__mux2_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11345__997 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__inv_2
XANTENNA__06939__S1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06604_ _03255_ _03260_ net746 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__mux2_4
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09323_ net1199 top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 top0.display.sclk sky130_fd_sc_hd__or2_2
X_07584_ _04239_ _04240_ net450 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a21oi_1
X_06535_ _03188_ _03191_ net752 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__mux2_1
XANTENNA__08466__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09254_ _04912_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__or2_1
X_11198__850 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1079_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06466_ top0.CPU.register.registers\[148\] top0.CPU.register.registers\[180\] top0.CPU.register.registers\[212\]
+ top0.CPU.register.registers\[244\] net918 net884 vssd1 vssd1 vccd1 vccd1 _03123_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09030__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ top0.CPU.internalMem.state\[1\] top0.CPU.internalMem.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _04850_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08218__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08205_ net3230 net421 _04695_ net491 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout504_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08136_ net3117 net215 net429 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
X_06397_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__inv_2
XANTENNA__08233__A3 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239__891 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__inv_2
XANTENNA__06875__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ net2847 net433 _04656_ net498 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a22o_1
X_07018_ net872 _03674_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__and2_1
XANTENNA__09718__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout873_A top0.CPU.decoder.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455__107 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__inv_2
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _04661_ net554 _04785_ net261 net3252 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__a32o_1
XANTENNA__05850__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370__22 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__inv_2
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11980_ net1672 _01619_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_80_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12601_ clknet_leaf_92_clk _02236_ net1083 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08457__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12532_ clknet_leaf_77_clk net3373 net1117 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05969__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ net2155 _02102_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[956\]
+ sky130_fd_sc_hd__dfrtp_1
X_11414_ clknet_leaf_77_clk _01062_ net1130 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08064__B net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09421__A2 _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ net2086 _02033_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[887\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06152__X _02809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08080__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07395__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ net30 net654 net593 top0.MMIO.WBData_i\[6\] vssd1 vssd1 vccd1 vccd1 _02273_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06618__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06094__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032__684 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__inv_2
X_10158_ top0.display.delayctr\[26\] _05613_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 top0.CPU.register.registers\[25\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05841__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10089_ _04967_ _05548_ top0.display.delayctr\[12\] vssd1 vssd1 vccd1 vccd1 _05563_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08696__A0 _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08160__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06320_ net726 _02976_ net736 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06251_ _02906_ _02907_ net580 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_2
XANTENNA__08255__A _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_100_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07671__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09948__B1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06182_ top0.CPU.register.registers\[917\] top0.CPU.register.registers\[949\] top0.CPU.register.registers\[981\]
+ top0.CPU.register.registers\[1013\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02839_
+ sky130_fd_sc_hd__mux4_1
X_10896__548 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__inv_2
Xhold436 top0.CPU.register.registers\[941\] vssd1 vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06857__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold414 top0.CPU.register.registers\[487\] vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 top0.CPU.register.registers\[569\] vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 top0.CPU.register.registers\[565\] vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold447 top0.CPU.register.registers\[638\] vssd1 vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09941_ _05430_ _05390_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__nand2b_1
X_10640__292 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__inv_2
Xhold469 top0.CPU.register.registers\[570\] vssd1 vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 top0.CPU.register.registers\[993\] vssd1 vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout905 net907 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
X_10937__589 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__inv_2
Xfanout916 net919 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
Xfanout949 top0.CPU.decoder.instruction\[10\] vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_2
Xfanout938 net941 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_2
X_09872_ net236 _05367_ _05368_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a31o_1
XANTENNA__06609__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout927 net929 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_4
Xhold1114 top0.CPU.intMem_out\[31\] vssd1 vssd1 vccd1 vccd1 net3336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1103 top0.CPU.register.registers\[137\] vssd1 vssd1 vccd1 vccd1 net3325 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08823_ net176 net672 net318 net287 net2633 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__a32o_1
XFILLER_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1158 _02175_ vssd1 vssd1 vccd1 vccd1 net3380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1125 top0.CPU.register.registers\[105\] vssd1 vssd1 vccd1 vccd1 net3347 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net180 net621 net322 net295 net2470 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__a32o_1
Xhold1147 top0.display.delayctr\[8\] vssd1 vssd1 vccd1 vccd1 net3369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 top0.display.dataforOutput\[2\] vssd1 vssd1 vccd1 vccd1 net3358 sky130_fd_sc_hd__dlygate4sd3_1
X_05966_ _02621_ _02622_ net725 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1169 top0.CPU.intMem_out\[19\] vssd1 vssd1 vccd1 vccd1 net3391 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _04357_ _04361_ _04360_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__or3b_1
XANTENNA__09025__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ net3288 net299 _04742_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a21o_1
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout454_A _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
X_05897_ _02552_ _02553_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08687__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08149__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06999__A1_N net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ _04248_ _04260_ _04275_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nor4_1
XFILLER_14_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout621_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ _04092_ _04223_ net461 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout719_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06518_ _03157_ net535 vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__nand2_1
X_09306_ _03700_ net550 net142 vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07340__Y _03997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09237_ net769 _04632_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nand2_1
X_07498_ _02514_ net529 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07500__C net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06449_ top0.CPU.register.registers\[406\] top0.CPU.register.registers\[438\] top0.CPU.register.registers\[470\]
+ top0.CPU.register.registers\[502\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03106_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09403__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ top0.CPU.register.registers\[45\] net572 net558 vssd1 vssd1 vccd1 vccd1 _04847_
+ sky130_fd_sc_hd__o21a_1
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08611__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ top0.CPU.register.registers\[92\] net565 vssd1 vssd1 vccd1 vccd1 _04825_
+ sky130_fd_sc_hd__or2_1
X_08119_ net3115 _04539_ net432 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XFILLER_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07965__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold970 top0.CPU.register.registers\[159\] vssd1 vssd1 vccd1 vccd1 net3192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 top0.CPU.register.registers\[395\] vssd1 vssd1 vccd1 vccd1 net3203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold992 top0.CPU.register.registers\[132\] vssd1 vssd1 vccd1 vccd1 net3214 sky130_fd_sc_hd__dlygate4sd3_1
X_11016__668 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__inv_2
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10012_ _05487_ _05490_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__nand2_1
XANTENNA__12588__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08914__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07025__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08059__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ net1655 _01602_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[456\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_83_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08678__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11894_ net1586 _01533_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07350__A0 _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08693__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583__235 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__inv_2
XANTENNA__09642__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_8_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08850__A0 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ net2207 _02154_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1008\]
+ sky130_fd_sc_hd__dfrtp_1
X_12446_ net2138 _02085_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[939\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624__276 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__inv_2
XANTENNA__09618__B _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ net2069 _02016_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07405__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08602__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07956__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08241__C net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06323__A top0.CPU.control.funct7\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357__9 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__inv_2
XANTENNA__06067__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08905__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05820_ _02471_ _02475_ net579 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_4
XFILLER_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07016__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
X_10518__170 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__inv_2
X_05751_ net943 net942 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__and2b_2
XANTENNA__08669__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ net199 net620 net398 net371 net2293 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a32o_1
X_05682_ top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__inv_2
XANTENNA__06144__A1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A0 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07892__A1 top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07421_ net337 _03979_ _04077_ net476 _03743_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_102_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07352_ net480 _03788_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09094__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__A2 _02766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06303_ net776 _02959_ _02956_ net741 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_135_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07283_ _03916_ _03917_ _03938_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07644__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ top0.CPU.register.registers\[147\] net576 vssd1 vssd1 vccd1 vccd1 _04803_
+ sky130_fd_sc_hd__or2_1
X_06234_ top0.CPU.register.registers\[664\] top0.CPU.register.registers\[696\] top0.CPU.register.registers\[728\]
+ top0.CPU.register.registers\[760\] net838 net803 vssd1 vssd1 vccd1 vccd1 _02891_
+ sky130_fd_sc_hd__mux4_1
X_06165_ top0.CPU.register.registers\[144\] top0.CPU.register.registers\[176\] top0.CPU.register.registers\[208\]
+ top0.CPU.register.registers\[240\] net844 net809 vssd1 vssd1 vccd1 vccd1 _02822_
+ sky130_fd_sc_hd__mux4_1
Xhold200 top0.CPU.register.registers\[615\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 top0.CPU.register.registers\[449\] vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 top0.CPU.register.registers\[489\] vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07947__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold233 top0.CPU.intMemAddr\[30\] vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 top0.CPU.register.registers\[459\] vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
X_06096_ _02751_ _02752_ net734 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
XANTENNA__05958__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05958__A1 top0.CPU.decoder.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 top0.CPU.register.registers\[583\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 top0.CPU.register.registers\[743\] vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 top0.CPU.register.registers\[930\] vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 top0.CPU.register.registers\[364\] vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 top0.CPU.register.registers\[101\] vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ top0.CPU.internalMem.pcOut\[22\] net646 _05419_ vssd1 vssd1 vccd1 vccd1 _02199_
+ sky130_fd_sc_hd__o21ba_1
Xfanout702 net704 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08859__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout713 net716 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
Xfanout724 net727 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_4
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ top0.CPU.internalMem.pcOut\[16\] _05343_ _05345_ vssd1 vssd1 vccd1 vccd1
+ _05356_ sky130_fd_sc_hd__a21o_1
Xfanout757 net759 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
Xfanout746 net748 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_8
Xfanout735 net740 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
XANTENNA__07616__X _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 top0.CPU.control.rs2\[3\] vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_4
Xfanout768 top0.CPU.internalMem.pcOut\[2\] vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout571_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout669_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _04714_ net307 net285 net2739 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a22o_1
X_09786_ top0.CPU.internalMem.pcOut\[11\] net652 _05283_ _05292_ vssd1 vssd1 vccd1
+ vccd1 _02188_ sky130_fd_sc_hd__a22o_1
XFILLER_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06998_ _03651_ _03654_ net862 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_65_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
X_08737_ _04679_ net314 net294 net2607 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__a22o_1
X_05949_ top0.CPU.register.registers\[129\] top0.CPU.register.registers\[161\] top0.CPU.register.registers\[193\]
+ top0.CPU.register.registers\[225\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02606_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout836_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__B2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _04660_ net314 net298 net3108 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a22o_1
X_07619_ net462 _03338_ net339 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ net3151 net329 net305 _04511_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a22o_1
X_10567__219 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__inv_2
XANTENNA__09085__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07511__B _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net1992 _01939_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[793\]
+ sky130_fd_sc_hd__dfrtp_1
X_12231_ net1923 _01870_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[724\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07938__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ net1854 _01801_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06297__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12093_ net1785 _01732_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[586\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__C1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08899__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A1 top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__B1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
X_11946_ net1638 _01585_ net984 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[439\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07323__A0 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ net1569 _01516_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[370\]
+ sky130_fd_sc_hd__dfrtp_1
X_11144__796 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05980__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06318__A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08418__A3 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08823__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12429_ net2121 _02068_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038__690 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__inv_2
XANTENNA__08051__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ net718 net506 net219 net547 net2325 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a32o_1
X_06921_ _03562_ _03571_ _03575_ _03155_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a211o_1
XANTENNA__09000__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06852_ top0.CPU.register.registers\[778\] top0.CPU.register.registers\[810\] top0.CPU.register.registers\[842\]
+ top0.CPU.register.registers\[874\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03509_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06365__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ _05141_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__and2_1
XANTENNA__10303__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10161__A2 _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05803_ _02458_ _02459_ net734 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
X_09571_ _05115_ _05116_ top0.CPU.internalMem.pcOut\[1\] vssd1 vssd1 vccd1 vccd1 _05118_
+ sky130_fd_sc_hd__a21o_1
X_06783_ top0.CPU.register.registers\[270\] top0.CPU.register.registers\[302\] top0.CPU.register.registers\[334\]
+ top0.CPU.register.registers\[366\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03440_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12021__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
X_05734_ net955 net950 net953 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__nand3_1
X_08522_ _04707_ net405 net364 net2918 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a22o_1
XFILLER_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05831__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08657__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08453_ net2941 net153 net374 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout152_A _04528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07404_ _04059_ _04060_ net345 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__mux2_1
XANTENNA__09067__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05876__B1 _02532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08384_ net160 net701 net391 net381 net2416 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a32o_1
XANTENNA__08814__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07335_ _03719_ _03815_ _03926_ _03933_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__o32ai_4
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout417_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ _03859_ _03922_ net465 vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__mux2_1
X_09005_ _02396_ net613 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__nand2_2
X_06217_ _02872_ _02873_ net731 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__mux2_1
X_07197_ _03055_ _03057_ _03074_ _03667_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__a211o_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07059__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06148_ top0.CPU.register.registers\[401\] top0.CPU.register.registers\[433\] top0.CPU.register.registers\[465\]
+ top0.CPU.register.registers\[497\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02805_
+ sky130_fd_sc_hd__mux4_1
X_06079_ top0.CPU.register.registers\[781\] top0.CPU.register.registers\[813\] top0.CPU.register.registers\[845\]
+ top0.CPU.register.registers\[877\] net850 net815 vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout786_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952__604 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__inv_2
Xfanout510 net511 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_2
X_09907_ _05402_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__xnor2_1
XANTENNA__05800__A0 _02446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout532 _03279_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
Xfanout521 _03637_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout953_A top0.CPU.decoder.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_2
Xfanout565 net567 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_4
Xfanout554 net556 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
XFILLER_132_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout576 _02388_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_2
X_09838_ _05294_ _05299_ _05309_ _05321_ _05308_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a32o_1
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_2
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11087__739 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__inv_2
X_09769_ _05273_ _05275_ net241 vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06108__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ net1492 _01439_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08648__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07856__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11731_ net1423 _01370_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[224\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07241__B _03073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11662_ net1354 _01301_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[155\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09058__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ net1285 _01232_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08805__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08072__B net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12214_ net1906 _01853_ net1002 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[707\]
+ sky130_fd_sc_hd__dfrtp_1
X_12145_ net1837 _01784_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[638\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06304__C _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10695__347 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__inv_2
XFILLER_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12076_ net1768 _01715_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[569\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08336__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06347__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10736__388 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__inv_2
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_88_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09190__Y top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10589__241 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__inv_2
X_11929_ net1621 _01568_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[422\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08247__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09049__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06048__A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05953__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ net473 net522 _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_99_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08272__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07051_ _03038_ _03669_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__or3b_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
X_06002_ net778 _02654_ _02657_ _02658_ net773 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09772__A1 top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06586__B2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07953_ net562 _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__or2_1
X_07884_ top0.CPU.intMem_out\[22\] net627 _04531_ _02382_ vssd1 vssd1 vccd1 vccd1
+ _04532_ sky130_fd_sc_hd__a211o_1
X_06904_ _03426_ _03445_ _03487_ _03560_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__or4_1
XFILLER_68_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_52_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08327__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06835_ top0.CPU.register.registers\[523\] top0.CPU.register.registers\[555\] top0.CPU.register.registers\[587\]
+ top0.CPU.register.registers\[619\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03492_
+ sky130_fd_sc_hd__mux4_1
X_09623_ net3304 net605 net658 net3330 net136 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__a221o_1
XFILLER_68_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06433__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06766_ top0.CPU.register.registers\[15\] top0.CPU.register.registers\[47\] top0.CPU.register.registers\[79\]
+ top0.CPU.register.registers\[111\] net934 net900 vssd1 vssd1 vccd1 vccd1 _03423_
+ sky130_fd_sc_hd__mux4_1
XFILLER_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ _02342_ net944 _04216_ net943 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__or4b_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09485_ top0.MMIO.WBData_i\[14\] net148 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__and2_1
X_05717_ top0.CPU.Op\[6\] top0.CPU.Op\[3\] top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1
+ _02374_ sky130_fd_sc_hd__nor3b_2
XANTENNA_fanout534_A _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ _04703_ net394 net366 net2697 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a22o_1
X_06697_ _03352_ _03353_ net765 vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__mux2_1
XFILLER_51_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08157__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ net2996 _04561_ net373 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
X_08367_ _04649_ net407 net384 net2765 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ _02578_ _03923_ _03838_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08263__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ net3326 net204 net414 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__mux2_1
X_07249_ net455 _03810_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__or2_1
XANTENNA__08015__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ _04938_ _05138_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or2_1
XANTENNA__06899__Y _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _04905_ net129 net121 net3300 net115 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a221o_1
XANTENNA__06121__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_2
XANTENNA__08112__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout384 _04723_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_4
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_4
Xfanout362 _04729_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_6_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_4
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_83_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ net1406 _01353_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[207\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ clknet_leaf_91_clk _02329_ net1084 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05978__Y _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05935__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ net1337 _01284_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[138\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ net1268 _01215_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06360__S0 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06017__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ net1820 _01767_ net1044 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[621\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_97_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12059_ net1751 _01698_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[552\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06620_ top0.CPU.register.registers\[5\] top0.CPU.register.registers\[37\] top0.CPU.register.registers\[69\]
+ top0.CPU.register.registers\[101\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03277_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06415__S1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06179__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ net866 _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__nor2_1
X_09270_ _04893_ _04898_ _04925_ _04928_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__or4bb_2
X_06482_ top0.CPU.register.registers\[661\] top0.CPU.register.registers\[693\] top0.CPU.register.registers\[725\]
+ top0.CPU.register.registers\[757\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03139_
+ sky130_fd_sc_hd__mux4_1
X_08221_ net506 net199 net683 net423 net2656 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a32o_1
XANTENNA__05926__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200__852 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__inv_2
XANTENNA__06506__A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ net2921 net425 _04676_ net494 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a22o_1
X_10446__98 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_9_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
X_08083_ net2923 net435 _04664_ net498 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a22o_1
X_07103_ net450 _03758_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__nand2_2
XANTENNA__08796__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ top0.CPU.register.registers\[927\] top0.CPU.register.registers\[959\] top0.CPU.register.registers\[991\]
+ top0.CPU.register.registers\[1023\] net852 net817 vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06103__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1024_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ top0.CPU.register.registers\[173\] net572 net558 vssd1 vssd1 vccd1 vccd1
+ _04792_ sky130_fd_sc_hd__o21a_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09028__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06654__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ top0.CPU.internalMem.pcOut\[14\] net639 net636 _04575_ vssd1 vssd1 vccd1
+ vccd1 _04576_ sky130_fd_sc_hd__o211a_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08181__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06406__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ net3002 net546 net493 _04517_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
X_06818_ top0.CPU.register.registers\[13\] top0.CPU.register.registers\[45\] top0.CPU.register.registers\[77\]
+ top0.CPU.register.registers\[109\] net934 net900 vssd1 vssd1 vccd1 vccd1 _03475_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09271__B _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07798_ _04378_ _04388_ _04400_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__or4_1
X_09606_ net577 _05141_ _05142_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and3b_1
XFILLER_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09537_ net940 _05058_ net126 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ _03387_ _03403_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout916_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ net130 net133 _05052_ net599 net3407 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__o32a_1
XANTENNA__09681__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09399_ _04893_ _04897_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ net153 net693 net394 net378 net2270 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11430_ clknet_leaf_65_clk _01078_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08236__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958__610 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__inv_2
XANTENNA__06798__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ _04863_ _04935_ _04851_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a21o_1
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08539__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ net16 net655 net594 top0.MMIO.WBData_i\[22\] vssd1 vssd1 vccd1 vccd1 _02289_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07518__Y _04175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1105 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_2
Xfanout1113 net1114 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_2
X_10174_ top0.display.delayctr\[29\] _05626_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__nand2_1
Xfanout1124 net1130 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
Xfanout192 _04587_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
Xfanout170 _04615_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout181 _04600_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
XFILLER_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08172__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06722__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05930__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05908__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ clknet_leaf_91_clk _02312_ net1084 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
X_11628_ net1320 _01267_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08778__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 top0.CPU.register.registers\[319\] vssd1 vssd1 vccd1 vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11559_ net1251 _01198_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[52\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold618 top0.CPU.register.registers\[923\] vssd1 vssd1 vccd1 vccd1 net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 top0.CPU.register.registers\[757\] vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08260__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09643__Y _05169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08950__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751__403 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__inv_2
X_05982_ _02637_ _02638_ net730 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
X_08770_ _04694_ net305 net289 net2763 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__a22o_1
X_07721_ net343 _04368_ _04369_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a31o_1
X_07652_ net448 _04218_ _03842_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__a21o_1
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06603_ _03256_ _03257_ _03259_ _03258_ net869 net749 vssd1 vssd1 vccd1 vccd1 _03260_
+ sky130_fd_sc_hd__mux4_1
X_07583_ _03758_ _04238_ net517 vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a21o_1
X_06534_ _03189_ _03190_ net762 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
X_09322_ top0.display.dataforOutput\[15\] top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1
+ top0.bitDataTFT sky130_fd_sc_hd__or2_1
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_105_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09253_ top0.CPU.internalMem.pcOut\[6\] top0.CPU.addrControl _04913_ _04914_ vssd1
+ vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__a22o_1
X_06465_ _03118_ _03119_ _03120_ _03121_ net758 net750 vssd1 vssd1 vccd1 vccd1 _03122_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_138_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06572__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08218__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06396_ net859 _03046_ _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a21oi_4
X_09184_ net156 net671 net273 net248 net2469 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a32o_1
X_08204_ net208 net679 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_138_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ net2915 net167 net430 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08769__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06875__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__A2 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ net211 net690 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ top0.CPU.register.registers\[927\] top0.CPU.register.registers\[959\] top0.CPU.register.registers\[991\]
+ top0.CPU.register.registers\[1023\] net936 net903 vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_8_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08170__B net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06401__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10494__146 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__inv_2
X_08968_ top0.CPU.register.registers\[183\] net564 vssd1 vssd1 vccd1 vccd1 _04785_
+ sky130_fd_sc_hd__or2_1
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08899_ net718 net187 net276 net283 net2484 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__a32o_1
X_07919_ net713 net222 vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__B _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_27_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535__187 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__inv_2
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ clknet_leaf_89_clk _02235_ net1087 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12531_ clknet_leaf_76_clk _02170_ net1123 vssd1 vssd1 vccd1 vccd1 top0.MISOtoMMIO\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08209__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ net2154 _02101_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[955\]
+ sky130_fd_sc_hd__dfrtp_1
X_11413_ clknet_leaf_69_clk _01061_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09421__A3 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__B1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06315__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ net2085 _02032_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[886\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10226_ net29 net657 net596 top0.MMIO.WBData_i\[5\] vssd1 vssd1 vccd1 vccd1 _02272_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08080__B net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06618__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08393__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10157_ top0.display.delayctr\[26\] _05613_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__or2_1
Xhold4 top0.CPU.register.registers\[29\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08300__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10088_ top0.display.delayctr\[12\] _04967_ _05548_ vssd1 vssd1 vccd1 vccd1 _05562_
+ sky130_fd_sc_hd__or3_2
XANTENNA__07424__B _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09920__A top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07440__A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06250_ net774 net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08255__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07671__A2 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10416__68 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__inv_2
XANTENNA__06306__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06181_ top0.CPU.register.registers\[789\] top0.CPU.register.registers\[821\] top0.CPU.register.registers\[853\]
+ top0.CPU.register.registers\[885\] net839 net804 vssd1 vssd1 vccd1 vccd1 _02838_
+ sky130_fd_sc_hd__mux4_1
X_11271__923 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__inv_2
XANTENNA__07586__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 top0.CPU.register.registers\[751\] vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06857__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 top0.CPU.register.registers\[628\] vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 top0.CPU.register.registers\[867\] vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold459 top0.CPU.register.registers\[463\] vssd1 vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 top0.CPU.register.registers\[805\] vssd1 vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _05400_ _05412_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__nand2_1
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 top0.CPU.register.registers\[610\] vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
XFILLER_131_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09176__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312__964 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__inv_2
XANTENNA__06609__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout939 net941 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
X_09871_ net239 _05369_ _05370_ net652 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a31o_1
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
Xfanout917 net919 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_4
XANTENNA__08384__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ net218 net674 net322 net288 net2505 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a32o_1
Xhold1115 top0.CPU.register.registers\[210\] vssd1 vssd1 vccd1 vccd1 net3337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1104 top0.CPU.register.registers\[789\] vssd1 vssd1 vccd1 vccd1 net3326 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net183 net621 net323 net295 net2361 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a32o_1
Xhold1126 top0.CPU.register.registers\[234\] vssd1 vssd1 vccd1 vccd1 net3348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1148 top0.CPU.register.registers\[254\] vssd1 vssd1 vccd1 vccd1 net3370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05834__S net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1137 top0.display.dataforOutput\[6\] vssd1 vssd1 vccd1 vccd1 net3359 sky130_fd_sc_hd__dlygate4sd3_1
X_05965_ top0.CPU.register.registers\[516\] top0.CPU.register.registers\[548\] top0.CPU.register.registers\[580\]
+ top0.CPU.register.registers\[612\] net830 net795 vssd1 vssd1 vccd1 vccd1 _02622_
+ sky130_fd_sc_hd__mux4_1
Xhold1159 top0.CPU.intMem_out\[12\] vssd1 vssd1 vccd1 vccd1 net3381 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout182_A _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ net450 _04102_ _03849_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09884__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ top0.CPU.register.registers\[424\] net573 net219 net695 _04736_ vssd1 vssd1
+ vccd1 vccd1 _04742_ sky130_fd_sc_hd__o2111a_1
X_05896_ top0.CPU.decoder.instruction\[10\] _02448_ _02535_ net781 net583 vssd1 vssd1
+ vccd1 vccd1 _02553_ sky130_fd_sc_hd__a221oi_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ _04285_ _04291_ _04281_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a21bo_2
XANTENNA_fanout447_A _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07566_ net532 net530 net470 vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
X_06517_ _03157_ net535 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__or2_1
X_09305_ net944 _02517_ _03709_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_62_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09041__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09100__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ top0.CPU.addrControl _04895_ _04896_ _04894_ vssd1 vssd1 vccd1 vccd1 _04898_
+ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07497_ _04139_ _04146_ _04151_ _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout614_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06448_ top0.CPU.register.registers\[278\] top0.CPU.register.registers\[310\] top0.CPU.register.registers\[342\]
+ top0.CPU.register.registers\[374\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03105_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06379_ _03032_ _03033_ _03034_ _03035_ net762 net865 vssd1 vssd1 vccd1 vccd1 _03036_
+ sky130_fd_sc_hd__mux4_1
X_10920__572 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__inv_2
X_09167_ _04719_ net274 net248 net2792 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a22o_1
XANTENNA__08611__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _04691_ net556 _04824_ net252 net3138 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a32o_1
X_08118_ net3172 net206 net432 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
X_08049_ net511 net181 net708 net438 net2326 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a32o_1
XFILLER_135_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430__82 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__inv_2
Xhold982 top0.CPU.register.registers\[400\] vssd1 vssd1 vccd1 vccd1 net3204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold971 top0.CPU.register.registers\[825\] vssd1 vssd1 vccd1 vccd1 net3193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold960 top0.CPU.register.registers\[504\] vssd1 vssd1 vccd1 vccd1 net3182 sky130_fd_sc_hd__dlygate4sd3_1
X_10011_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__inv_2
XANTENNA__08375__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold993 top0.CPU.register.registers\[153\] vssd1 vssd1 vccd1 vccd1 net3215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_73_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08914__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08120__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07025__S1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__C net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ net1654 _01601_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12557__RESET_B net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11893_ net1585 _01532_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[386\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07350__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06575__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ net2206 _02153_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1007\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11255__907 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__inv_2
X_12445_ net2137 _02084_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[938\]
+ sky130_fd_sc_hd__dfrtp_1
X_12376_ net2068 _02015_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09158__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08366__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11149__801 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__inv_2
X_10209_ net2808 net123 net116 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a21o_1
XFILLER_121_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09193__Y top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05750_ net942 net943 net945 top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__or4b_1
XANTENNA__07016__S1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05681_ top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__inv_2
XANTENNA__07341__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07892__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07420_ _04034_ _04076_ net458 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
XANTENNA__06775__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863__515 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07170__A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07351_ net480 _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nand2_1
X_06302_ _02957_ _02958_ net726 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__mux2_1
X_10904__556 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07282_ _03916_ _03917_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o21a_1
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05896__Y _02553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06233_ _02497_ _02834_ _02870_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__nor4_1
X_09021_ net223 net3308 net349 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__mux2_1
X_06164_ net778 _02816_ net773 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__o21ai_1
Xhold201 top0.CPU.register.registers\[934\] vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold212 top0.CPU.register.registers\[613\] vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 top0.CPU.register.registers\[102\] vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 top0.CPU.register.registers\[356\] vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 top0.CPU.register.registers\[332\] vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
X_06095_ top0.CPU.register.registers\[524\] top0.CPU.register.registers\[556\] top0.CPU.register.registers\[588\]
+ top0.CPU.register.registers\[620\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02752_
+ sky130_fd_sc_hd__mux4_1
Xhold278 top0.CPU.register.registers\[874\] vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 top0.CPU.register.registers\[557\] vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 top0.CPU.register.registers\[425\] vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold289 top0.CPU.register.registers\[744\] vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net238 _05415_ _05418_ _05110_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__o22a_1
Xfanout703 net704 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_2
Xfanout714 net716 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09149__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__inv_2
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_8
Xfanout725 net727 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_4
Xfanout736 net740 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout397_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
X_08805_ _04713_ net314 net286 net2874 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold1212_A top0.CPU.intMem_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ _05290_ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__or2_1
X_06997_ _03652_ _03653_ net756 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout564_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ _04678_ net305 net293 net2601 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__a22o_1
X_05948_ _02601_ _02604_ net776 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05879_ top0.CPU.decoder.instruction\[10\] _02448_ _02535_ net781 vssd1 vssd1 vccd1
+ vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08667_ _04659_ net306 net297 net2917 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a22o_1
XANTENNA__06766__S0 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09609__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ net344 _04272_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout829_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ net2928 net329 net307 _04505_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _04204_ _04205_ _04153_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__A2 _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10647__299 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__inv_2
X_09219_ top0.CPU.intMemAddr\[12\] top0.CPU.intMemAddr\[11\] top0.CPU.intMemAddr\[21\]
+ top0.CPU.intMemAddr\[16\] vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net1922 _01869_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[723\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07079__X _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08596__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08115__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07239__B _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ net1853 _01800_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[654\]
+ sky130_fd_sc_hd__dfrtp_1
X_12092_ net1784 _01731_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[585\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold790 top0.CPU.register.registers\[277\] vssd1 vssd1 vccd1 vccd1 net3012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08348__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08899__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09848__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550__202 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__inv_2
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ net1637 _01584_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[438\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07323__A1 _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07874__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ net1568 _01515_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[369\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06509__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05980__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12428_ net2120 _02067_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ net2051 _01998_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[852\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06920_ _03155_ _03246_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__or2_1
XANTENNA__08339__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06851_ top0.CPU.register.registers\[906\] top0.CPU.register.registers\[938\] top0.CPU.register.registers\[970\]
+ top0.CPU.register.registers\[1002\] net933 net899 vssd1 vssd1 vccd1 vccd1 _03508_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06996__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05802_ top0.CPU.register.registers\[531\] top0.CPU.register.registers\[563\] top0.CPU.register.registers\[595\]
+ top0.CPU.register.registers\[627\] net856 net821 vssd1 vssd1 vccd1 vccd1 _02459_
+ sky130_fd_sc_hd__mux4_1
X_09570_ top0.CPU.internalMem.pcOut\[1\] _05115_ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_
+ sky130_fd_sc_hd__and3_1
X_06782_ top0.CPU.register.registers\[398\] top0.CPU.register.registers\[430\] top0.CPU.register.registers\[462\]
+ top0.CPU.register.registers\[494\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03439_
+ sky130_fd_sc_hd__mux4_1
X_08521_ net151 net675 net405 net363 net2711 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a32o_1
X_05733_ net954 net950 net952 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__and3_1
XANTENNA__08106__A3 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08708__B net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ net3062 net159 net373 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07403_ net537 net536 net447 _03129_ net467 net459 vssd1 vssd1 vccd1 vccd1 _04060_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05876__B2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ net166 net705 net389 net381 net2316 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a32o_1
XANTENNA__07617__A2 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _03809_ _03823_ net479 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07265_ net538 net521 net473 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1054_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ top0.CPU.decoder.instruction\[11\] _04725_ vssd1 vssd1 vccd1 vccd1 _04797_
+ sky130_fd_sc_hd__nor2_4
X_11318__970 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__inv_2
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06216_ top0.CPU.register.registers\[534\] top0.CPU.register.registers\[566\] top0.CPU.register.registers\[598\]
+ top0.CPU.register.registers\[630\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02873_
+ sky130_fd_sc_hd__mux4_1
X_07196_ _03074_ _03667_ _03055_ _03057_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_57_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10991__643 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__inv_2
X_06147_ _02802_ _02803_ net726 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
X_06078_ top0.CPU.register.registers\[909\] top0.CPU.register.registers\[941\] top0.CPU.register.registers\[973\]
+ top0.CPU.register.registers\[1005\] net850 net815 vssd1 vssd1 vccd1 vccd1 _02735_
+ sky130_fd_sc_hd__mux4_1
XFILLER_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09555__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_A top0.CPU.control.rs2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net515 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
X_10400__52 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__inv_2
X_09906_ _05387_ _05392_ _05386_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a21bo_1
Xfanout533 _03241_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout681_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
Xfanout522 _03617_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1107_X net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout544 _02433_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
Xfanout599 _04948_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_2
X_09837_ top0.CPU.internalMem.pcOut\[15\] _05328_ _05318_ vssd1 vssd1 vccd1 vccd1
+ _05339_ sky130_fd_sc_hd__a21o_1
Xfanout577 _04936_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
Xfanout588 _02417_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08345__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A_N net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09768_ _05273_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__or2_1
XANTENNA__08750__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ net180 net3196 net359 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__mux2_1
XANTENNA__07803__A _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ net1422 _01369_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[223\]
+ sky130_fd_sc_hd__dfrtp_1
X_09699_ top0.CPU.internalMem.pcOut\[5\] _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__xor2_1
XANTENNA__07081__Y _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08502__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ net1353 _01300_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[154\]
+ sky130_fd_sc_hd__dfrtp_1
X_11592_ net1284 _01231_ net1070 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08033__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ net1905 _01852_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[706\]
+ sky130_fd_sc_hd__dfrtp_1
X_11070__722 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__inv_2
X_12144_ net1836 _01783_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10128__B1 _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ net1767 _01714_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[568\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11111__763 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08741__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06978__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07713__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ net1620 _01567_ net1030 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[421\]
+ sky130_fd_sc_hd__dfrtp_1
X_11859_ net1551 _01498_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[352\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05953__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07050_ _03704_ _03706_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08272__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__X _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08009__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06001_ net725 _02655_ net737 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a21o_1
X_10975__627 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__inv_2
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__09772__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08980__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07952_ _03989_ net234 net229 vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and3_1
XANTENNA__10119__B1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ _02386_ _02871_ _04476_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__a2bb2o_1
X_06903_ _03505_ _03521_ _03542_ _03559_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_52_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06834_ top0.CPU.register.registers\[651\] top0.CPU.register.registers\[683\] top0.CPU.register.registers\[715\]
+ top0.CPU.register.registers\[747\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03491_
+ sky130_fd_sc_hd__mux4_1
X_09622_ _02715_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nor2_1
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08732__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ top0.CPU.control.funct7\[6\] _05061_ net126 vssd1 vssd1 vccd1 vccd1 _01122_
+ sky130_fd_sc_hd__mux2_1
X_10869__521 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__inv_2
X_08504_ net197 net686 net404 net367 net2706 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a32o_1
X_06765_ top0.CPU.register.registers\[143\] top0.CPU.register.registers\[175\] top0.CPU.register.registers\[207\]
+ top0.CPU.register.registers\[239\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03422_
+ sky130_fd_sc_hd__mux4_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09484_ top0.MMIO.WBData_i\[0\] net139 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__or2_1
X_05716_ top0.CPU.Op\[2\] top0.CPU.Op\[1\] top0.CPU.Op\[0\] vssd1 vssd1 vccd1 vccd1
+ _02373_ sky130_fd_sc_hd__nand3b_1
XFILLER_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06239__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ top0.CPU.register.registers\[256\] top0.CPU.register.registers\[288\] top0.CPU.register.registers\[320\]
+ top0.CPU.register.registers\[352\] net921 net887 vssd1 vssd1 vccd1 vccd1 _03353_
+ sky130_fd_sc_hd__mux4_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ net2795 _04555_ net375 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout527_A _03463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08366_ _04648_ net392 net382 net3105 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08799__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ _02533_ _03504_ net339 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08263__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ net3067 net206 net414 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__mux2_1
X_07248_ net455 _03813_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout896_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08015__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__inv_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054__706 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__inv_2
XANTENNA__09763__A2 _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _04901_ net129 net121 net3361 net115 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a221o_1
XANTENNA__06026__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377__29 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__inv_2
XFILLER_2_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06121__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 net332 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_8
Xfanout341 _03741_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout352 _04798_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_4
Xfanout374 net376 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_6
XANTENNA__05880__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_6_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout385 net387 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_2
XFILLER_74_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07533__A _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ clknet_leaf_93_clk _02328_ net1081 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XFILLER_42_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11713_ net1405 _01352_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[206\]
+ sky130_fd_sc_hd__dfrtp_1
X_11644_ net1336 _01283_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[137\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05935__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10662__314 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__inv_2
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
X_11575_ net1267 _01214_ net970 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08254__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06360__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367__1019 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__inv_2
X_10703__355 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__inv_2
XANTENNA__06017__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08303__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net1819 _01766_ net1097 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[620\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05871__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ net1750 _01697_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[551\]
+ sky130_fd_sc_hd__dfrtp_1
X_10391__43 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__inv_2
XANTENNA__06059__A2_N _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08714__A0 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06550_ _03205_ _03206_ net758 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06179__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06481_ net753 _03137_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or2_1
XANTENNA__08493__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08220_ net3223 net421 _04702_ net494 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a22o_1
XANTENNA__05926__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08151_ net210 net617 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__and2_1
XANTENNA__10052__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ net223 net692 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__and2_1
X_07102_ _02428_ _02431_ _03710_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__or3_2
XANTENNA__08796__A3 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07033_ top0.CPU.register.registers\[799\] top0.CPU.register.registers\[831\] top0.CPU.register.registers\[863\]
+ top0.CPU.register.registers\[895\] net852 net817 vssd1 vssd1 vccd1 vccd1 _03690_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06008__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06103__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ _04667_ net274 net262 net2745 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1017_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07935_ _04476_ _04573_ _04574_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a21o_1
XANTENNA__05862__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ _02634_ _05007_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__nor2_1
XFILLER_56_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_3_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06668__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ net716 net208 vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__and2_1
XANTENNA__09044__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06817_ top0.CPU.register.registers\[141\] top0.CPU.register.registers\[173\] top0.CPU.register.registers\[205\]
+ top0.CPU.register.registers\[237\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03474_
+ sky130_fd_sc_hd__mux4_1
X_07797_ _04411_ _04421_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__or3_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06192__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ net3398 _05065_ net126 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
X_06748_ _03387_ _03403_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nor2_1
X_09467_ top0.MMIO.WBData_i\[27\] net145 net135 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__o21a_1
XANTENNA__09130__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08418_ net159 net690 net386 net377 net2592 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08484__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06679_ _03334_ _03335_ net756 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__mux2_1
X_09398_ _04918_ _04920_ _04927_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_22_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08349_ net714 net213 net391 net410 net2519 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a32o_1
XFILLER_138_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08787__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ net2419 net117 net111 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a21o_1
X_10242_ net15 net657 net596 top0.MMIO.WBData_i\[21\] vssd1 vssd1 vccd1 vccd1 _02288_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07528__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__A1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08123__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1103 net1105 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08944__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ top0.display.delayctr\[29\] _05626_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__or2_1
XANTENNA__05853__S0 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1125 net1130 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_2
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_2
Xfanout182 _04596_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout171 _04611_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
Xfanout160 net163 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
Xfanout193 net195 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XANTENNA__06578__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08172__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182__834 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__inv_2
XFILLER_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08078__B net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09121__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06030__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223__875 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__inv_2
XANTENNA__08475__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05908__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ clknet_leaf_81_clk _02311_ net1112 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__10129__A _02850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11627_ net1319 _01266_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_11558_ net1250 _01197_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold608 top0.CPU.register.registers\[920\] vssd1 vssd1 vccd1 vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ clknet_leaf_79_clk top0.display.next_state\[1\] net1111 vssd1 vssd1 vccd1
+ vccd1 top0.display.state\[1\] sky130_fd_sc_hd__dfrtp_1
Xhold619 top0.CPU.register.registers\[337\] vssd1 vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06097__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08935__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05844__S0 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06410__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10790__442 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__inv_2
X_05981_ top0.CPU.register.registers\[773\] top0.CPU.register.registers\[805\] top0.CPU.register.registers\[837\]
+ top0.CPU.register.registers\[869\] net848 net814 vssd1 vssd1 vccd1 vccd1 _02638_
+ sky130_fd_sc_hd__mux4_1
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07720_ _04376_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__inv_2
XANTENNA__06488__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _03562_ _03571_ _03573_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831__483 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__inv_2
XANTENNA__07910__B2 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ top0.CPU.register.registers\[7\] top0.CPU.register.registers\[39\] top0.CPU.register.registers\[71\]
+ top0.CPU.register.registers\[103\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03259_
+ sky130_fd_sc_hd__mux4_1
X_07582_ net489 _04237_ _04238_ _03837_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__o2bb2a_1
X_06533_ top0.CPU.register.registers\[18\] top0.CPU.register.registers\[50\] top0.CPU.register.registers\[82\]
+ top0.CPU.register.registers\[114\] net931 net897 vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__mux4_1
X_09321_ net662 _04959_ _04972_ net603 vssd1 vssd1 vccd1 vccd1 top0.display.next_state\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_105_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08466__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ net769 top0.CPU.intMemAddr\[6\] net610 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__o21a_1
X_06464_ top0.CPU.register.registers\[532\] top0.CPU.register.registers\[564\] top0.CPU.register.registers\[596\]
+ top0.CPU.register.registers\[628\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03121_
+ sky130_fd_sc_hd__mux4_1
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06572__S1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06395_ net746 _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__and2_1
X_08203_ net3259 net421 _04694_ net491 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
X_09183_ net157 net668 _04849_ net247 net3302 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a32o_1
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08134_ net2878 net173 net430 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ net3147 net436 _04655_ net503 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a22o_1
XANTENNA__09179__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ top0.CPU.register.registers\[799\] top0.CPU.register.registers\[831\] top0.CPU.register.registers\[863\]
+ top0.CPU.register.registers\[895\] net937 net903 vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09039__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07635__X _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166__818 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__inv_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A top0.CPU.decoder.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ _04660_ net275 net262 net3036 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__a22o_1
X_08898_ net723 net190 net280 net284 net2289 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__a32o_1
X_07918_ top0.CPU.internalMem.pcOut\[17\] net639 net633 _04560_ vssd1 vssd1 vccd1
+ vccd1 _04561_ sky130_fd_sc_hd__o211a_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07849_ net563 _04500_ _04501_ net626 vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o211a_1
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_67_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08154__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207__859 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__inv_2
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366__1018 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__inv_2
XANTENNA__06260__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _05092_ _05093_ _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__and3_1
XANTENNA__09103__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08457__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ net2222 _02169_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1023\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06012__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07530__B _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08209__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12461_ net2153 _02100_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[954\]
+ sky130_fd_sc_hd__dfrtp_1
X_11412_ clknet_leaf_77_clk _01060_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06861__S net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06315__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net2084 _02031_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08090__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06079__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ net28 net655 net594 net3322 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__o22a_1
XANTENNA__08917__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774__426 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__inv_2
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ _02942_ net551 net141 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__o21ai_1
Xhold5 top0.CPU.internalMem.load2Ct\[0\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
X_10361__13 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__inv_2
X_10087_ net3362 net665 net603 _05561_ _05161_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a221o_1
X_10815__467 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__inv_2
XANTENNA__09342__B1 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07424__C _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09920__B top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10668__320 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__inv_2
XFILLER_90_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06003__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12659_ clknet_leaf_66_clk _02294_ net1103 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10709__361 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__inv_2
XANTENNA__07120__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06306__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06180_ _02835_ _02836_ net732 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__mux2_1
Xhold416 top0.CPU.register.registers\[127\] vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 top0.CPU.register.registers\[453\] vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08271__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold427 top0.CPU.register.registers\[81\] vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold449 top0.CPU.register.registers\[634\] vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 top0.CPU.register.registers\[675\] vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout907 top0.CPU.decoder.instruction\[16\] vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_4
XANTENNA__08908__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09870_ top0.CPU.internalMem.pcOut\[18\] _05359_ vssd1 vssd1 vccd1 vccd1 _05370_
+ sky130_fd_sc_hd__or2_1
XANTENNA__10306__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout929 net938 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
X_08821_ net180 net674 net322 net287 net2616 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a32o_1
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_2
XANTENNA__08698__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold1105 net91 vssd1 vssd1 vccd1 vccd1 net3327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 top0.CPU.intMem_out\[17\] vssd1 vssd1 vccd1 vccd1 net3360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 top0.CPU.intMem_out\[30\] vssd1 vssd1 vccd1 vccd1 net3349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 net38 vssd1 vssd1 vccd1 vccd1 net3338 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net187 net619 net321 net295 net2760 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__a32o_1
Xhold1149 top0.display.delayctr\[14\] vssd1 vssd1 vccd1 vccd1 net3371 sky130_fd_sc_hd__dlygate4sd3_1
X_05964_ top0.CPU.register.registers\[644\] top0.CPU.register.registers\[676\] top0.CPU.register.registers\[708\]
+ top0.CPU.register.registers\[740\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02621_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06490__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ net179 net696 net322 net299 net2467 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_107_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07703_ net486 _03720_ _03816_ _04358_ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o311a_1
X_05895_ _02544_ _02550_ net580 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08687__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ _03758_ _04286_ _04288_ _04290_ _03840_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a311o_1
XANTENNA__06242__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07631__A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ net245 _04219_ _04220_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__o211a_1
X_06516_ net748 _03172_ _03165_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a21oi_4
X_09304_ net577 _04952_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_62_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1084_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07496_ _03960_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__and2_1
XFILLER_110_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09235_ top0.CPU.addrControl _04895_ _04896_ _04894_ vssd1 vssd1 vccd1 vccd1 _04897_
+ sky130_fd_sc_hd__o31a_1
X_06447_ net753 _03099_ net859 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout607_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09166_ net196 net676 net279 net249 net2641 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a32o_1
X_06378_ top0.CPU.register.registers\[286\] top0.CPU.register.registers\[318\] top0.CPU.register.registers\[350\]
+ top0.CPU.register.registers\[382\] net937 net901 vssd1 vssd1 vccd1 vccd1 _03035_
+ sky130_fd_sc_hd__mux4_1
X_10461__113 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__inv_2
XANTENNA__09277__B _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ top0.CPU.register.registers\[93\] net569 vssd1 vssd1 vccd1 vccd1 _04824_
+ sky130_fd_sc_hd__or2_1
X_08117_ net2810 _04528_ net429 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
X_08048_ net509 net184 net708 net438 net2618 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a32o_1
XANTENNA__06622__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout976_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 top0.CPU.register.registers\[924\] vssd1 vssd1 vccd1 vccd1 net3183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold950 top0.CPU.register.registers\[918\] vssd1 vssd1 vccd1 vccd1 net3172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 top0.CPU.register.registers\[793\] vssd1 vssd1 vccd1 vccd1 net3194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold983 top0.CPU.register.registers\[143\] vssd1 vssd1 vccd1 vccd1 net3205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 top0.CPU.register.registers\[136\] vssd1 vssd1 vccd1 vccd1 net3216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ _05497_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10502__154 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__inv_2
XFILLER_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09999_ _05487_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07806__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08914__A3 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__A1 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ net1653 _01600_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[454\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07350__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net1584 _01531_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[385\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12597__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ net2205 _02152_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1006\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294__946 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__inv_2
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12444_ net2136 _02083_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[937\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ net2067 _02014_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08602__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08091__B net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11335__987 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__inv_2
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08311__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188__840 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__inv_2
XANTENNA__08905__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ net2843 net117 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__and2_1
XFILLER_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10139_ top0.display.delayctr\[22\] net663 _05141_ _05599_ _05602_ vssd1 vssd1 vccd1
+ vccd1 _02231_ sky130_fd_sc_hd__a221o_1
XFILLER_95_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11408__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229__881 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__inv_2
XFILLER_75_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08669__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05680_ top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__inv_2
XANTENNA__07341__A2 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06775__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07170__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ _03053_ net538 net521 net520 net474 net465 vssd1 vssd1 vccd1 vccd1 _04007_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09094__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06301_ top0.CPU.register.registers\[27\] top0.CPU.register.registers\[59\] top0.CPU.register.registers\[91\]
+ top0.CPU.register.registers\[123\] net826 net793 vssd1 vssd1 vccd1 vccd1 _02958_
+ sky130_fd_sc_hd__mux4_1
X_07281_ _03931_ _03932_ _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__and4_1
X_10943__595 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__inv_2
X_09020_ net204 net2892 net350 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06232_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__inv_2
X_06163_ net737 _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__nor2_1
XANTENNA__09097__B net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08054__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 top0.CPU.register.registers\[929\] vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 top0.CPU.register.registers\[460\] vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 top0.CPU.register.registers\[845\] vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06536__A1_N net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold213 top0.CPU.register.registers\[868\] vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_11365__1017 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__inv_2
X_06094_ top0.CPU.register.registers\[652\] top0.CPU.register.registers\[684\] top0.CPU.register.registers\[716\]
+ top0.CPU.register.registers\[748\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02751_
+ sky130_fd_sc_hd__mux4_1
Xhold257 top0.CPU.register.registers\[719\] vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 top0.CPU.register.registers\[289\] vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 top0.CPU.register.registers\[963\] vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _05416_ _05417_ net646 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__o21a_1
Xhold279 top0.CPU.register.registers\[614\] vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout704 net712 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_2
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_2
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_113_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09853_ net587 _04557_ _05351_ top0.CPU.internalMem.pcOut\[17\] vssd1 vssd1 vccd1
+ vccd1 _05354_ sky130_fd_sc_hd__a211o_1
Xfanout748 _02346_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_A _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _05272_ _05276_ _05289_ net240 vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a31o_1
XFILLER_105_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout759 _02344_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07345__B _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ _04712_ net306 net285 net2794 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__a22o_1
XANTENNA__08109__A1 _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08735_ _04677_ net305 net293 net2583 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__a22o_1
X_06996_ top0.CPU.register.registers\[282\] top0.CPU.register.registers\[314\] top0.CPU.register.registers\[346\]
+ top0.CPU.register.registers\[378\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03653_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout557_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05947_ _02602_ _02603_ net782 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold1205_A top0.CPU.intMem_out\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05878_ _02376_ _02447_ _02450_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__nand3_4
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06215__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _04658_ net305 net297 net3122 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a22o_1
XANTENNA__06676__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09609__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07617_ _04264_ _04273_ _04271_ _04270_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__o211a_1
X_08597_ net2881 net329 net311 _04499_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _02831_ _04149_ _03241_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout724_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09085__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ _02908_ _03617_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__nor2_1
X_11022__674 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__inv_2
X_09218_ top0.CPU.intMemAddr\[23\] _04876_ _02337_ vssd1 vssd1 vccd1 vccd1 _04880_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08045__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09149_ _04708_ net556 _04843_ net248 net3229 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a32o_1
X_12160_ net1852 _01799_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__A0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ net1783 _01730_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[584\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold791 top0.CPU.register.registers\[539\] vssd1 vssd1 vccd1 vccd1 net3013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold780 top0.CPU.register.registers\[1017\] vssd1 vssd1 vccd1 vccd1 net3002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08131__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07020__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06206__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10886__538 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__inv_2
X_11944_ net1636 _01583_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[437\]
+ sky130_fd_sc_hd__dfrtp_1
X_11875_ net1567 _01514_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[368\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630__282 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09076__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927__579 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__inv_2
XANTENNA__08823__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09198__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09697__A_N _04127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ net2119 _02066_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[920\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09784__B1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12358_ net2050 _01997_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08051__A3 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12289_ net1981 _01928_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06693__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06350__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09000__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ _02730_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__xnor2_2
X_05801_ top0.CPU.register.registers\[659\] top0.CPU.register.registers\[691\] top0.CPU.register.registers\[723\]
+ top0.CPU.register.registers\[755\] net856 net821 vssd1 vssd1 vccd1 vccd1 _02458_
+ sky130_fd_sc_hd__mux4_1
XFILLER_83_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06996__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ net866 _03437_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__nor2_1
X_05732_ net955 net952 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__nand2_1
X_08520_ net948 _02400_ _04705_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__or3_4
XANTENNA__07181__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ net2788 net160 net373 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__mux2_1
XFILLER_51_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ net535 net534 _03221_ net533 net467 net459 vssd1 vssd1 vccd1 vccd1 _04059_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_34_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09067__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006__658 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__inv_2
X_08382_ net213 net702 net391 net382 net2593 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a32o_1
XANTENNA__08814__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08275__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ _03521_ _03968_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_124_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07264_ net345 _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__or2_1
X_06215_ top0.CPU.register.registers\[662\] top0.CPU.register.registers\[694\] top0.CPU.register.registers\[726\]
+ top0.CPU.register.registers\[758\] net837 net802 vssd1 vssd1 vccd1 vccd1 _02872_
+ sky130_fd_sc_hd__mux4_1
X_09003_ net156 net693 net273 net262 net2276 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1047_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ _03669_ _03786_ _03845_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A3 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06146_ top0.CPU.register.registers\[17\] top0.CPU.register.registers\[49\] top0.CPU.register.registers\[81\]
+ top0.CPU.register.registers\[113\] net826 net791 vssd1 vssd1 vccd1 vccd1 _02803_
+ sky130_fd_sc_hd__mux4_1
XFILLER_104_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06077_ net943 _02474_ _02472_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a21o_2
XANTENNA__09555__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06684__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_2
XFILLER_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09527__A0 top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__inv_2
Xfanout523 _03600_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_4
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _02400_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout534 _03193_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout556 _04754_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
X_10573__225 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__inv_2
X_09836_ _05226_ _05244_ _05245_ _05296_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a2111o_1
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_2
Xfanout567 _02388_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
XANTENNA__06761__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _05250_ _05252_ _05260_ _05262_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout841_A top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ _03632_ _03633_ _03634_ _03635_ net758 net863 vssd1 vssd1 vccd1 vccd1 _03636_
+ sky130_fd_sc_hd__mux4_1
X_08718_ net182 net3234 net359 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout939_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ top0.CPU.control.funct7\[0\] net632 _02453_ _05210_ vssd1 vssd1 vccd1 vccd1
+ _05211_ sky130_fd_sc_hd__a31o_1
XANTENNA__07803__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ net182 net708 net323 net303 net2523 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a32o_1
X_10614__266 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__inv_2
XANTENNA__06739__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07091__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__A _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09058__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11660_ net1352 _01299_ net968 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08266__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ net1283 _01230_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[84\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_115_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08805__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08281__A3 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10508__160 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__inv_2
XANTENNA__08569__A1 _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12212_ net1904 _01851_ net960 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[705\]
+ sky130_fd_sc_hd__dfrtp_1
X_12143_ net1835 _01782_ net997 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[636\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11753__RESET_B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06675__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ net1766 _01713_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06427__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06978__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__12541__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11927_ net1619 _01566_ net973 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[420\]
+ sky130_fd_sc_hd__dfrtp_1
X_11364__1016 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__inv_2
X_11858_ net1550 _01497_ net1053 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09049__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11789_ net1481 _01428_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[282\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_106_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10064__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06345__A top0.CPU.control.funct7\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06000_ net782 _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__and2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__06666__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557__209 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__inv_2
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ _02385_ net628 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nor2_4
XANTENNA__06586__A3 _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10119__A1 _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06902_ net524 _03557_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06991__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _04363_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07904__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06833_ _02533_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__xnor2_1
X_09621_ net577 _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__or2_1
XFILLER_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06764_ top0.CPU.register.registers\[399\] top0.CPU.register.registers\[431\] top0.CPU.register.registers\[463\]
+ top0.CPU.register.registers\[495\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03421_
+ sky130_fd_sc_hd__mux4_1
X_09552_ top0.CPU.control.funct7\[5\] _05067_ net126 vssd1 vssd1 vccd1 vccd1 _01121_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07940__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07623__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ net199 net687 net399 net367 net2598 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a32o_1
X_05715_ top0.CPU.Op\[2\] top0.CPU.Op\[1\] top0.CPU.Op\[0\] vssd1 vssd1 vccd1 vccd1
+ _02372_ sky130_fd_sc_hd__and3b_1
X_09483_ top0.MMIO.WBData_i\[26\] net137 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout255_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08496__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06695_ top0.CPU.register.registers\[384\] top0.CPU.register.registers\[416\] top0.CPU.register.registers\[448\]
+ top0.CPU.register.registers\[480\] net921 net887 vssd1 vssd1 vccd1 vccd1 _03352_
+ sky130_fd_sc_hd__mux4_1
X_08434_ net3139 _04548_ net376 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__mux2_1
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05711__X _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ _04647_ net396 net382 net2768 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
XANTENNA__08454__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _02534_ net526 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout422_A _04689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ net3020 net152 net413 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
X_11093__745 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__inv_2
X_07247_ net455 _03807_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ net490 net518 vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout791_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06657__S0 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06129_ _02782_ _02783_ _02784_ _02785_ net733 net780 vssd1 vssd1 vccd1 vccd1 _02786_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout889_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134__786 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__inv_2
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_4
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout364 _04729_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_8
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 net354 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_8
XANTENNA__05880__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _05320_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__and2_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07373__X _04030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout397 net408 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_4
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_2
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11712_ net1404 _01351_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[205\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11028__680 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__inv_2
X_12692_ clknet_leaf_93_clk _02327_ net1082 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11643_ net1335 _01282_ net1009 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[136\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_11574_ net1266 _01213_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06896__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10742__394 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__inv_2
XANTENNA__10306__C_N _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ net1818 _01765_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[619\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06104__S net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05871__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ net1749 _01696_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[550\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09911__A0 top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__10150__A _02924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06480_ _03135_ _03136_ net764 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_1
XFILLER_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05898__B _02553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08150_ net3207 net425 _04675_ net499 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a22o_1
X_07101_ _02423_ _02427_ _02430_ _03711_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__o211a_4
X_11077__729 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__inv_2
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08650__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06887__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08081_ net2943 net436 _04663_ net501 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
X_07032_ _03687_ _03688_ net730 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__mux2_1
XANTENNA__07525__A2_N _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08402__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ net196 net697 net278 net260 net2392 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__a32o_1
XANTENNA__09833__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ top0.CPU.intMem_out\[14\] net627 _02773_ net591 net642 vssd1 vssd1 vccd1
+ vccd1 _04574_ sky130_fd_sc_hd__a221o_1
XANTENNA__05862__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06949__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__B1 top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ top0.CPU.internalMem.pcOut\[25\] net638 net633 _04515_ vssd1 vssd1 vccd1
+ vccd1 _04516_ sky130_fd_sc_hd__o211a_2
XFILLER_56_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout372_A _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _04952_ net660 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_3_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06816_ _03469_ _03470_ _03471_ _03472_ net762 net752 vssd1 vssd1 vccd1 vccd1 _03473_
+ sky130_fd_sc_hd__mux4_1
X_07796_ _04432_ _04442_ _04452_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__or3_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06192__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09535_ top0.CPU.control.funct3\[1\] _05081_ net125 vssd1 vssd1 vccd1 vccd1 _01104_
+ sky130_fd_sc_hd__mux2_1
X_06747_ _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__inv_2
XANTENNA__08469__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685__337 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__inv_2
X_09466_ net130 net134 _05051_ net597 net3417 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__o32a_1
X_06678_ top0.CPU.register.registers\[257\] top0.CPU.register.registers\[289\] top0.CPU.register.registers\[321\]
+ top0.CPU.register.registers\[353\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07692__A1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08417_ net160 net690 net391 net377 net2352 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a32o_1
XANTENNA__08484__A3 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ _05000_ _05001_ _05005_ _04949_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a31o_1
XANTENNA__07692__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ net721 net169 net402 net411 net2548 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a32o_1
X_10437__89 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__inv_2
X_10726__378 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__inv_2
XANTENNA__08236__A3 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06878__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08641__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ net504 net177 net672 net419 net2696 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a32o_1
X_10310_ _02359_ _05640_ _05639_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__o21ai_1
X_10241_ net14 net655 net594 top0.MMIO.WBData_i\[20\] vssd1 vssd1 vccd1 vccd1 _02287_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579__231 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__inv_2
X_11363__1015 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__inv_2
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__buf_2
X_10172_ _02992_ _03001_ _05577_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05853__S1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1129 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_4
Xfanout1115 net1132 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_4
Xfanout183 _04596_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_1
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
Xfanout172 _04611_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout161 net163 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
XANTENNA__06802__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09657__C1 _02532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05930__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08475__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06030__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ clknet_leaf_82_clk _02310_ net1109 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07683__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08227__A3 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10129__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11626_ net1318 _01265_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06869__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ net1249 _01196_ net1040 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08632__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold609 top0.CPU.register.registers\[221\] vssd1 vssd1 vccd1 vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08314__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ clknet_leaf_81_clk top0.display.next_state\[0\] net1111 vssd1 vssd1 vccd1
+ vccd1 top0.display.state\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__10145__A _02906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06097__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__A2 _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05844__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05980_ top0.CPU.register.registers\[901\] top0.CPU.register.registers\[933\] top0.CPU.register.registers\[965\]
+ top0.CPU.register.registers\[997\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02637_
+ sky130_fd_sc_hd__mux4_1
X_12109_ net1801 _01748_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07650_ net342 _04297_ _04298_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ top0.CPU.register.registers\[135\] top0.CPU.register.registers\[167\] top0.CPU.register.registers\[199\]
+ top0.CPU.register.registers\[231\] net927 net893 vssd1 vssd1 vccd1 vccd1 _03258_
+ sky130_fd_sc_hd__mux4_1
X_07581_ net488 _03894_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__or2_1
XANTENNA__08556__Y _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06532_ top0.CPU.register.registers\[146\] top0.CPU.register.registers\[178\] top0.CPU.register.registers\[210\]
+ top0.CPU.register.registers\[242\] net931 net897 vssd1 vssd1 vccd1 vccd1 _03189_
+ sky130_fd_sc_hd__mux4_1
X_09320_ _04966_ _04969_ _04970_ _04971_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_105_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09251_ _04106_ net232 net227 _02337_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__a31o_1
XFILLER_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06517__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07674__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06463_ top0.CPU.register.registers\[660\] top0.CPU.register.registers\[692\] top0.CPU.register.registers\[724\]
+ top0.CPU.register.registers\[756\] net918 net884 vssd1 vssd1 vccd1 vccd1 _03120_
+ sky130_fd_sc_hd__mux4_1
X_08202_ net209 net679 vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_138_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06882__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09415__A2 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08218__A3 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06394_ _03047_ _03048_ _03050_ _03049_ net870 net754 vssd1 vssd1 vccd1 vccd1 _03051_
+ sky130_fd_sc_hd__mux4_1
X_09182_ top0.CPU.register.registers\[33\] net564 net552 vssd1 vssd1 vccd1 vccd1 _04849_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_138_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout120_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ net2685 net177 net429 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
XANTENNA__08623__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05780__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout218_A _04603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08064_ net224 net693 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and2_1
X_07015_ _03670_ _03671_ net763 vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__mux2_1
XANTENNA__09179__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07348__B _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09563__B _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06679__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _04659_ net267 net259 net2732 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net719 net193 _04767_ net283 net3312 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__a32o_1
X_07917_ _04476_ _04557_ _04558_ _04559_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_95_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08154__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07848_ net591 _02946_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__nand2_1
XFILLER_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06260__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11246__898 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09518_ top0.MMIO.WBData_i\[23\] top0.MMIO.WBData_i\[19\] top0.MMIO.WBData_i\[1\]
+ _02358_ net137 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__a41o_1
X_07779_ _02578_ _03720_ _03877_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or3_1
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06708__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06267__X _02924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ top0.MMIO.WBData_i\[18\] net146 net135 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06012__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099__751 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__inv_2
X_12460_ net2152 _02099_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[953\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08614__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11411_ clknet_leaf_77_clk _01059_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12391_ net2083 _02030_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[884\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07098__X _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08090__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05979__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06079__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ net27 net657 net596 top0.MMIO.WBData_i\[3\] vssd1 vssd1 vccd1 vccd1 _02270_
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ net3426 net663 net602 _05615_ _05612_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a221o_1
XANTENNA__08393__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
X_10086_ _04967_ _05548_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__o21ai_1
Xhold6 top0.CPU.register.registers\[20\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06156__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08309__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__A0 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ clknet_leaf_66_clk _02293_ net1104 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ net1301 _01248_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06616__C1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09648__B top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ clknet_leaf_84_clk _02224_ net1107 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_10_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold417 top0.CPU.register.registers\[455\] vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold406 top0.CPU.register.registers\[381\] vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold439 top0.CPU.register.registers\[239\] vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 top0.CPU.register.registers\[164\] vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08908__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ net183 net676 net323 net287 net2461 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a32o_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout919 net941 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_2
Xfanout908 net910 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_4
XANTENNA__08384__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 top0.display.dataforOutput\[12\] vssd1 vssd1 vccd1 vccd1 net3328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07592__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08751_ net191 net624 net327 net296 net2521 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_77_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
Xhold1139 net37 vssd1 vssd1 vccd1 vccd1 net3361 sky130_fd_sc_hd__dlygate4sd3_1
X_05963_ top0.CPU.decoder.instruction\[11\] _02448_ _02535_ net774 net583 vssd1 vssd1
+ vccd1 vccd1 _02620_ sky130_fd_sc_hd__a221o_1
Xhold1128 top0.display.dataforOutput\[3\] vssd1 vssd1 vccd1 vccd1 net3350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 top0.CPU.register.registers\[260\] vssd1 vssd1 vccd1 vccd1 net3339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06490__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08682_ net182 net696 net323 net299 net2549 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_107_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09333__A1 _04292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ _03740_ _04141_ _04142_ net442 vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05894_ _02544_ _02550_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__nand2_1
X_10948__600 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__inv_2
XANTENNA__07912__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ net517 _04286_ _04287_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout168_A _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06242__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ net344 net441 _03810_ _03357_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__a22o_1
X_06515_ _03168_ _03171_ net754 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
X_09303_ net577 _04952_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11362__1014 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__inv_2
X_07495_ _02496_ _03193_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout335_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ _02337_ top0.CPU.intMemAddr\[10\] vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06446_ net866 _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1077_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09165_ net200 net673 _04846_ net249 net3236 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_32_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1185_A top0.CPU.intMem_out\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06377_ top0.CPU.register.registers\[414\] top0.CPU.register.registers\[446\] top0.CPU.register.registers\[478\]
+ top0.CPU.register.registers\[510\] net935 net903 vssd1 vssd1 vccd1 vccd1 _03034_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ net2830 net207 net432 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
X_10407__59 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__inv_2
XANTENNA_fanout502_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10797__449 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__inv_2
X_09096_ _04690_ net558 _04823_ net254 net3090 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__a32o_1
X_08047_ net504 net188 net706 net438 net2322 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a32o_1
Xhold940 top0.CPU.register.registers\[250\] vssd1 vssd1 vccd1 vccd1 net3162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 top0.CPU.register.registers\[527\] vssd1 vssd1 vccd1 vccd1 net3184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold951 net101 vssd1 vssd1 vccd1 vccd1 net3173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 top0.CPU.register.registers\[985\] vssd1 vssd1 vccd1 vccd1 net3195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold984 top0.CPU.register.registers\[261\] vssd1 vssd1 vccd1 vccd1 net3206 sky130_fd_sc_hd__dlygate4sd3_1
X_10541__193 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__inv_2
XFILLER_103_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout871_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 top0.CPU.register.registers\[667\] vssd1 vssd1 vccd1 vccd1 net3217 sky130_fd_sc_hd__dlygate4sd3_1
X_09998_ top0.CPU.internalMem.pcOut\[28\] _05486_ vssd1 vssd1 vccd1 vccd1 _05488_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_73_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07583__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ net176 net706 _04781_ net265 net3346 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_68_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
X_11960_ net1652 _01599_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11891_ net1583 _01530_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[384\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07541__B _03037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09088__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07350__A3 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A0 _04498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ net2204 _02151_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1005\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_100_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12443_ net2135 _02082_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[936\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08063__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07269__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12374_ net2066 _02013_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[867\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12566__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09484__A top0.MMIO.WBData_i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421__73 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__inv_2
XANTENNA__06901__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08366__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ net44 net121 net115 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a21o_1
XFILLER_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10138_ _05600_ _05601_ net600 vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_59_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
X_10069_ top0.display.delayctr\[7\] _05545_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__or2_2
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05951__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09079__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07341__A3 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05983__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08826__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ _03760_ _03927_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__or2_1
X_06300_ top0.CPU.register.registers\[155\] top0.CPU.register.registers\[187\] top0.CPU.register.registers\[219\]
+ top0.CPU.register.registers\[251\] net828 net791 vssd1 vssd1 vccd1 vccd1 _02957_
+ sky130_fd_sc_hd__mux4_1
X_06231_ _02871_ _02887_ net583 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux2_2
X_10484__136 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06162_ _02817_ _02818_ net784 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XANTENNA__08054__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10525__177 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__inv_2
Xhold214 top0.CPU.register.registers\[360\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 top0.CPU.register.registers\[304\] vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
X_06093_ net581 _02734_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__o21ai_4
Xhold225 top0.CPU.register.registers\[193\] vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 top0.CPU.register.registers\[972\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09394__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold269 top0.CPU.intMemAddr\[12\] vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ top0.CPU.internalMem.pcOut\[21\] _05394_ top0.CPU.internalMem.pcOut\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06160__S0 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 top0.CPU.register.registers\[967\] vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 top0.CPU.register.registers\[32\] vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12236__RESET_B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06060__A1_N _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 net712 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_4
XANTENNA__09003__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout738 net740 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_113_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ top0.CPU.internalMem.pcOut\[17\] _05352_ vssd1 vssd1 vccd1 vccd1 _05353_
+ sky130_fd_sc_hd__nand2_1
Xfanout727 _02349_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
Xfanout749 net755 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_4
Xfanout716 net723 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_2
X_09783_ _05272_ _05276_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a21oi_1
X_08803_ _04711_ net305 net285 net2967 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a22o_1
XFILLER_100_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09306__A1 _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _04676_ net308 net293 net2876 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__a22o_1
X_06995_ top0.CPU.register.registers\[410\] top0.CPU.register.registers\[442\] top0.CPU.register.registers\[474\]
+ top0.CPU.register.registers\[506\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03652_
+ sky130_fd_sc_hd__mux4_1
XFILLER_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05946_ top0.CPU.register.registers\[897\] top0.CPU.register.registers\[929\] top0.CPU.register.registers\[961\]
+ top0.CPU.register.registers\[993\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02603_
+ sky130_fd_sc_hd__mux4_1
X_05877_ _02532_ net579 top0.CPU.control.funct7\[6\] _02518_ vssd1 vssd1 vccd1 vccd1
+ _02534_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout452_A _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06215__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _04657_ net308 net297 net2735 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a22o_1
XFILLER_54_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07616_ _03759_ _04266_ _04267_ _03747_ _03841_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o221a_1
X_08596_ net3061 net330 net317 _04493_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ _02812_ _03222_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__nor2_1
XANTENNA__05974__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07096__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ _02925_ net523 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__xnor2_1
X_09217_ _04877_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__or2_1
X_06429_ net750 _03085_ net858 vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08045__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ top0.CPU.register.registers\[61\] _02396_ vssd1 vssd1 vccd1 vccd1 _04843_
+ sky130_fd_sc_hd__or2_1
X_09079_ net186 net619 _04819_ net257 net3284 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08596__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07376__X _04033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold781 top0.CPU.intMemAddr\[28\] vssd1 vssd1 vccd1 vccd1 net3003 sky130_fd_sc_hd__dlygate4sd3_1
X_12090_ net1782 _01729_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[583\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06721__A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 top0.CPU.register.registers\[150\] vssd1 vssd1 vccd1 vccd1 net2992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold792 top0.CPU.register.registers\[883\] vssd1 vssd1 vccd1 vccd1 net3014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08899__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261__913 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__inv_2
XANTENNA__06206__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ net1635 _01582_ net999 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[436\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11874_ net1566 _01513_ net1047 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07271__B _03092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05965__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08808__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302__954 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__inv_2
XANTENNA__08823__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06455__X _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06390__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ net2118 _02065_ net995 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[919\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12357_ net2049 _01996_ net1036 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06142__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12288_ net1980 _01927_ net1044 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06693__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361__1013 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__inv_2
XANTENNA__08339__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09000__A3 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05800_ _02446_ _02456_ net580 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_2
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06780_ _03435_ _03436_ net765 vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__mux2_1
X_10910__562 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__inv_2
X_05731_ net652 _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__nor2_4
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08511__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ net2863 net166 net373 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__mux2_1
XANTENNA__07181__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08381_ net169 net709 net402 net383 net2358 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a32o_1
X_07401_ net245 _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07332_ _03971_ _03985_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__nand3_2
X_11045__697 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__inv_2
XANTENNA__09389__A _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ _03918_ _03919_ net459 vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__mux2_1
X_06214_ net787 net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a21oi_2
X_07194_ net453 net518 _03747_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a21o_1
X_09002_ net157 net690 net267 net259 net2589 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__a32o_1
XANTENNA__09775__A1 top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06145_ top0.CPU.register.registers\[145\] top0.CPU.register.registers\[177\] top0.CPU.register.registers\[209\]
+ top0.CPU.register.registers\[241\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02802_
+ sky130_fd_sc_hd__mux4_1
X_06076_ _02619_ _02686_ _02731_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_57_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06684__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_2
X_09904_ _05399_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__nand2_1
Xfanout524 _03556_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _05294_ _05309_ _05320_ _05330_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__nand4_1
Xfanout557 net560 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07924__X _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 _03173_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07002__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 net548 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_4
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout579 _02422_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_2
XANTENNA__06761__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _05250_ _05260_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__nand2_1
XANTENNA__08750__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06978_ top0.CPU.register.registers\[283\] top0.CPU.register.registers\[315\] top0.CPU.register.registers\[347\]
+ top0.CPU.register.registers\[379\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03635_
+ sky130_fd_sc_hd__mux4_1
X_09697_ _04127_ net233 net228 net589 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__and4b_1
X_08717_ net186 net3203 net359 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout834_A top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07803__C _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05929_ net786 _02583_ net780 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__o21a_1
X_08648_ net186 net706 net318 net303 net2444 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a32o_1
XFILLER_42_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08502__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ net2839 net181 net336 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__mux2_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ net1282 _01229_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09299__A top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06372__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ net1903 _01850_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[704\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06722__Y _03379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ net1834 _01781_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[635\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06675__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10853__505 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__inv_2
X_12073_ net1765 _01712_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[566\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09762__A top0.CPU.control.funct7\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10128__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06427__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08741__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11926_ net1618 _01565_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[419\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ net1549 _01496_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[350\]
+ sky130_fd_sc_hd__dfrtp_1
X_11788_ net1480 _01427_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08317__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07465__C1 _03743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
X_12409_ net2101 _02048_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06666__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ net723 net513 net190 net549 net2391 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a32o_1
XFILLER_114_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596__248 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__inv_2
XANTENNA__08980__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10119__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ net524 _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__or2_1
XANTENNA__06991__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07881_ net3219 net546 net492 _04529_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
X_10637__289 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__inv_2
XANTENNA__07904__B _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09620_ _02343_ _05006_ net550 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o21a_1
X_06832_ _02619_ _02686_ _02718_ _02730_ net540 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_52_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08732__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06763_ top0.CPU.register.registers\[271\] top0.CPU.register.registers\[303\] top0.CPU.register.registers\[335\]
+ top0.CPU.register.registers\[367\] net936 net902 vssd1 vssd1 vccd1 vccd1 _03420_
+ sky130_fd_sc_hd__mux4_1
X_09551_ top0.CPU.control.funct7\[4\] _05086_ net125 vssd1 vssd1 vccd1 vccd1 _01120_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07940__B1 _02734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05714_ top0.CPU.Op\[6\] top0.CPU.Op\[3\] vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__or2_1
X_08502_ _04702_ net388 net365 net3073 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__a22o_1
X_09482_ top0.MMIO.WBData_i\[27\] net137 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__or2_1
X_06694_ _03349_ _03350_ net764 vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__mux2_1
X_08433_ net2916 net223 net374 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
XANTENNA__08248__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _04646_ net395 net382 net2578 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a22o_1
XANTENNA__08799__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _03727_ _03926_ _03946_ net484 vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__o22a_1
XANTENNA__07456__C1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06354__S0 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ net3063 net207 net414 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__mux2_1
X_07246_ _03760_ _03895_ _03896_ _03851_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o221a_1
XANTENNA__06106__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07177_ net485 _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__nor2_1
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06657__S1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06128_ top0.CPU.register.registers\[270\] top0.CPU.register.registers\[302\] top0.CPU.register.registers\[334\]
+ top0.CPU.register.registers\[366\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02785_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout784_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06059_ top0.CPU.control.funct7\[3\] _02518_ _02715_ net579 vssd1 vssd1 vccd1 vccd1
+ _02716_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__08971__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout332 _04735_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
Xfanout321 net326 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_4
Xfanout310 net313 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_2
XANTENNA__08184__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout951_A top0.CPU.decoder.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__A4 _02355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout343 _03716_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
Xfanout354 _04752_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_8
Xfanout365 _04728_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_8
Xfanout376 _04726_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_4
X_09818_ _05300_ _05321_ _05308_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__o21a_1
Xfanout398 net399 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout387 net393 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_2
X_09749_ _04044_ net234 net229 net631 vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a31o_1
XANTENNA__09279__A3 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11711_ net1403 _01350_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[204\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10294__A1 _02446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12691_ clknet_leaf_93_clk _02326_ net1082 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XFILLER_42_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11360__1012 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__inv_2
X_11642_ net1334 _01281_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[135\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08137__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06446__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07998__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09987__B2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11573_ net1265 _01212_ net970 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06896__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ net1817 _01764_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[618\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06648__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12056_ net1748 _01695_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[549\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output44_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11308__960 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__inv_2
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10150__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ net1601 _01548_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[402\]
+ sky130_fd_sc_hd__dfrtp_1
X_10981__633 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__inv_2
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_44_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09978__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ net347 _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__or3_1
XANTENNA__06887__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08080_ net204 net700 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__and2_1
X_07031_ top0.CPU.register.registers\[543\] top0.CPU.register.registers\[575\] top0.CPU.register.registers\[607\]
+ top0.CPU.register.registers\[639\] net851 net817 vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__mux4_1
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08982_ net200 net694 _04791_ net260 net3310 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__a32o_1
XANTENNA__08953__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07933_ _04331_ net231 net226 vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__and3_1
X_07864_ top0.CPU.intMem_out\[25\] net627 _04514_ net642 vssd1 vssd1 vccd1 vccd1 _04515_
+ sky130_fd_sc_hd__a211o_1
X_10382__34 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__inv_2
X_06815_ top0.CPU.register.registers\[525\] top0.CPU.register.registers\[557\] top0.CPU.register.registers\[589\]
+ top0.CPU.register.registers\[621\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03472_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08181__A3 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ top0.display.dataforOutput\[3\] net604 net658 top0.display.dataforOutput\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ net342 _04443_ _04444_ _04451_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout365_A _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ top0.CPU.control.funct3\[0\] _05075_ net126 vssd1 vssd1 vccd1 vccd1 _01103_
+ sky130_fd_sc_hd__mux2_1
X_06746_ net745 _03402_ _03395_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__a21oi_4
X_09465_ top0.MMIO.WBData_i\[26\] net145 net135 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__o21a_1
XANTENNA__09130__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060__712 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__inv_2
XANTENNA_fanout532_A _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06677_ top0.CPU.register.registers\[385\] top0.CPU.register.registers\[417\] top0.CPU.register.registers\[449\]
+ top0.CPU.register.registers\[481\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03334_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08416_ net166 net693 net392 net377 net2660 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a32o_1
X_09396_ _02408_ _05000_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__or2_1
XANTENNA__07692__A2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11101__753 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__inv_2
X_08347_ net715 net173 net390 net409 net2497 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06878__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06101__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__C net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ net506 net220 net672 net419 net2387 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a32o_1
X_07229_ _03853_ _03855_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07809__B _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ net12 net656 net595 top0.MMIO.WBData_i\[19\] vssd1 vssd1 vccd1 vccd1 _02286_
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07097__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net3414 net664 net661 _05625_ _05628_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a221o_1
XANTENNA__07825__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1127 net1129 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout140 _05013_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1116 net1118 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout151 _04482_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
Xfanout173 _04611_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_2
Xfanout184 _04596_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
Xfanout195 _04582_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08172__A3 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06802__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965__617 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__inv_2
XFILLER_55_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09121__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ clknet_leaf_81_clk _02309_ net1109 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ net1317 _01264_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06869__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07435__A2 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ net1248 _01195_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10859__511 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__inv_2
X_11487_ clknet_leaf_83_clk _01129_ net1111 vssd1 vssd1 vccd1 vccd1 top0.display.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08396__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08935__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12108_ net1800 _01747_ net968 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[601\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05954__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ net1731 _01678_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[532\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09950__A top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06600_ top0.CPU.register.registers\[391\] top0.CPU.register.registers\[423\] top0.CPU.register.registers\[455\]
+ top0.CPU.register.registers\[487\] net915 net881 vssd1 vssd1 vccd1 vccd1 _03257_
+ sky130_fd_sc_hd__mux4_1
X_07580_ _04051_ _04060_ net478 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
X_06531_ _03186_ _03187_ net871 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09250_ top0.CPU.internalMem.pcOut\[7\] top0.CPU.addrControl _04910_ _04911_ vssd1
+ vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a22o_1
XANTENNA__06557__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06462_ top0.CPU.register.registers\[788\] top0.CPU.register.registers\[820\] top0.CPU.register.registers\[852\]
+ top0.CPU.register.registers\[884\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03119_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07725__A1_N net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08201_ net3127 net421 _04693_ net494 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
XANTENNA__06309__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09181_ net163 net669 net270 net247 net2533 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__a32o_1
X_06393_ top0.CPU.register.registers\[29\] top0.CPU.register.registers\[61\] top0.CPU.register.registers\[93\]
+ top0.CPU.register.registers\[125\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03050_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08132_ net3126 net219 net430 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XANTENNA__08623__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05780__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ net2775 net434 _04654_ net514 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07014_ top0.CPU.register.registers\[543\] top0.CPU.register.registers\[575\] top0.CPU.register.registers\[607\]
+ top0.CPU.register.registers\[639\] net937 net902 vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout113_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__B _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07348__C _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06025__S net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05864__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _04658_ net267 net259 net2799 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__a22o_1
XFILLER_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07916_ _02386_ _02793_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nor2_1
XANTENNA__07364__B _03540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10652__304 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__inv_2
X_08896_ top0.CPU.register.registers\[237\] net572 net558 vssd1 vssd1 vccd1 vccd1
+ _04767_ sky130_fd_sc_hd__o21a_1
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _04378_ net231 net226 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_67_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06796__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ _04286_ _04287_ net453 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09517_ _05091_ _05095_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__and3_1
X_06729_ _03250_ _03261_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__or2_1
XANTENNA__09103__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__S0 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ net131 net133 _05042_ net598 net3360 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__o32a_1
X_09379_ net2624 _04518_ net606 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08614__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ net2082 _02029_ net1129 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[883\]
+ sky130_fd_sc_hd__dfrtp_1
X_11410_ clknet_leaf_87_clk _01058_ net1090 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08923__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05979__A2 _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__S0 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ net24 net656 net595 top0.MMIO.WBData_i\[2\] vssd1 vssd1 vccd1 vccd1 _02269_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08917__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ _05613_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08003__X _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold7 top0.CPU.register.registers\[18\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ top0.display.delayctr\[11\] _05557_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__nand2_1
XANTENNA__09770__A top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07353__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08550__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07290__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07105__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__A2 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06313__C1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12657_ clknet_leaf_66_clk _02292_ net1101 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11608_ net1300 _01247_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06193__X _02850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12588_ clknet_leaf_84_clk _02223_ net1107 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06634__A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 top0.CPU.register.registers\[338\] vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 top0.CPU.register.registers\[349\] vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
X_11539_ net1231 _01178_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08081__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold429 top0.CPU.register.registers\[906\] vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10176__B1 _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_4
XANTENNA__08384__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1118 top0.CPU.register.registers\[74\] vssd1 vssd1 vccd1 vccd1 net3340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1107 top0.CPU.register.registers\[69\] vssd1 vssd1 vccd1 vccd1 net3329 sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ net193 net620 _04748_ net295 net3318 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__a32o_1
Xhold1129 _01133_ vssd1 vssd1 vccd1 vccd1 net3351 sky130_fd_sc_hd__dlygate4sd3_1
X_05962_ net476 net471 net462 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_107_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ net186 net694 net318 net299 net2286 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a32o_1
XFILLER_66_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07701_ _02888_ _03112_ net446 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__or3_1
X_05893_ net772 _02549_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__or2_2
XANTENNA__08541__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07912__B _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07632_ _03758_ _04286_ _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__and3_1
XANTENNA__06778__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09302_ top0.display.state\[1\] top0.display.state\[2\] top0.display.state\[0\] vssd1
+ vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__or3b_2
X_07563_ _03738_ _04171_ _04170_ net339 vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__o2bb2a_1
X_06514_ _03169_ _03170_ net766 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07494_ _04149_ _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nor2_1
XFILLER_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09233_ net769 _04593_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__and2_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06445_ _03100_ _03101_ net764 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout328_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09164_ top0.CPU.register.registers\[48\] net570 net558 vssd1 vssd1 vccd1 vccd1 _04846_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06376_ top0.CPU.register.registers\[30\] top0.CPU.register.registers\[62\] top0.CPU.register.registers\[94\]
+ top0.CPU.register.registers\[126\] net937 net901 vssd1 vssd1 vccd1 vccd1 _03033_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06544__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08115_ net3087 net208 net429 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
X_09095_ top0.CPU.register.registers\[94\] net572 vssd1 vssd1 vccd1 vccd1 _04823_
+ sky130_fd_sc_hd__or2_1
X_11172__824 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__inv_2
X_08046_ net513 net190 net710 net440 net2480 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a32o_1
Xhold930 net95 vssd1 vssd1 vccd1 vccd1 net3152 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold941 top0.CPU.register.registers\[777\] vssd1 vssd1 vccd1 vccd1 net3163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 top0.CPU.register.registers\[188\] vssd1 vssd1 vccd1 vccd1 net3174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 top0.CPU.register.registers\[571\] vssd1 vssd1 vccd1 vccd1 net3185 sky130_fd_sc_hd__dlygate4sd3_1
X_11213__865 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__inv_2
Xhold974 top0.CPU.register.registers\[393\] vssd1 vssd1 vccd1 vccd1 net3196 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08375__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 top0.CPU.register.registers\[892\] vssd1 vssd1 vccd1 vccd1 net3207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold996 top0.CPU.register.registers\[49\] vssd1 vssd1 vccd1 vccd1 net3218 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout864_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ top0.CPU.internalMem.pcOut\[28\] _05486_ vssd1 vssd1 vccd1 vccd1 _05487_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_73_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07583__A1 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ top0.CPU.register.registers\[199\] net570 net557 vssd1 vssd1 vccd1 vccd1
+ _04781_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09590__A _02596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ net2960 net282 net267 _04529_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__a22o_1
XFILLER_84_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08532__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__A1 _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ net1582 _01529_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ net2203 _02150_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1004\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ net2134 _02081_ net981 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[935\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780__432 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__inv_2
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08063__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06173__B _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07269__B net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12373_ net2065 _02012_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[866\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08239__C_N net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09765__A top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07837__X _04492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821__473 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__inv_2
XFILLER_109_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ net2800 net123 net116 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a21o_1
XFILLER_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ top0.display.delayctr\[22\] _05596_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nand2_1
XFILLER_0_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08771__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ net3419 net664 net602 _05547_ _05147_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08523__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07224__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09005__A _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05983__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08826__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09659__B _05169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06230_ net742 _02886_ _02879_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__a21oi_4
XANTENNA__06932__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06364__A _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156__808 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09251__A1 _04106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06161_ top0.CPU.register.registers\[912\] top0.CPU.register.registers\[944\] top0.CPU.register.registers\[976\]
+ top0.CPU.register.registers\[1008\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02818_
+ sky130_fd_sc_hd__mux4_1
Xhold204 top0.CPU.register.registers\[594\] vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
X_06092_ net581 _02748_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__nand2_1
Xhold215 top0.CPU.register.registers\[715\] vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 top0.CPU.register.registers\[738\] vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07262__A0 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09394__B top0.CPU.control.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 top0.CPU.register.registers\[361\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 top0.CPU.register.registers\[461\] vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ top0.CPU.internalMem.pcOut\[22\] top0.CPU.internalMem.pcOut\[21\] _05394_
+ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__and3_1
XANTENNA__06160__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold259 top0.CPU.register.registers\[483\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09003__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10149__B1 _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout739 net740 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_113_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout728 net730 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_4
X_09851_ net587 _04557_ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a21o_1
XANTENNA__07565__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 net723 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_4
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09782_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__and2_1
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06994_ _03649_ _03650_ net756 vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__mux2_1
X_08802_ _04710_ net308 net285 net2824 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a22o_1
XANTENNA__08762__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09306__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ _04675_ net311 net293 net2678 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a22o_1
X_05945_ top0.CPU.register.registers\[769\] top0.CPU.register.registers\[801\] top0.CPU.register.registers\[833\]
+ top0.CPU.register.registers\[865\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02602_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout180_A _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08514__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05876_ top0.CPU.control.funct7\[6\] _02518_ _02532_ net579 vssd1 vssd1 vccd1 vccd1
+ _02533_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08664_ _04656_ net311 net297 net2936 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a22o_1
X_08595_ net3257 net331 net324 _04488_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__a22o_1
XANTENNA__05879__A1 top0.CPU.decoder.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05879__B2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout445_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07615_ _03320_ _03360_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10764__416 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__inv_2
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07546_ _04130_ _04197_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__a21o_1
XANTENNA__05974__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06973__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ _04475_ _04494_ _04506_ _04512_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__or4_1
X_07477_ _04132_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08192__C net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805__457 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__inv_2
X_06428_ _03083_ _03084_ net869 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
X_09147_ _04707_ net279 net250 net2460 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__a22o_1
X_06359_ top0.CPU.register.registers\[414\] top0.CPU.register.registers\[446\] top0.CPU.register.registers\[478\]
+ top0.CPU.register.registers\[510\] net850 net818 vssd1 vssd1 vccd1 vccd1 _03016_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07089__B net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ top0.CPU.register.registers\[107\] net570 net557 vssd1 vssd1 vccd1 vccd1
+ _04819_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_75_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08029_ net3260 net437 _04645_ net492 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
Xhold760 top0.CPU.register.registers\[499\] vssd1 vssd1 vccd1 vccd1 net2982 sky130_fd_sc_hd__dlygate4sd3_1
X_10658__310 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__inv_2
Xhold782 top0.CPU.register.registers\[567\] vssd1 vssd1 vccd1 vccd1 net3004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 top0.CPU.register.registers\[771\] vssd1 vssd1 vccd1 vccd1 net2993 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 net98 vssd1 vssd1 vccd1 vccd1 net3015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08753__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__A1 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ net1634 _01581_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[435\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07044__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ net1565 _01512_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[366\]
+ sky130_fd_sc_hd__dfrtp_1
X_11341__993 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__inv_2
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05965__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06390__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12425_ net2117 _02064_ net1074 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[918\]
+ sky130_fd_sc_hd__dfrtp_1
X_12356_ net2048 _01995_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08992__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06142__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12287_ net1979 _01926_ net1094 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[780\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06123__S net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08744__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451__103 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__inv_2
X_05730_ _02375_ _02376_ _02380_ net640 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__and4_1
XFILLER_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__A3 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06793__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08380_ net173 net703 net391 net381 net2524 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a32o_1
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ _03906_ _03926_ _04056_ net484 vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_34_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07331_ _02533_ _03504_ net444 _03986_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ net522 net537 net467 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__mux2_1
X_06213_ _02852_ _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_1
X_09001_ net160 net691 net270 net259 net2303 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__a32o_1
X_07193_ net490 _03758_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nand2_2
XANTENNA__08027__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06144_ net736 _02800_ net772 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08983__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07637__B _04127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06075_ _02619_ _02686_ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_57_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_2
X_09903_ net586 _04535_ _05398_ top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1
+ vccd1 _05400_ sky130_fd_sc_hd__a211o_1
XANTENNA__05892__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout503 net516 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_9_0_clk_X clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_4
X_09834_ net652 _05333_ _05335_ _05336_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__o31a_1
XFILLER_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout525 _03540_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08735__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 _03112_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284__936 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__inv_2
Xfanout569 _02388_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold1210_A top0.CPU.intMem_out\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ top0.CPU.internalMem.pcOut\[10\] _05271_ vssd1 vssd1 vccd1 vccd1 _05273_
+ sky130_fd_sc_hd__xor2_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06977_ top0.CPU.register.registers\[411\] top0.CPU.register.registers\[443\] top0.CPU.register.registers\[475\]
+ top0.CPU.register.registers\[507\] net911 net879 vssd1 vssd1 vccd1 vccd1 _03634_
+ sky130_fd_sc_hd__mux4_1
XFILLER_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08716_ _04586_ net3314 net360 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__mux2_1
X_09696_ top0.CPU.internalMem.pcOut\[4\] net650 _05209_ vssd1 vssd1 vccd1 vccd1 _02181_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07803__D net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05928_ net733 _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__or2_1
X_08647_ net191 net710 net327 net304 net2446 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a32o_1
XANTENNA__09160__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325__977 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__inv_2
X_05859_ _02338_ net626 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ net2835 net184 net336 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07529_ _02750_ _03483_ _04185_ _02769_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__o22a_1
X_11178__830 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__inv_2
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06372__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ net1902 _01849_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[703\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08931__B net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219__871 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__inv_2
XANTENNA__08423__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10892__544 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__inv_2
X_10388__40 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__inv_2
XANTENNA__07547__B _03222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10254__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net1833 _01780_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[634\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold590 top0.CPU.register.registers\[330\] vssd1 vssd1 vccd1 vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05883__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ net1764 _01711_ net1077 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[565\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07529__B2 _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10933__585 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__inv_2
XFILLER_92_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_88_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11925_ net1617 _01564_ net977 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ net1548 _01495_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[349\]
+ sky130_fd_sc_hd__dfrtp_1
X_11787_ net1479 _01426_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06268__A1 _02924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12408_ net2100 _02047_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[901\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XANTENNA__08965__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ net2031 _01978_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05874__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06900_ _02716_ _03522_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__xnor2_1
X_07880_ net716 net152 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__and2_1
X_06831_ _03426_ _03445_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__or3_1
XFILLER_56_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_52_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11012__664 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__inv_2
X_06762_ net865 _03414_ _03417_ _03418_ net861 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__o221a_1
X_09550_ top0.CPU.control.funct7\[3\] _05079_ net126 vssd1 vssd1 vccd1 vccd1 _01119_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07940__B2 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09481_ _02336_ net148 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__nand2_1
X_08501_ _04556_ net684 net406 net367 net2426 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a32o_1
X_05713_ top0.CPU.Op\[0\] top0.CPU.Op\[1\] vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__nand2_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06051__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08496__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06693_ top0.CPU.register.registers\[0\] top0.CPU.register.registers\[32\] top0.CPU.register.registers\[64\]
+ top0.CPU.register.registers\[96\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__mux4_1
X_08432_ net3070 net204 net374 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__mux2_1
XANTENNA__06027__A1_N top0.CPU.control.funct7\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout143_A _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08248__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ _04645_ net387 net381 net2927 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
X_07314_ _03505_ _03520_ _03969_ _03970_ net344 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a311o_1
X_08294_ net3194 net208 net413 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
X_07245_ net477 _03892_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a21o_1
XFILLER_118_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout310_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06106__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876__528 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__inv_2
X_07176_ _03789_ _03831_ net347 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a21o_1
XFILLER_117_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06127_ top0.CPU.register.registers\[398\] top0.CPU.register.registers\[430\] top0.CPU.register.registers\[462\]
+ top0.CPU.register.registers\[494\] net836 net800 vssd1 vssd1 vccd1 vccd1 _02784_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08956__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06058_ net743 _02714_ _02707_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a21oi_4
X_10620__272 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__inv_2
Xfanout300 _04741_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
Xfanout322 net326 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout311 net313 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_2
X_10917__569 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__inv_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_8
Xfanout344 _03715_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_4
Xfanout333 _04733_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_6
Xfanout366 _04728_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06698__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ top0.CPU.internalMem.pcOut\[12\] _05293_ _05307_ vssd1 vssd1 vccd1 vccd1
+ _05321_ sky130_fd_sc_hd__a21bo_1
XFILLER_101_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout377 net378 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_4
XANTENNA__06195__A0 _02850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout388 net393 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_4
X_09748_ top0.CPU.internalMem.pcOut\[8\] net650 _05257_ vssd1 vssd1 vccd1 vccd1 _02185_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA__08198__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06290__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09133__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ top0.CPU.internalMem.pcOut\[3\] net768 vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nand2_1
XANTENNA__09684__B2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__A1 top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ net1402 _01349_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10294__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ clknet_leaf_92_clk _02325_ net1082 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
X_11641_ net1333 _01280_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ net1264 _01211_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[65\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08947__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ net1816 _01763_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ net1747 _01694_ net974 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05806__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08175__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06281__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09124__B1 _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08478__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06033__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ net1600 _01547_ net988 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[401\]
+ sky130_fd_sc_hd__dfrtp_1
X_11839_ net1531 _01478_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09300__X _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563__215 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__inv_2
XANTENNA__08650__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07030_ top0.CPU.register.registers\[671\] top0.CPU.register.registers\[703\] top0.CPU.register.registers\[735\]
+ top0.CPU.register.registers\[767\] net852 net817 vssd1 vssd1 vccd1 vccd1 _03687_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08938__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604__256 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08981_ top0.CPU.register.registers\[176\] net571 net560 vssd1 vssd1 vccd1 vccd1
+ _04791_ sky130_fd_sc_hd__o21a_1
XFILLER_130_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07932_ net721 net510 net196 net547 net2420 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a32o_1
XFILLER_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07863_ net561 _04512_ _04513_ net625 vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o211a_1
XANTENNA__08166__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06814_ top0.CPU.register.registers\[653\] top0.CPU.register.registers\[685\] top0.CPU.register.registers\[717\]
+ top0.CPU.register.registers\[749\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03471_
+ sky130_fd_sc_hd__mux4_1
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07913__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ top0.display.dataforOutput\[2\] net604 net658 net3350 _05139_ vssd1 vssd1
+ vccd1 vccd1 _01133_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06272__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ top0.CPU.decoder.instruction\[11\] _05077_ net125 vssd1 vssd1 vccd1 vccd1
+ _01102_ sky130_fd_sc_hd__mux2_1
XANTENNA__09115__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07794_ _03774_ _03882_ _04162_ net441 _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o221ai_2
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06745_ _03398_ _03401_ net862 vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout358_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08469__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ net131 net133 _05050_ net597 net3442 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__o32a_1
XANTENNA__09130__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06676_ _03331_ _03332_ net756 vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__mux2_1
X_09395_ net550 _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_65_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ net215 net691 net391 net378 net2356 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a32o_1
XANTENNA__07141__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_A _03540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ net714 net175 net390 net410 net2499 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140__792 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ net511 net181 net674 net420 net2600 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a32o_1
XANTENNA__08641__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07228_ _03849_ _03863_ _03882_ _03720_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__o221a_1
XFILLER_4_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__C net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ _03809_ _03815_ net348 vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__mux2_1
XANTENNA__08929__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358__10 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__inv_2
X_10170_ _05626_ _05627_ net600 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08701__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07825__B _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_2
Xfanout1106 net1132 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_2
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_2
Xfanout130 net132 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout174 _04611_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_1
Xfanout141 _04956_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout163 _04626_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout152 _04528_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
Xfanout196 net198 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
Xfanout185 _04596_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06263__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__B1 _02571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__A1 _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06015__S0 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_12673_ clknet_leaf_82_clk _02308_ net1108 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XFILLER_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11624_ net1316 _01263_ net1068 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08093__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11555_ net1247 _01194_ net1017 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08632__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11486_ clknet_leaf_81_clk _01128_ net1111 vssd1 vssd1 vccd1 vccd1 top0.display.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10898__550 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__inv_2
XFILLER_109_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10939__591 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__inv_2
X_10299_ _02942_ net551 net144 vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__o21ai_1
X_12107_ net1799 _01746_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[600\]
+ sky130_fd_sc_hd__dfrtp_1
X_12038_ net1730 _01677_ net1128 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[531\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08148__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06254__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__A _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083__735 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__inv_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06530_ top0.CPU.register.registers\[402\] top0.CPU.register.registers\[434\] top0.CPU.register.registers\[466\]
+ top0.CPU.register.registers\[498\] net931 net897 vssd1 vssd1 vccd1 vccd1 _03187_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06006__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06461_ top0.CPU.register.registers\[916\] top0.CPU.register.registers\[948\] top0.CPU.register.registers\[980\]
+ top0.CPU.register.registers\[1012\] net918 net884 vssd1 vssd1 vccd1 vccd1 _03118_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06557__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124__776 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__inv_2
XANTENNA_max_cap578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08200_ net210 net682 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__and2_1
XANTENNA__06882__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06309__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ net165 net669 net272 net247 net2283 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__a32o_1
X_06392_ top0.CPU.register.registers\[157\] top0.CPU.register.registers\[189\] top0.CPU.register.registers\[221\]
+ top0.CPU.register.registers\[253\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03049_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08131_ net2754 net181 net430 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
XANTENNA__07831__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ net212 net695 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__and2_1
XANTENNA__07198__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07013_ top0.CPU.register.registers\[671\] top0.CPU.register.registers\[703\] top0.CPU.register.registers\[735\]
+ top0.CPU.register.registers\[767\] net937 net902 vssd1 vssd1 vccd1 vccd1 _03670_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442__94 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__inv_2
XANTENNA__09179__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11018__670 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__inv_2
XFILLER_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ _04657_ net274 net259 net2858 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__a22o_1
X_07915_ top0.CPU.intMem_out\[17\] net628 net643 vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a21o_1
XANTENNA__08139__A1 _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691__343 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__inv_2
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08895_ net2908 _04753_ net274 _04577_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__a22o_1
XANTENNA__07898__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ net3009 net546 net498 _04499_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06245__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06796__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732__384 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__inv_2
XANTENNA_fanout642_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _03242_ _03941_ _03572_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_67_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09516_ _05057_ _05058_ _05085_ _05087_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__and4_1
XFILLER_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06728_ _03250_ _03261_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__nor2_1
X_09447_ top0.MMIO.WBData_i\[17\] _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and2_1
XFILLER_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06277__A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06659_ _03312_ _03315_ net862 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ net2989 _04524_ net608 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__mux2_1
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06564__X _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ net3057 net410 net395 _04523_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08090__A3 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__S1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ net13 net656 net595 top0.MMIO.WBData_i\[1\] vssd1 vssd1 vccd1 vccd1 _02268_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09527__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07555__B _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ top0.display.delayctr\[24\] _05604_ top0.display.delayctr\[25\] vssd1 vssd1
+ vccd1 vccd1 _05614_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11535__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10084_ net3403 net665 net603 _05559_ _05159_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold8 top0.CPU.register.registers\[21\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
X_11067__719 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07290__B _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08302__A1 _04561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12656_ clknet_leaf_71_clk _02291_ net1121 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_12587_ clknet_leaf_84_clk _02222_ net1107 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11607_ net1299 _01246_ net970 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06616__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08605__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11538_ net1230 _01177_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold408 top0.CPU.register.registers\[701\] vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 top0.CPU.register.registers\[47\] vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ clknet_leaf_60_clk _01117_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct7\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09945__B top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675__327 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__inv_2
XFILLER_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold1108 top0.display.dataforOutput\[8\] vssd1 vssd1 vccd1 vccd1 net3330 sky130_fd_sc_hd__dlygate4sd3_1
X_05961_ net477 net471 net463 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__and3_1
Xhold1119 net88 vssd1 vssd1 vccd1 vccd1 net3341 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ _04103_ _04356_ net452 vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07329__C1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ net191 net699 net327 net300 net2530 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a32o_1
X_05892_ _02545_ _02546_ _02548_ _02547_ net782 net735 vssd1 vssd1 vccd1 vccd1 _02549_
+ sky130_fd_sc_hd__mux4_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06227__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10716__368 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06778__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ net485 _04027_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XANTENNA__06809__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07562_ _02578_ _03906_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__or2_1
XANTENNA__08864__X _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06513_ top0.CPU.register.registers\[19\] top0.CPU.register.registers\[51\] top0.CPU.register.registers\[83\]
+ top0.CPU.register.registers\[115\] net940 net906 vssd1 vssd1 vccd1 vccd1 _03170_
+ sky130_fd_sc_hd__mux4_1
X_09301_ top0.display.state\[1\] top0.display.state\[2\] top0.display.state\[0\] vssd1
+ vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__nor3b_1
X_10569__221 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__inv_2
XFILLER_34_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07493_ _02831_ net533 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__xor2_1
X_09232_ top0.CPU.internalMem.pcOut\[10\] net609 vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__or2_1
X_06444_ top0.CPU.register.registers\[534\] top0.CPU.register.registers\[566\] top0.CPU.register.registers\[598\]
+ top0.CPU.register.registers\[630\] net922 net889 vssd1 vssd1 vccd1 vccd1 _03101_
+ sky130_fd_sc_hd__mux4_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06375_ top0.CPU.register.registers\[158\] top0.CPU.register.registers\[190\] top0.CPU.register.registers\[222\]
+ top0.CPU.register.registers\[254\] net935 net903 vssd1 vssd1 vccd1 vccd1 _03032_
+ sky130_fd_sc_hd__mux4_1
X_09163_ _04718_ net552 _04845_ net247 net3218 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__a32o_1
XANTENNA__08057__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_A _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08114_ net3055 _04510_ net429 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
X_09094_ net151 net688 net280 net254 net2588 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a32o_1
Xhold920 top0.CPU.register.registers\[755\] vssd1 vssd1 vccd1 vccd1 net3142 sky130_fd_sc_hd__dlygate4sd3_1
X_08045_ net511 net194 net709 net438 net2380 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a32o_1
Xhold931 net84 vssd1 vssd1 vccd1 vccd1 net3153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 top0.CPU.register.registers\[265\] vssd1 vssd1 vccd1 vccd1 net3175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 top0.CPU.register.registers\[1022\] vssd1 vssd1 vccd1 vccd1 net3164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 top0.CPU.register.registers\[391\] vssd1 vssd1 vccd1 vccd1 net3186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold986 top0.CPU.register.registers\[243\] vssd1 vssd1 vccd1 vccd1 net3208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold975 top0.CPU.register.registers\[540\] vssd1 vssd1 vccd1 vccd1 net3197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 top0.CPU.register.registers\[1015\] vssd1 vssd1 vccd1 vccd1 net3219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ net585 _04494_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_73_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07806__D net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net218 net706 net277 net265 net2430 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__a32o_1
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ net2972 net284 net274 _04523_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__a22o_1
X_07829_ net563 _04483_ _04484_ net626 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__o211a_1
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09088__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__Q top0.CPU.intMem_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ net2202 _02149_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1003\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08426__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ net2133 _02080_ net1012 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[934\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09796__B1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11787__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ net2064 _02011_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[865\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__A0 top0.CPU.control.funct7\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ net2985 net117 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10136_ top0.display.delayctr\[22\] _05596_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__or2_1
X_10067_ _05545_ _05546_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__nand2_1
XANTENNA__06209__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12575__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__A1_N net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09005__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09079__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08826__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06932__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ clknet_leaf_71_clk _02274_ net1119 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11195__847 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__inv_2
XANTENNA__06364__B _03020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06160_ top0.CPU.register.registers\[784\] top0.CPU.register.registers\[816\] top0.CPU.register.registers\[848\]
+ top0.CPU.register.registers\[880\] net844 net809 vssd1 vssd1 vccd1 vccd1 _02817_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08054__A3 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold205 top0.CPU.register.registers\[106\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
X_06091_ net773 _02739_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a21oi_4
Xhold216 top0.CPU.register.registers\[232\] vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06696__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07262__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__A0 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 top0.CPU.register.registers\[62\] vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 top0.CPU.register.registers\[585\] vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 top0.CPU.intMemAddr\[3\] vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_11236__888 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__inv_2
X_10412__64 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__inv_2
XFILLER_113_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__C _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06448__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout729 net730 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
Xfanout718 net722 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_4
Xfanout707 net711 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_4
X_09850_ net587 _02793_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__nor2_1
X_09781_ top0.CPU.internalMem.pcOut\[11\] _05284_ _05286_ vssd1 vssd1 vccd1 vccd1
+ _05288_ sky130_fd_sc_hd__nand3_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08801_ _04709_ net311 net285 net2766 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a22o_1
X_06993_ top0.CPU.register.registers\[26\] top0.CPU.register.registers\[58\] top0.CPU.register.registers\[90\]
+ top0.CPU.register.registers\[122\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03650_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06222__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11089__741 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__inv_2
X_08732_ _04674_ net317 net294 net2628 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a22o_1
X_05944_ _02599_ _02600_ net724 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
XANTENNA__07317__A2 _03504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08663_ _04655_ net317 net298 net2825 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a22o_1
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout173_A _04611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05875_ net743 _02531_ _02522_ _02526_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__o2bb2a_2
X_08594_ net2938 net332 _04738_ net722 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a22o_1
XANTENNA__06620__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07614_ net441 _04168_ _04268_ net245 vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_37_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08817__A2 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07545_ _03704_ _04198_ _04201_ _04128_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__o211ai_1
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_127_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout438_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_clk_X clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07476_ _02944_ net520 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__xnor2_1
XANTENNA_hold1190_A top0.CPU.intMem_out\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09215_ _04483_ _04489_ _04500_ _04518_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__or4_1
X_06427_ top0.CPU.register.registers\[919\] top0.CPU.register.registers\[951\] top0.CPU.register.registers\[983\]
+ top0.CPU.register.registers\[1015\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03084_
+ sky130_fd_sc_hd__mux4_1
X_10844__496 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__inv_2
X_09146_ net150 net675 net280 net250 net2528 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__a32o_1
X_06358_ top0.CPU.register.registers\[286\] top0.CPU.register.registers\[318\] top0.CPU.register.registers\[350\]
+ top0.CPU.register.registers\[382\] net850 net815 vssd1 vssd1 vccd1 vccd1 _03015_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08045__A3 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__B1 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09077_ net191 net624 net280 net258 net2331 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__a32o_1
X_06289_ top0.CPU.control.funct7\[2\] net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02946_
+ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_75_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06687__S0 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08028_ net152 net701 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__and2_1
Xhold761 top0.CPU.register.registers\[655\] vssd1 vssd1 vccd1 vccd1 net2983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold772 top0.CPU.register.registers\[146\] vssd1 vssd1 vccd1 vccd1 net2994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold750 top0.CPU.register.registers\[248\] vssd1 vssd1 vccd1 vccd1 net2972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 top0.CPU.register.registers\[778\] vssd1 vssd1 vccd1 vccd1 net3005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 net77 vssd1 vssd1 vccd1 vccd1 net3016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ top0.CPU.internalMem.pcOut\[26\] net645 _05470_ vssd1 vssd1 vccd1 vccd1 _02203_
+ sky130_fd_sc_hd__o21a_1
XFILLER_77_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10738__390 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__inv_2
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11941_ net1633 _01580_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[434\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11872_ net1564 _01511_ net1034 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09540__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08269__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08009__X _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__A3 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09769__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ net2116 _02063_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[917\]
+ sky130_fd_sc_hd__dfrtp_1
X_12355_ net2047 _01994_ net1013 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07244__A1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06678__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12286_ net1978 _01925_ net1013 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[779\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _02471_ net550 net141 vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__o21ai_1
X_10490__142 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__inv_2
XANTENNA__06507__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787__439 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__inv_2
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_109_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_34_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07330_ net443 _03973_ _03974_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531__183 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__inv_2
XFILLER_32_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08275__A3 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__A_N _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ net164 net692 net272 net259 net2342 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__a32o_1
X_07261_ net520 net523 net467 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__mux2_1
X_06212_ _02853_ _02868_ net582 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__mux2_2
X_07192_ net517 _03847_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__nand2_2
XANTENNA__06669__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06143_ _02798_ _02799_ net783 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
XANTENNA__05719__A top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06074_ _02534_ _02698_ _02717_ _02730_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_57_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_4
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _05397_ _05398_ top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1
+ _05399_ sky130_fd_sc_hd__o21ai_1
Xfanout504 net507 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
XANTENNA__05892__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09833_ top0.CPU.internalMem.pcOut\[15\] net647 vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or2_1
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
Xfanout526 _03504_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout537 _03092_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout290_A _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__RESET_B net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _05271_ top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 _05272_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_67_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06976_ top0.CPU.register.registers\[27\] top0.CPU.register.registers\[59\] top0.CPU.register.registers\[91\]
+ top0.CPU.register.registers\[123\] net913 net877 vssd1 vssd1 vccd1 vccd1 _03633_
+ sky130_fd_sc_hd__mux4_1
XFILLER_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08715_ _04581_ net3209 net359 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
X_09695_ _05204_ _05205_ _05208_ net237 net651 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__o221a_1
XANTENNA__08499__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05927_ top0.CPU.register.registers\[896\] top0.CPU.register.registers\[928\] top0.CPU.register.registers\[960\]
+ top0.CPU.register.registers\[992\] net836 net801 vssd1 vssd1 vccd1 vccd1 _02584_
+ sky130_fd_sc_hd__mux4_1
X_08646_ net193 net707 net319 net303 net2459 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a32o_1
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05858_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__inv_2
XFILLER_54_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout722_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ net2951 net188 net335 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05789_ net741 _02445_ _02440_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a21oi_4
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06825__A1_N net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09299__C _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__A3 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07528_ net527 _04162_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__nand2_1
X_07459_ _03403_ net532 net470 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__mux2_1
XANTENNA__08671__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ net182 net686 _04836_ net254 net3340 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__a32o_1
XANTENNA__07387__Y _04044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12140_ net1832 _01779_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09518__A3 top0.MMIO.WBData_i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ net1763 _01710_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[564\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold580 top0.CPU.register.registers\[772\] vssd1 vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05883__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 top0.CPU.register.registers\[776\] vssd1 vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07934__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06737__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10474__126 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__inv_2
XFILLER_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05960__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11924_ net1616 _01563_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515__167 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__inv_2
X_11855_ net1547 _01494_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[348\]
+ sky130_fd_sc_hd__dfrtp_1
X_11786_ net1478 _01425_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08662__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06673__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ net2099 _02046_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07217__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08414__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10221__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__A2 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
X_12338_ net2030 _01977_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05874__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ net1961 _01908_ net958 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06830_ _03466_ _03484_ _03485_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_52_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06761_ net762 _03415_ net752 vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__a21o_1
X_08500_ _04701_ net408 net368 net2748 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a22o_1
X_09480_ top0.MMIO.WBData_i\[1\] net139 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__or2_1
X_05712_ _02366_ _02367_ _02364_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__o21ai_1
X_06692_ top0.CPU.register.registers\[128\] top0.CPU.register.registers\[160\] top0.CPU.register.registers\[192\]
+ top0.CPU.register.registers\[224\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03349_
+ sky130_fd_sc_hd__mux4_1
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08431_ net2834 net206 net374 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__mux2_1
XANTENNA__06051__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11819__RESET_B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06009__A2_N net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ _04644_ net396 net382 net2950 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a22o_1
X_07313_ _03520_ _03969_ _03505_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08653__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ net3050 net209 net413 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XANTENNA__08591__Y _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11401__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ net485 _03890_ _03891_ net338 net244 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a221o_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251__903 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__inv_2
XFILLER_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout303_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08405__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__inv_2
XANTENNA__07759__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06126_ top0.CPU.register.registers\[14\] top0.CPU.register.registers\[46\] top0.CPU.register.registers\[78\]
+ top0.CPU.register.registers\[110\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02783_
+ sky130_fd_sc_hd__mux4_1
X_06057_ _02710_ _02713_ net737 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
Xfanout323 net326 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
Xfanout301 net302 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_8
Xfanout356 _04752_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_4
XANTENNA_fanout672_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout334 _04733_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_4
XANTENNA__06814__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _05318_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__nor2_1
Xfanout378 net380 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_8
Xfanout389 net393 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_2
X_09747_ _05252_ _05253_ _05256_ _05110_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06290__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ _03612_ _03613_ _03614_ _03615_ net764 net866 vssd1 vssd1 vccd1 vccd1 _03616_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout937_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07144__A0 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _05187_ _05191_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__o21a_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08629_ _04638_ net324 net303 net2741 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__a22o_1
XANTENNA__08892__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07695__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ net1332 _01279_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08644__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ net1263 _01210_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07998__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08434__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900__552 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__inv_2
XFILLER_109_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09773__B top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ net1815 _01762_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[616\]
+ sky130_fd_sc_hd__dfrtp_1
X_11035__687 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__inv_2
X_12054_ net1746 _01693_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[547\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08175__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06281__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_4_13_0_clk_X clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_125_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08478__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06033__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ net1599 _01546_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[400\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07686__A1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08883__B1 _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ net1530 _01477_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09013__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08635__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
X_11769_ net1461 _01408_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07989__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08650__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07101__X _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10643__295 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__inv_2
XANTENNA__09060__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07610__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08980_ _04666_ net269 net261 net2845 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__a22o_1
X_07931_ net634 _04571_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__and2_1
X_07862_ net591 _02910_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nand2_1
XANTENNA__08166__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ top0.CPU.register.registers\[781\] top0.CPU.register.registers\[813\] top0.CPU.register.registers\[845\]
+ top0.CPU.register.registers\[877\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03470_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07913__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _04957_ _05138_ net661 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__o21a_1
XANTENNA__06272__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ net948 _05057_ net125 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07793_ net449 _04447_ _04449_ _04446_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o211a_1
XANTENNA__07931__B _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06744_ _03399_ _03400_ net758 vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout253_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ top0.MMIO.WBData_i\[25\] net145 net135 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__o21a_1
XANTENNA__09204__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ top0.CPU.register.registers\[1\] top0.CPU.register.registers\[33\] top0.CPU.register.registers\[65\]
+ top0.CPU.register.registers\[97\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03332_
+ sky130_fd_sc_hd__mux4_1
X_08414_ net170 net696 net403 net380 net2688 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a32o_1
X_09394_ net942 top0.CPU.control.funct3\[1\] _02517_ vssd1 vssd1 vccd1 vccd1 _05006_
+ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_65_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08345_ net718 net217 net399 net411 net2511 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08626__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout420_A _04706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout518_A _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08276_ net509 net184 net674 net420 net2609 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a32o_1
XANTENNA__06101__A1 top0.CPU.control.rs2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ net446 _03856_ _03858_ _03875_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__D net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__inv_2
X_06109_ net781 _02761_ _02764_ _02765_ net744 vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__o221a_1
XANTENNA__10197__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ _02428_ net578 _03712_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_2
Xfanout1129 net1130 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1131 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_4
Xfanout1107 net1115 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout120 net124 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
Xfanout142 _04956_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
Xfanout164 _04622_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_2
XFILLER_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10373__25 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__inv_2
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
Xfanout186 net189 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_2
Xfanout175 net178 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_2
XFILLER_59_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06263__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08429__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06015__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12672_ clknet_leaf_82_clk _02307_ net1108 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
X_10586__238 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09409__A2 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11623_ net1315 _01262_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08617__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ net1246 _01193_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08093__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10627__279 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__inv_2
X_11485_ clknet_leaf_81_clk _01127_ net1112 vssd1 vssd1 vccd1 vccd1 top0.display.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08396__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10298_ net3027 net118 net111 _05668_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a22o_1
X_12106_ net1798 _01745_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[599\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12037_ net1729 _01676_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[530\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_89_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08148__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07591__X _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06254__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07108__A0 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06006__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06460_ _02869_ _03116_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ net2651 net184 net430 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
XANTENNA__08608__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_06391_ top0.CPU.register.registers\[413\] top0.CPU.register.registers\[445\] top0.CPU.register.registers\[477\]
+ top0.CPU.register.registers\[509\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03048_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06383__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08061_ net512 net150 net697 net435 net2369 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_60_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ _03056_ _03074_ _03667_ _03057_ _03039_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__o311a_1
XANTENNA__06190__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_69_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08963_ _04656_ net554 _04784_ net259 net3174 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__a32o_1
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07914_ _04442_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__and3_2
XFILLER_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08894_ net721 net196 net278 net283 net2661 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1008_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ net713 net211 vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__and2_1
XANTENNA__06245__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07776_ _03223_ _03224_ _03242_ _03941_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_67_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09515_ top0.MMIO.WBData_i\[28\] top0.MMIO.WBData_i\[26\] top0.MMIO.WBData_i\[11\]
+ _02355_ net137 vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a41o_1
XANTENNA__08847__A0 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06727_ _03280_ _03380_ _03281_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o21a_1
X_09446_ _04933_ _05036_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout635_A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06658_ _03313_ _03314_ net757 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ net2545 _04530_ net606 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__mux2_1
X_06589_ _03177_ _03198_ _03244_ _03245_ _03174_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout802_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10418__70 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__inv_2
X_08328_ net3098 net409 net386 _04517_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XANTENNA__08614__A3 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ net500 net206 net671 net418 net2267 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a32o_1
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09024__A0 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06181__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08378__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ net2 net655 net594 top0.MMIO.WBData_i\[0\] vssd1 vssd1 vccd1 vccd1 _02267_
+ sky130_fd_sc_hd__o22a_1
X_10971__623 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__inv_2
XFILLER_106_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10152_ top0.display.delayctr\[24\] top0.display.delayctr\[25\] _05604_ vssd1 vssd1
+ vccd1 vccd1 _05613_ sky130_fd_sc_hd__or3_1
X_10083_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__nand2_1
XANTENNA__09543__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 top0.CPU.register.registers\[28\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07852__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__A0 _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11504__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05995__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11147__799 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__inv_2
XFILLER_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06313__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12655_ clknet_leaf_71_clk _02290_ net1119 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09263__B1 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12586_ clknet_leaf_84_clk _02221_ net1110 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11606_ net1298 _01245_ net982 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ net1229 _01176_ net1050 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 top0.CPU.intMemAddr\[9\] vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11468_ clknet_leaf_67_clk _01116_ net1103 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.funct7\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09015__B1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ clknet_leaf_57_clk _01047_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11050__702 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1109 top0.CPU.register.registers\[274\] vssd1 vssd1 vccd1 vccd1 net3331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05960_ net584 _02614_ _02615_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a21boi_2
Xclkbuf_leaf_2_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05891_ top0.CPU.register.registers\[3\] top0.CPU.register.registers\[35\] top0.CPU.register.registers\[67\]
+ top0.CPU.register.registers\[99\] net831 net796 vssd1 vssd1 vccd1 vccd1 _02548_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06227__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06001__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ net489 _04025_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__or2_1
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08829__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ _04052_ _04061_ net488 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__mux2_1
X_06512_ top0.CPU.register.registers\[147\] top0.CPU.register.registers\[179\] top0.CPU.register.registers\[211\]
+ top0.CPU.register.registers\[243\] net940 net906 vssd1 vssd1 vccd1 vccd1 _03169_
+ sky130_fd_sc_hd__mux4_1
X_09300_ _04865_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__or2_1
X_10352__4 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__inv_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08593__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07492_ _04147_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and2_1
X_09231_ _04871_ _04884_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__o21a_1
X_06443_ top0.CPU.register.registers\[662\] top0.CPU.register.registers\[694\] top0.CPU.register.registers\[726\]
+ top0.CPU.register.registers\[758\] net923 net889 vssd1 vssd1 vccd1 vccd1 _03100_
+ sky130_fd_sc_hd__mux4_1
X_06374_ net754 _03030_ net860 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__o21ai_1
X_09162_ top0.CPU.register.registers\[49\] net564 vssd1 vssd1 vccd1 vccd1 _04845_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08057__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08113_ net2840 _04504_ net429 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09093_ net948 _04688_ _04732_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__or3_4
XANTENNA__09006__A0 _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_A _04618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 top0.CPU.register.registers\[927\] vssd1 vssd1 vccd1 vccd1 net3132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 top0.CPU.register.registers\[167\] vssd1 vssd1 vccd1 vccd1 net3143 sky130_fd_sc_hd__dlygate4sd3_1
X_10955__607 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__inv_2
XANTENNA__07937__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net3032 net440 _04651_ net502 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
Xhold943 top0.CPU.register.registers\[144\] vssd1 vssd1 vccd1 vccd1 net3165 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold932 top0.CPU.register.registers\[284\] vssd1 vssd1 vccd1 vccd1 net3154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 top0.CPU.register.registers\[151\] vssd1 vssd1 vccd1 vccd1 net3176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 top0.CPU.register.registers\[389\] vssd1 vssd1 vccd1 vccd1 net3220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 top0.CPU.register.registers\[397\] vssd1 vssd1 vccd1 vccd1 net3209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_clkbuf_4_1_0_clk_X clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 top0.CPU.register.registers\[145\] vssd1 vssd1 vccd1 vccd1 net3198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 top0.CPU.register.registers\[981\] vssd1 vssd1 vccd1 vccd1 net3187 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08780__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ net585 _02981_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__nor2_1
XANTENNA__06240__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net180 net708 net277 net265 net2518 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout752_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _04517_ net552 _04759_ net282 net3045 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__a32o_1
X_10849__501 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__inv_2
XANTENNA__08487__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ net591 _03009_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__nand2_1
XFILLER_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08532__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07740__B1 _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _02852_ net447 _03739_ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__o31a_1
XANTENNA__09088__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08707__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ net3408 net599 net132 _05030_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__o22a_1
XFILLER_9_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ net2132 _02079_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[933\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06059__B1 _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12371_ net2063 _02010_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08442__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ net2734 net123 net116 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a21o_1
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__B1 _04175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08220__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ _02887_ _05577_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08771__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06209__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ top0.display.delayctr\[6\] _05542_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08523__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05968__S0 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08826__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__12544__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ clknet_leaf_71_clk _02273_ net1120 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06393__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_135_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12569_ clknet_leaf_57_clk _02208_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06145__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 top0.CPU.register.registers\[73\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 top0.CPU.internalMem.load2Ct\[1\] vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
X_06090_ net778 _02742_ _02745_ _02746_ net744 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__o221a_1
XANTENNA__06661__A _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06696__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 top0.CPU.register.registers\[298\] vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07476__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold228 top0.CPU.register.registers\[736\] vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09003__A3 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_4
Xfanout719 net722 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
X_08800_ _04708_ net317 net286 net3072 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a22o_1
XANTENNA__06448__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _05284_ _05286_ top0.CPU.internalMem.pcOut\[11\] vssd1 vssd1 vccd1 vccd1
+ _05287_ sky130_fd_sc_hd__a21o_1
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06992_ top0.CPU.register.registers\[154\] top0.CPU.register.registers\[186\] top0.CPU.register.registers\[218\]
+ top0.CPU.register.registers\[250\] net908 net874 vssd1 vssd1 vccd1 vccd1 _03649_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08762__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ _04673_ net324 net296 net2666 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
XANTENNA__07970__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05943_ top0.CPU.register.registers\[513\] top0.CPU.register.registers\[545\] top0.CPU.register.registers\[577\]
+ top0.CPU.register.registers\[609\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02600_
+ sky130_fd_sc_hd__mux4_1
X_08662_ _04654_ net324 net299 net2837 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a22o_1
XANTENNA__08514__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05724__B top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09911__S net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05874_ _02527_ _02528_ _02530_ _02529_ net784 net737 vssd1 vssd1 vccd1 vccd1 _02531_
+ sky130_fd_sc_hd__mux4_1
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ net479 _03317_ net444 _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__o31a_1
X_08593_ net634 _04481_ net327 vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__and3_2
XANTENNA__06620__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout166_A _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07544_ _04199_ _04200_ _03704_ _03829_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__a211o_1
XANTENNA__05740__A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ _02962_ _03637_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09214_ net770 top0.CPU.intMemAddr\[31\] _04874_ _04875_ vssd1 vssd1 vccd1 vccd1
+ _04876_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout333_A _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06426_ top0.CPU.register.registers\[791\] top0.CPU.register.registers\[823\] top0.CPU.register.registers\[855\]
+ top0.CPU.register.registers\[887\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03083_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09778__A1 top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ net949 _04705_ _04732_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__or3_4
X_06357_ _03010_ _03011_ _03012_ _03013_ net730 net740 vssd1 vssd1 vccd1 vccd1 _03014_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09778__B2 top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09076_ net193 net622 _04818_ net257 net3272 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__a32o_1
XANTENNA__05739__X _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06288_ net580 _02928_ _02943_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a21boi_1
XANTENNA__06687__S1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08027_ net3088 net440 _04644_ net500 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a22o_1
Xhold740 top0.CPU.register.registers\[851\] vssd1 vssd1 vccd1 vccd1 net2962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 top0.CPU.register.registers\[912\] vssd1 vssd1 vccd1 vccd1 net2973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 top0.CPU.register.registers\[423\] vssd1 vssd1 vccd1 vccd1 net2995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 top0.CPU.register.registers\[122\] vssd1 vssd1 vccd1 vccd1 net2984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 top0.CPU.register.registers\[252\] vssd1 vssd1 vccd1 vccd1 net3006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 top0.CPU.register.registers\[280\] vssd1 vssd1 vccd1 vccd1 net3017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net235 _05465_ _05466_ _05469_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a31o_1
XFILLER_77_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07961__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _04647_ net274 net264 net2582 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08505__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11940_ net1632 _01579_ net993 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[433\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06516__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11871_ net1563 _01510_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[364\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05921__Y _02578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06375__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ net2115 _02062_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06127__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12354_ net2046 _01993_ net1046 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06481__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08992__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12285_ net1977 _01924_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[778\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06204__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ net3418 net665 net662 _05582_ _05585_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a221o_1
XANTENNA__05963__C1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06507__A1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10049_ top0.display.delayctr\[0\] top0.display.delayctr\[1\] top0.display.delayctr\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__or3_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11162__814 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__inv_2
XANTENNA__06602__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203__855 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__inv_2
X_07260_ _03094_ _03114_ _03915_ net344 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__a31o_1
XANTENNA__06943__X _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08590__B net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06211_ net742 _02867_ _02862_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a21oi_2
X_07191_ _03747_ _03846_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__nor2_1
XANTENNA__06118__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06669__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06142_ top0.CPU.register.registers\[913\] top0.CPU.register.registers\[945\] top0.CPU.register.registers\[977\]
+ top0.CPU.register.registers\[1009\] net828 net793 vssd1 vssd1 vccd1 vccd1 _02799_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08983__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06073_ top0.CPU.control.funct7\[5\] _02518_ _02729_ net581 vssd1 vssd1 vccd1 vccd1
+ _02730_ sky130_fd_sc_hd__a22o_2
X_09901_ net585 _02851_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_57_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout505 net507 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout516 _02405_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
X_09832_ top0.CPU.internalMem.pcOut\[15\] _05325_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05335_ sky130_fd_sc_hd__a21oi_1
Xfanout527 _03463_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_4
Xfanout538 _03073_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06746__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08735__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _02392_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_8
XANTENNA__05735__A top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ net588 _04016_ net234 net229 _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__a41oi_2
XTAP_TAPCELL_ROW_70_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10770__422 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__inv_2
XANTENNA__06330__S net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06975_ top0.CPU.register.registers\[155\] top0.CPU.register.registers\[187\] top0.CPU.register.registers\[219\]
+ top0.CPU.register.registers\[251\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03632_
+ sky130_fd_sc_hd__mux4_1
X_08714_ _04576_ net3064 net358 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__mux2_1
X_09694_ _05206_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__or2_1
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05926_ top0.CPU.register.registers\[768\] top0.CPU.register.registers\[800\] top0.CPU.register.registers\[832\]
+ top0.CPU.register.registers\[864\] net836 net801 vssd1 vssd1 vccd1 vccd1 _02583_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09160__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811__463 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__inv_2
X_05857_ net581 _02513_ _02512_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout450_A _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ _04651_ net316 net302 net2517 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a22o_1
XFILLER_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ net3035 _04586_ net336 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07527_ _04179_ _04180_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__and3_1
XFILLER_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05788_ _02441_ _02442_ _02443_ _02444_ net724 net776 vssd1 vssd1 vccd1 vccd1 _02445_
+ sky130_fd_sc_hd__mux4_2
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06357__S0 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07458_ net482 _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__and2_1
X_07389_ net342 _03967_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nand2_1
XANTENNA__06682__B1 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06409_ net863 _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__nor2_1
XANTENNA__07668__Y _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ top0.CPU.register.registers\[74\] net573 net559 vssd1 vssd1 vccd1 vccd1 _04836_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07548__C_N _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09059_ top0.CPU.register.registers\[120\] net568 vssd1 vssd1 vccd1 vccd1 _04813_
+ sky130_fd_sc_hd__or2_1
X_12070_ net1762 _01709_ net1128 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08720__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 net63 vssd1 vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 top0.CPU.register.registers\[46\] vssd1 vssd1 vccd1 vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold592 top0.CPU.register.registers\[190\] vssd1 vssd1 vccd1 vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09923__B2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08187__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06737__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05960__A2 _02614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net1615 _01562_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[416\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06596__S0 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ net1546 _01493_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07071__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ net1477 _01424_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[278\]
+ sky130_fd_sc_hd__dfrtp_1
X_12406_ net2098 _02045_ net988 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[899\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11771__RESET_B net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ net2029 _01976_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10221__B2 top0.MMIO.WBData_i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379__31 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__inv_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_1
XANTENNA__08965__A2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ net1960 _01907_ net967 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[761\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08178__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754__406 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__inv_2
XANTENNA__08193__A3 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net1891 _01838_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[692\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06150__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ net872 _03416_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__and2_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_05711_ _02366_ _02367_ _02364_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__o21a_1
XANTENNA__10288__A1 _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07770__A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06691_ net866 _03343_ net859 vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08430_ net2807 _04528_ net373 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XANTENNA__08350__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648__300 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__inv_2
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08102__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _04643_ net386 net381 net2770 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a22o_1
X_07312_ _03567_ _03967_ _03521_ _03541_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__a211o_1
X_08292_ net2723 _04504_ net413 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
X_07243_ net341 _03897_ _03898_ net442 _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o221a_1
X_11290__942 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__inv_2
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ net466 net518 vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__or2_1
X_06125_ top0.CPU.register.registers\[142\] top0.CPU.register.registers\[174\] top0.CPU.register.registers\[206\]
+ top0.CPU.register.registers\[238\] net835 net801 vssd1 vssd1 vccd1 vccd1 _02782_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08956__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06056_ _02711_ _02712_ net728 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1038_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10497__149 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__inv_2
XFILLER_87_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08169__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 _04737_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
Xfanout302 net304 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331__983 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__inv_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_8
Xfanout324 net326 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
X_09815_ top0.CPU.internalMem.pcOut\[14\] _05317_ vssd1 vssd1 vccd1 vccd1 _05319_
+ sky130_fd_sc_hd__nor2_1
XFILLER_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_8
Xfanout346 net348 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08184__A3 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 _04728_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
XANTENNA__06814__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _05254_ _05255_ net650 vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__o21a_1
XANTENNA__09669__B1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06958_ top0.CPU.register.registers\[280\] top0.CPU.register.registers\[312\] top0.CPU.register.registers\[344\]
+ top0.CPU.register.registers\[376\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03615_
+ sky130_fd_sc_hd__mux4_1
X_09677_ _05187_ _05191_ net241 vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09133__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05909_ net725 _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__or2_1
XANTENNA__08341__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ net710 _04738_ net304 net2783 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__a22o_1
X_06889_ top0.CPU.register.registers\[776\] top0.CPU.register.registers\[808\] top0.CPU.register.registers\[840\]
+ top0.CPU.register.registers\[872\] net929 net895 vssd1 vssd1 vccd1 vccd1 _03546_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout832_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ net2999 _04492_ net334 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
X_11570_ net1262 _01209_ net1053 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08715__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__11529__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08016__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06502__S0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09546__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12122_ net1814 _01761_ net1006 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[615\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08450__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ net1745 _01692_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[546\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07907__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout880 net882 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout891 net892 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09124__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ net1598 _01545_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[399\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06569__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11837_ net1529 _01476_ net1024 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[330\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_44_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ net1460 _01407_ net1044 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06934__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07843__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274__926 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__inv_2
X_11699_ net1391 _01338_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[192\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11315__967 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07930_ top0.CPU.internalMem.pcOut\[15\] net642 _04569_ _04570_ vssd1 vssd1 vccd1
+ vccd1 _04571_ sky130_fd_sc_hd__a22o_2
XFILLER_69_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07484__B _03112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168__820 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__inv_2
X_07861_ _04400_ net231 net226 vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__and3_1
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06812_ top0.CPU.register.registers\[909\] top0.CPU.register.registers\[941\] top0.CPU.register.registers\[973\]
+ top0.CPU.register.registers\[1005\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03469_
+ sky130_fd_sc_hd__mux4_1
XFILLER_84_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ _02551_ _05007_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__nor2_1
X_07792_ net483 _04109_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a21o_1
X_09531_ net951 _05070_ net125 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XANTENNA__09115__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06743_ top0.CPU.register.registers\[262\] top0.CPU.register.registers\[294\] top0.CPU.register.registers\[326\]
+ top0.CPU.register.registers\[358\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03400_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08323__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11209__861 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__inv_2
XANTENNA__05732__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ net132 net134 _05049_ net599 net3441 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__o32a_1
XFILLER_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07677__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06674_ top0.CPU.register.registers\[129\] top0.CPU.register.registers\[161\] top0.CPU.register.registers\[193\]
+ top0.CPU.register.registers\[225\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03331_
+ sky130_fd_sc_hd__mux4_1
X_09393_ _04988_ _05003_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nand2b_1
X_10882__534 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__inv_2
X_08413_ net171 net692 net390 net377 net2294 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a32o_1
X_08344_ net720 net179 net401 net411 net2486 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08626__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08275_ net506 net188 net672 net419 net2287 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a32o_1
XANTENNA__06732__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout413_A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923__575 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__inv_2
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07226_ _03005_ _03054_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__xnor2_1
X_07157_ net455 _03813_ _03811_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21a_1
XANTENNA__08929__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06108_ net787 _02762_ net740 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a21o_1
X_07088_ _02431_ _03742_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout782_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_4
X_06039_ _02692_ _02693_ _02694_ _02695_ net728 net778 vssd1 vssd1 vccd1 vccd1 _02696_
+ sky130_fd_sc_hd__mux4_1
Xfanout121 net123 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1108 net1115 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
Xfanout143 _04953_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
Xfanout132 _05024_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout165 _04622_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
Xfanout154 net156 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
Xfanout198 _04572_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XANTENNA__06799__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 net189 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
Xfanout176 net178 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07365__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ top0.CPU.internalMem.pcOut\[7\] _05228_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__and2_1
XANTENNA__05915__A2 _02563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06325__C1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12671_ clknet_leaf_91_clk _02306_ net1085 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
X_11622_ net1314 _01261_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08617__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06971__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08445__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002__654 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__inv_2
X_11553_ net1245 _01192_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_11484_ clknet_leaf_81_clk _01126_ net1109 vssd1 vssd1 vccd1 vccd1 top0.display.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xteam_07_1190 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] team_07_1190/LO sky130_fd_sc_hd__conb_1
XANTENNA__10188__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12105_ net1797 _01744_ net1071 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[598\]
+ sky130_fd_sc_hd__dfrtp_1
X_10297_ net144 _05611_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07872__X _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12036_ net1728 _01675_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[529\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07356__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08553__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07108__A1 _03221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866__518 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__inv_2
X_10907__559 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__inv_2
XANTENNA__08608__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610__262 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__inv_2
X_06390_ top0.CPU.register.registers\[285\] top0.CPU.register.registers\[317\] top0.CPU.register.registers\[349\]
+ top0.CPU.register.registers\[381\] net926 net892 vssd1 vssd1 vccd1 vccd1 _03047_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07479__B _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ net946 _02399_ net699 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__nand3_1
X_07011_ _03056_ _03074_ _03667_ _03057_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__o31a_1
XANTENNA__06190__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07495__A _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08792__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ top0.CPU.register.registers\[188\] net566 vssd1 vssd1 vccd1 vccd1 _04784_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12239__RESET_B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08893_ net718 net200 _04766_ net283 net3264 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__a32o_1
X_07913_ net719 net508 net203 net547 net2543 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a32o_1
XANTENNA__08544__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07844_ top0.CPU.internalMem.pcOut\[28\] net638 net634 _04497_ vssd1 vssd1 vccd1
+ vccd1 _04498_ sky130_fd_sc_hd__o211a_2
XANTENNA__05743__A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ net343 _03914_ _04422_ _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a31o_1
XFILLER_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_27_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09514_ _05080_ _05081_ _05082_ _05088_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__and4_1
X_06726_ _03282_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__nor2_1
XFILLER_37_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09445_ net131 _05038_ net133 net597 net3412 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__o32a_1
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06657_ top0.CPU.register.registers\[258\] top0.CPU.register.registers\[290\] top0.CPU.register.registers\[322\]
+ top0.CPU.register.registers\[354\] net916 net882 vssd1 vssd1 vccd1 vccd1 _03314_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout530_A _03379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ net2382 _04535_ net607 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__mux2_1
X_06588_ _03157_ net535 _03196_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ net3000 net409 net385 _04511_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
XANTENNA__08075__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06861__X _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ net3135 net417 _04714_ net494 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
XFILLER_20_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout997_A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06181__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07209_ net466 _03770_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__nand2_1
X_10433__85 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__inv_2
X_10220_ net767 net657 top0.wishbone0.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05648_
+ sky130_fd_sc_hd__or3b_1
X_08189_ net495 net153 net617 net426 net2386 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ net141 _05611_ net660 vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09109__B net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ top0.display.delayctr\[10\] _05554_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553__205 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__inv_2
XANTENNA__07338__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06101__X _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_122_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05995__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06849__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05940__X _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ clknet_leaf_74_clk _02289_ net1124 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09446__A_N _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12585_ clknet_leaf_83_clk _02220_ net1110 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11605_ net1297 _01244_ net969 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06077__A1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ net1228 _01175_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_13_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11467_ clknet_leaf_74_clk _01115_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.rs2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11398_ clknet_leaf_59_clk _01046_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08774__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10349_ net2250 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08526__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ net1711 _01658_ net1059 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[512\]
+ sky130_fd_sc_hd__dfrtp_1
X_11130__782 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__inv_2
XANTENNA__06001__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05890_ top0.CPU.register.registers\[131\] top0.CPU.register.registers\[163\] top0.CPU.register.registers\[195\]
+ top0.CPU.register.registers\[227\] net831 net796 vssd1 vssd1 vccd1 vccd1 _02547_
+ sky130_fd_sc_hd__mux4_1
XFILLER_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08541__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _03705_ _04216_ _04128_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__a21bo_1
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06511_ _03166_ _03167_ net873 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__mux2_1
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08593__B _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ net607 _04889_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__or3_1
X_07491_ _02810_ _02811_ _03221_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_62_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06442_ _03097_ _03098_ net764 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
XFILLER_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06373_ _03028_ _03029_ net873 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
X_09161_ _04730_ _04731_ net250 net2875 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__a22o_1
XANTENNA__08057__A2 _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09092_ net155 net617 _04821_ net256 net3226 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a32o_1
XANTENNA__07265__A0 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08112_ net3183 net211 net429 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
X_08043_ net221 net705 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and2_1
Xhold922 top0.CPU.register.registers\[286\] vssd1 vssd1 vccd1 vccd1 net3144 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10994__646 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__inv_2
XANTENNA_fanout209_A _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold911 top0.CPU.register.registers\[55\] vssd1 vssd1 vccd1 vccd1 net3133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07937__B _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold900 top0.CPU.register.registers\[442\] vssd1 vssd1 vccd1 vccd1 net3122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 top0.CPU.register.registers\[531\] vssd1 vssd1 vccd1 vccd1 net3177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05738__A top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold944 top0.CPU.register.registers\[980\] vssd1 vssd1 vccd1 vccd1 net3166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A1 _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 top0.CPU.register.registers\[256\] vssd1 vssd1 vccd1 vccd1 net3155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 top0.CPU.register.registers\[266\] vssd1 vssd1 vccd1 vccd1 net3210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12632__Q top0.MMIO.WBData_i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold966 top0.CPU.register.registers\[141\] vssd1 vssd1 vccd1 vccd1 net3188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09994_ _05437_ _05480_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a21o_1
Xhold977 top0.CPU.register.registers\[129\] vssd1 vssd1 vccd1 vccd1 net3199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07953__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__A2 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold999 top0.CPU.register.registers\[38\] vssd1 vssd1 vccd1 vccd1 net3221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06240__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ net182 net708 _04780_ net265 net3307 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__a32o_1
XANTENNA__08517__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ top0.CPU.register.registers\[249\] net564 vssd1 vssd1 vccd1 vccd1 _04759_
+ sky130_fd_sc_hd__or2_1
X_07827_ _03852_ net231 net226 vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__and3_1
XFILLER_57_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10888__540 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__inv_2
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout745_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ _02852_ _03150_ net341 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06709_ top0.CPU.register.registers\[900\] top0.CPU.register.registers\[932\] top0.CPU.register.registers\[964\]
+ top0.CPU.register.registers\[996\] net916 net882 vssd1 vssd1 vccd1 vccd1 _03366_
+ sky130_fd_sc_hd__mux4_1
X_07689_ _03427_ _03444_ _04321_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10929__581 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__inv_2
XANTENNA_fanout912_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ top0.MMIO.WBData_i\[10\] net146 _05028_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__o21a_1
XFILLER_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ net2585 _04616_ net609 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ net2062 _02009_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06059__B2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08723__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11073__725 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__inv_2
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08024__A _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ net2708 net123 net116 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a21o_1
XFILLER_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08756__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06231__A1 _02887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ net3428 net663 net602 _05598_ _05595_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a221o_1
X_11114__766 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__inv_2
XANTENNA__08220__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08508__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ top0.display.delayctr\[6\] _05542_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__or2_1
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09720__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05968__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__A top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008__660 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__inv_2
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ clknet_leaf_75_clk _02272_ net1125 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09236__A1 top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06393__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07103__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681__333 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__inv_2
XFILLER_12_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12568_ clknet_leaf_57_clk _02207_ net1092 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08995__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06145__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11519_ net1211 _01158_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold207 top0.CPU.register.registers\[841\] vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_12499_ net2191 _02138_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[992\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold229 top0.CPU.intMemAddr\[26\] vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_10722__374 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__inv_2
Xhold218 top0.CPU.register.registers\[995\] vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08747__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 net711 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05992__S net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06222__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08211__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07970__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ net749 _03647_ net858 vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08762__A3 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ net624 _04738_ net296 net2621 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a22o_1
X_05942_ top0.CPU.register.registers\[641\] top0.CPU.register.registers\[673\] top0.CPU.register.registers\[705\]
+ top0.CPU.register.registers\[737\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02599_
+ sky130_fd_sc_hd__mux4_1
X_08661_ net699 _04738_ net300 net2579 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a22o_1
XANTENNA__09172__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05724__C top0.CPU.Op\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05873_ top0.CPU.register.registers\[11\] top0.CPU.register.registers\[43\] top0.CPU.register.registers\[75\]
+ top0.CPU.register.registers\[107\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02530_
+ sky130_fd_sc_hd__mux4_1
XFILLER_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06081__S0 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ net479 _03317_ net339 vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a21o_1
X_08592_ _02404_ _04732_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__nor2_4
XFILLER_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07543_ _02983_ _03883_ _03073_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__or3b_1
XANTENNA__05740__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06289__A1 top0.CPU.control.funct7\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _02962_ net521 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__and2_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout159_A _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ top0.CPU.intMemAddr\[30\] top0.CPU.intMemAddr\[29\] top0.CPU.intMemAddr\[28\]
+ top0.CPU.intMemAddr\[27\] vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__or4_1
X_06425_ net862 _03081_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout326_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ net155 net682 _04841_ net252 net3275 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a32o_1
X_06356_ top0.CPU.register.registers\[542\] top0.CPU.register.registers\[574\] top0.CPU.register.registers\[606\]
+ top0.CPU.register.registers\[638\] net853 net818 vssd1 vssd1 vccd1 vccd1 _03013_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09778__A2 top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057__709 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__inv_2
X_09075_ top0.CPU.register.registers\[109\] net572 net558 vssd1 vssd1 vccd1 vccd1
+ _04818_ sky130_fd_sc_hd__o21a_1
XANTENNA__08986__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout114_X net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06287_ net580 _02928_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a21bo_2
XANTENNA__07159__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ net207 net705 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__and2_1
Xhold730 top0.CPU.register.registers\[501\] vssd1 vssd1 vccd1 vccd1 net2952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 top0.CPU.register.registers\[735\] vssd1 vssd1 vccd1 vccd1 net2974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout695_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold763 net42 vssd1 vssd1 vccd1 vccd1 net2985 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold741 top0.CPU.register.registers\[246\] vssd1 vssd1 vccd1 vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
X_10403__55 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__inv_2
Xhold796 top0.CPU.register.registers\[862\] vssd1 vssd1 vccd1 vccd1 net3018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 top0.CPU.register.registers\[134\] vssd1 vssd1 vccd1 vccd1 net3007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06998__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold774 top0.CPU.register.registers\[657\] vssd1 vssd1 vccd1 vccd1 net2996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07961__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net235 _05467_ _05468_ net645 vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout862_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06299__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ _04646_ net273 net264 net2736 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__a22o_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09163__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ net213 net3339 net353 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__mux2_1
XANTENNA__08910__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ net1562 _01509_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[363\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665__317 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06375__S1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ net2114 _02061_ net1127 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[915\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706__358 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__inv_2
XANTENNA__08453__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06127__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12353_ net2045 _01992_ net1061 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[846\]
+ sky130_fd_sc_hd__dfrtp_1
X_12284_ net1976 _01923_ net1025 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06204__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10559__211 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__inv_2
XFILLER_136_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10117_ _05583_ _05584_ net601 vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10048_ top0.display.delayctr\[1\] net664 net602 _05532_ _05135_ vssd1 vssd1 vccd1
+ vccd1 _02210_ sky130_fd_sc_hd__a221o_1
XFILLER_48_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__09154__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08901__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 top0.CPU.register.registers\[737\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06063__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05810__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11999_ net1691 _01638_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[492\]
+ sky130_fd_sc_hd__dfrtp_1
X_11242__894 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__inv_2
XANTENNA__08680__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06210_ _02863_ _02864_ _02866_ _02865_ net783 net736 vssd1 vssd1 vccd1 vccd1 _02867_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08871__B net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07190_ net451 _03748_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__or2_2
XANTENNA__06118__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__A1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06141_ top0.CPU.register.registers\[785\] top0.CPU.register.registers\[817\] top0.CPU.register.registers\[849\]
+ top0.CPU.register.registers\[881\] net827 net792 vssd1 vssd1 vccd1 vccd1 _02798_
+ sky130_fd_sc_hd__mux4_1
X_06072_ _02723_ _02728_ net743 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_4
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08983__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09900_ net586 _04421_ net234 net229 vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__and4_1
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_2
XANTENNA__06611__S net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ top0.CPU.internalMem.pcOut\[15\] _05325_ net239 vssd1 vssd1 vccd1 vccd1 _05334_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkload13_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout539 _03037_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
Xfanout528 _03443_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
X_09762_ top0.CPU.control.funct7\[5\] net631 _02453_ vssd1 vssd1 vccd1 vccd1 _05270_
+ sky130_fd_sc_hd__and3_1
X_06974_ net753 _03630_ top0.CPU.decoder.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ _03631_ sky130_fd_sc_hd__o21ai_1
X_08713_ _04571_ net3243 net359 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
XFILLER_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07790__X _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05925_ _02580_ _02581_ net733 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__mux2_1
X_09693_ top0.CPU.internalMem.pcOut\[4\] top0.CPU.internalMem.pcOut\[3\] net768 vssd1
+ vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and3_1
XFILLER_82_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout276_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net198 net709 net325 net303 net2681 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a32o_1
XANTENNA__06054__S0 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05856_ net941 _02474_ _02472_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a21o_1
XFILLER_54_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ net2818 _04581_ net335 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XANTENNA__05801__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05787_ top0.CPU.register.registers\[279\] top0.CPU.register.registers\[311\] top0.CPU.register.registers\[343\]
+ top0.CPU.register.registers\[375\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02444_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_85_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07526_ _04083_ _04096_ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or3_1
XANTENNA__07459__A0 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06357__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07457_ _04036_ _04038_ net345 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__mux2_1
X_07388_ _03385_ _03407_ _03409_ _03559_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__o31a_1
X_06408_ _03063_ _03064_ net759 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XANTENNA__08959__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ net186 net683 _04835_ net253 net3342 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a32o_1
X_06339_ top0.CPU.register.registers\[413\] top0.CPU.register.registers\[445\] top0.CPU.register.registers\[477\]
+ top0.CPU.register.registers\[509\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02996_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07965__X _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09058_ _04678_ net552 _04812_ net255 net3150 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ top0.CPU.internalMem.pcOut\[0\] net640 _04633_ _04634_ net635 vssd1 vssd1
+ vccd1 vccd1 _04635_ sky130_fd_sc_hd__o221a_2
XANTENNA__08187__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 top0.CPU.register.registers\[731\] vssd1 vssd1 vccd1 vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 top0.CPU.register.registers\[1014\] vssd1 vssd1 vccd1 vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11388__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 top0.CPU.register.registers\[52\] vssd1 vssd1 vccd1 vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 top0.CPU.register.registers\[945\] vssd1 vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06293__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185__837 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__inv_2
XANTENNA__11436__Q top0.CPU.intMem_out\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ net1614 _01561_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[415\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11226__878 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__inv_2
XANTENNA__06596__S1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11853_ net1545 _01492_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[346\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ net1476 _01423_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[277\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08111__A1 _04492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08662__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07870__B1 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06673__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079__731 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__inv_2
X_12405_ net2097 _02044_ net978 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[898\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08414__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10221__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
X_12336_ net2028 _01975_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[829\]
+ sky130_fd_sc_hd__dfrtp_1
X_12267_ net1959 _01906_ net1072 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[760\]
+ sky130_fd_sc_hd__dfrtp_1
X_12198_ net1890 _01837_ net1128 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[691\]
+ sky130_fd_sc_hd__dfrtp_1
X_10394__46 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__inv_2
X_10793__445 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__inv_2
XANTENNA__08212__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__06284__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10834__486 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__inv_2
XANTENNA__08866__B _04732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05710_ top0.CPU.internalMem.state\[1\] top0.CPU.internalMem.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _02367_ sky130_fd_sc_hd__or2_1
XANTENNA__06036__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ net753 _03346_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__nor2_1
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08350__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ _04642_ net385 net381 net2958 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a22o_1
X_07311_ _03567_ _03967_ _03541_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08102__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08653__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ net2852 _04498_ net413 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__mux2_1
X_07242_ _02983_ net538 net446 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__or3_1
X_10728__380 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__inv_2
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ _03740_ _03828_ _03829_ net443 _03827_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a221o_1
XANTENNA__08405__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06124_ net739 _02780_ net771 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10212__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__A3 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06055_ top0.CPU.register.registers\[8\] top0.CPU.register.registers\[40\] top0.CPU.register.registers\[72\]
+ top0.CPU.register.registers\[104\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02712_
+ sky130_fd_sc_hd__mux4_1
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08169__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout314 net317 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_2
Xfanout336 _04733_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_4
X_09814_ top0.CPU.internalMem.pcOut\[14\] _05317_ vssd1 vssd1 vccd1 vccd1 _05318_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11481__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06275__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09652__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _04727_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_8
Xfanout358 net360 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout560_A _04754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ top0.CPU.internalMem.pcOut\[8\] _05240_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06957_ top0.CPU.register.registers\[408\] top0.CPU.register.registers\[440\] top0.CPU.register.registers\[472\]
+ top0.CPU.register.registers\[504\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03614_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05752__Y _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ _05189_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nand2b_1
X_06888_ _03543_ _03544_ net760 vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__mux2_1
XANTENNA__09133__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05908_ top0.CPU.register.registers\[386\] top0.CPU.register.registers\[418\] top0.CPU.register.registers\[450\]
+ top0.CPU.register.registers\[482\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02565_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08341__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ net947 net710 _04734_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__nand3_1
XFILLER_82_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05839_ net582 _02495_ _02494_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__o21ai_4
XFILLER_55_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout825_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ net2932 _04487_ net335 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08644__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ _04690_ net405 net367 net2726 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
X_07509_ net454 net530 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_25_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10480__132 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__inv_2
XANTENNA__08016__B net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10203__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10777__429 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__inv_2
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07855__B _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ net1813 _01760_ net979 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[614\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold390 top0.CPU.register.registers\[222\] vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
X_10521__173 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__inv_2
XANTENNA__06251__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ net1744 _01691_ net957 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[545\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10281__B _05169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 top0.CPU.decoder.instruction\[17\] vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net907 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_125_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 top0.CPU.register.registers\[237\] vssd1 vssd1 vccd1 vccd1 net3312 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06569__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11905_ net1597 _01544_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[398\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12357__RESET_B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08883__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11836_ net1528 _01475_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08096__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net1459 _01406_ net971 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[260\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08635__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06493__Y _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10439__91 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__inv_2
X_11698_ net1390 _01337_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__A3 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net2011 _01958_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07359__C1 _04015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07860_ net3321 net546 net491 _04511_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XANTENNA__06257__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06582__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ net540 _02770_ _03446_ _02750_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__a211o_1
XANTENNA__07374__A2 _04030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07781__A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07791_ net488 _04114_ _03841_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a21o_1
X_09530_ net953 _05072_ net125 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06742_ top0.CPU.register.registers\[390\] top0.CPU.register.registers\[422\] top0.CPU.register.registers\[454\]
+ top0.CPU.register.registers\[486\] net918 net884 vssd1 vssd1 vccd1 vccd1 _03399_
+ sky130_fd_sc_hd__mux4_1
X_09461_ top0.MMIO.WBData_i\[24\] _05041_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06397__A _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06334__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06673_ net749 _03325_ _03328_ _03329_ net745 vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__a221o_1
X_09392_ _02338_ net629 _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07005__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ net177 net691 net390 net378 net2662 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a32o_1
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ net720 net185 net402 net411 net2390 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a32o_1
XANTENNA__09823__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ net515 net190 net677 net420 net2365 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10464__116 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__inv_2
XANTENNA__06732__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07225_ _03878_ _03881_ net487 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__mux2_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1050_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ _02579_ _02597_ _03318_ _03812_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o31a_1
X_06107_ net734 _02763_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__and2_1
XFILLER_106_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505__157 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__inv_2
X_07087_ net578 _03743_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nor2_1
X_06038_ top0.CPU.register.registers\[265\] top0.CPU.register.registers\[297\] top0.CPU.register.registers\[329\]
+ top0.CPU.register.registers\[361\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02695_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07167__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout122 net123 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_93_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1109 net1115 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_2
Xfanout111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xfanout144 _04937_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
Xfanout155 net156 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
XANTENNA__06799__S1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout199 net201 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
Xfanout177 net178 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
XFILLER_47_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
Xfanout166 _04622_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
XANTENNA__08562__A1 _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _05234_ _05235_ _05237_ net241 vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a31o_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07989_ net714 net497 net216 net546 net2299 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_2_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06100__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _05162_ _05169_ _05175_ net142 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__and4b_1
XANTENNA__06325__B1 _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ clknet_leaf_91_clk _02305_ net1085 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08726__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297__949 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__inv_2
X_11621_ net1313 _01260_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06971__S1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11041__693 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__inv_2
XANTENNA__08093__A3 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ net1244 _01191_ net1030 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10276__B _05162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12772__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11483_ clknet_leaf_81_clk _01125_ net1109 vssd1 vssd1 vccd1 vccd1 top0.display.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_07_1180 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] team_07_1180/LO sky130_fd_sc_hd__conb_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07866__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1191 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] team_07_1191/LO sky130_fd_sc_hd__conb_1
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06487__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ net1796 _01743_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[597\]
+ sky130_fd_sc_hd__dfrtp_1
X_10296_ net3058 net118 net111 _05607_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22o_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12035_ net1727 _01674_ net1033 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[528\]
+ sky130_fd_sc_hd__dfrtp_1
X_10364__16 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__inv_2
XANTENNA__09145__X _04842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09305__B _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06411__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946__598 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ net1511 _01458_ net1070 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[312\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05848__X _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ _03621_ _03659_ _03661_ _03665_ _03076_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a311oi_4
X_10799__451 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__inv_2
XANTENNA__07044__A1 _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07495__B _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__S0 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08792__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08961_ _04655_ net275 net262 net2762 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__a22o_1
X_08892_ top0.CPU.register.registers\[240\] net571 net557 vssd1 vssd1 vccd1 vccd1
+ _04766_ sky130_fd_sc_hd__o21a_1
X_07912_ net633 _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__and2_1
X_07843_ top0.CPU.intMem_out\[28\] net627 _04496_ net642 vssd1 vssd1 vccd1 vccd1 _04497_
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout189_A _04592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _04426_ _04427_ _04429_ _04430_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__or4_1
XFILLER_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_27_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06650__S0 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09513_ top0.MMIO.WBData_i\[27\] top0.MMIO.WBData_i\[6\] top0.MMIO.WBData_i\[2\]
+ _02356_ net140 vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a41o_1
X_06725_ _03380_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nand2b_1
XFILLER_37_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout356_A _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ top0.MMIO.WBData_i\[15\] _04933_ net143 net139 _05039_ vssd1 vssd1 vccd1
+ vccd1 _05040_ sky130_fd_sc_hd__o2111a_1
X_06656_ top0.CPU.register.registers\[386\] top0.CPU.register.registers\[418\] top0.CPU.register.registers\[450\]
+ top0.CPU.register.registers\[482\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03313_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ net2288 _04541_ net606 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__mux2_1
X_06587_ _03223_ _03243_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__or2_1
X_11025__677 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__inv_2
XANTENNA_fanout523_A _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08326_ net3068 net409 net388 _04505_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08480__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08257_ net152 net670 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_95_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ net493 net159 net614 net425 net2259 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a32o_1
X_07208_ _03861_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06469__S0 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07139_ _03792_ _03795_ net347 vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08232__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05918__B _02574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _02924_ net551 vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_7_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ top0.display.delayctr\[10\] _05554_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__or2_1
X_10592__244 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__inv_2
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07338__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__B _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06641__S0 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12767__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10633__285 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__inv_2
XFILLER_28_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ clknet_leaf_71_clk _02288_ net1122 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ clknet_leaf_82_clk _02219_ net1109 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10409__61 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__inv_2
X_11604_ net1296 _01243_ net959 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08471__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07274__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11535_ net1227 _01174_ net1001 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ clknet_leaf_67_clk _01114_ net1119 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.rs2\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09015__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11397_ clknet_leaf_59_clk _01045_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08204__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10348_ net2255 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08774__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10279_ net2987 net118 net112 _05661_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a22o_1
X_12018_ net1710 _01657_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[511\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09035__B net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06632__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08829__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06510_ top0.CPU.register.registers\[403\] top0.CPU.register.registers\[435\] top0.CPU.register.registers\[467\]
+ top0.CPU.register.registers\[499\] net940 net906 vssd1 vssd1 vccd1 vccd1 _03167_
+ sky130_fd_sc_hd__mux4_1
X_07490_ _02810_ _02811_ _03221_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08874__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__C net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06441_ top0.CPU.register.registers\[790\] top0.CPU.register.registers\[822\] top0.CPU.register.registers\[854\]
+ top0.CPU.register.registers\[886\] net923 net888 vssd1 vssd1 vccd1 vccd1 _03098_
+ sky130_fd_sc_hd__mux4_1
XFILLER_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ _04717_ net281 net250 net2308 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__a22o_1
X_06372_ top0.CPU.register.registers\[926\] top0.CPU.register.registers\[958\] top0.CPU.register.registers\[990\]
+ top0.CPU.register.registers\[1022\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03029_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08057__A3 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ net3156 _04492_ net432 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XANTENNA__08462__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ top0.CPU.register.registers\[96\] net568 net555 vssd1 vssd1 vccd1 vccd1 _04821_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07265__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08042_ net510 net196 net709 net438 net2811 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06681__Y _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold912 top0.CPU.register.registers\[517\] vssd1 vssd1 vccd1 vccd1 net3134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold901 top0.CPU.register.registers\[37\] vssd1 vssd1 vccd1 vccd1 net3123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 net66 vssd1 vssd1 vccd1 vccd1 net3145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 net59 vssd1 vssd1 vccd1 vccd1 net3167 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold934 top0.CPU.register.registers\[925\] vssd1 vssd1 vccd1 vccd1 net3156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 top0.CPU.register.registers\[272\] vssd1 vssd1 vccd1 vccd1 net3189 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _05450_ _05463_ _05479_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a31o_1
Xhold989 net83 vssd1 vssd1 vccd1 vccd1 net3211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 top0.CPU.register.registers\[92\] vssd1 vssd1 vccd1 vccd1 net3200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 top0.CPU.register.registers\[387\] vssd1 vssd1 vccd1 vccd1 net3178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06871__S0 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ top0.CPU.register.registers\[202\] net573 net559 vssd1 vssd1 vccd1 vccd1
+ _04780_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_90_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10576__228 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__inv_2
XANTENNA__09226__A top0.CPU.internalMem.pcOut\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05754__A top0.CPU.control.funct7\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06528__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _04511_ net552 _04758_ net282 net3162 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__a32o_1
X_07826_ net721 net512 net150 net548 net2483 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a32o_1
XANTENNA_hold1219_A top0.CPU.intMem_out\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10617__269 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__inv_2
XFILLER_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ net453 _04111_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ net454 _03247_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07688_ _03444_ _04321_ _03427_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout905_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ net3404 net598 net131 _05029_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__B1 _03356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06639_ _03294_ _03295_ net869 vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__mux2_1
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08048__A3 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ net2449 _04619_ net609 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XFILLER_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ net3005 net185 net416 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__mux2_1
X_09289_ _04944_ _04945_ _04946_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.loadCt_n\[1\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_119_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08024__B net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ net2836 net123 net115 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a21o_1
XANTENNA__11439__Q top0.CPU.intMem_out\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ _05596_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__nand2_1
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10064_ net3430 net664 net603 _05544_ _05145_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a221o_1
XANTENNA__05727__D1 top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09181__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11765__RESET_B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08692__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12636_ clknet_leaf_74_clk _02271_ net1125 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07103__B _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xnet1023_2 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ clknet_leaf_57_clk _02206_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12498_ net2190 _02137_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[991\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold208 top0.CPU.register.registers\[200\] vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_11518_ net1210 _01157_ net1007 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11449_ clknet_leaf_69_clk _01097_ net1118 vssd1 vssd1 vccd1 vccd1 top0.CPU.Op\[6\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold219 top0.CPU.register.registers\[978\] vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373__1025 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06853__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06990_ _03645_ _03646_ net869 vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05941_ _02579_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__nor2_1
X_08660_ net947 net699 _04734_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__nand3_1
XFILLER_94_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05872_ top0.CPU.register.registers\[139\] top0.CPU.register.registers\[171\] top0.CPU.register.registers\[203\]
+ top0.CPU.register.registers\[235\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02529_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06081__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ net477 _03814_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__nand2_1
X_08591_ _02398_ _02404_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__nor2_2
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08278__A3 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07542_ _03005_ _03054_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__or2_1
XANTENNA__08683__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07473_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961__613 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__inv_2
X_09212_ top0.CPU.intMemAddr\[26\] top0.CPU.intMemAddr\[25\] top0.CPU.intMemAddr\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__or3_1
X_06424_ _03079_ _03080_ net758 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
X_06355_ top0.CPU.register.registers\[670\] top0.CPU.register.registers\[702\] top0.CPU.register.registers\[734\]
+ top0.CPU.register.registers\[766\] net850 net815 vssd1 vssd1 vccd1 vccd1 _03012_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09143_ top0.CPU.register.registers\[64\] net568 net555 vssd1 vssd1 vccd1 vccd1 _04841_
+ sky130_fd_sc_hd__o21a_1
XFILLER_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10242__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11096__748 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__inv_2
XANTENNA__07789__A2 _03482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05749__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06286_ net584 _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__nand2_1
X_09074_ _04686_ net274 net256 net2507 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__a22o_1
Xhold720 top0.CPU.register.registers\[534\] vssd1 vssd1 vccd1 vccd1 net2942 sky130_fd_sc_hd__dlygate4sd3_1
X_08025_ net3195 net437 _04643_ net493 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a22o_1
X_11137__789 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__inv_2
Xhold742 top0.CPU.register.registers\[421\] vssd1 vssd1 vccd1 vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09655__S _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold764 top0.CPU.register.registers\[884\] vssd1 vssd1 vccd1 vccd1 net2986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 top0.CPU.register.registers\[305\] vssd1 vssd1 vccd1 vccd1 net2975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 top0.CPU.register.registers\[953\] vssd1 vssd1 vccd1 vccd1 net2953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 top0.CPU.register.registers\[358\] vssd1 vssd1 vccd1 vccd1 net3019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 top0.CPU.register.registers\[259\] vssd1 vssd1 vccd1 vccd1 net3008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 top0.CPU.register.registers\[437\] vssd1 vssd1 vccd1 vccd1 net2997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09976_ top0.CPU.internalMem.pcOut\[26\] _05455_ vssd1 vssd1 vccd1 vccd1 _05468_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06844__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout855_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ _04645_ net267 net263 net2859 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__a22o_1
X_08858_ net168 net3206 net356 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__mux2_1
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08910__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07809_ net530 _03403_ net528 net527 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ net176 net683 net318 net291 net2646 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a32o_1
XANTENNA__08269__A3 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07204__A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12421_ net2113 _02060_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[914\]
+ sky130_fd_sc_hd__dfrtp_1
X_10745__397 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__inv_2
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12352_ net2044 _01991_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[845\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net1975 _01922_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[776\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10598__250 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__inv_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06835__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05963__A1 top0.CPU.decoder.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ top0.display.delayctr\[18\] _05579_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05963__B2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ top0.display.delayctr\[0\] top0.display.delayctr\[1\] vssd1 vssd1 vccd1 vccd1
+ _05532_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07165__A0 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10639__291 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__inv_2
Xhold91 top0.CPU.register.registers\[1001\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 top0.CPU.register.registers\[871\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06063__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05810__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ net1690 _01637_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[491\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_34_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07468__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08680__A3 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ clknet_leaf_74_clk _02254_ net1127 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08417__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10224__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06140_ net777 _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__nor2_1
X_06071_ _02724_ _02725_ _02727_ _02726_ net784 net738 vssd1 vssd1 vccd1 vccd1 _02728_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_74_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ net236 _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_2
Xfanout529 _03425_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
Xfanout518 _03685_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_2
XANTENNA__05735__C net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09761_ top0.CPU.internalMem.pcOut\[9\] net650 _05266_ _05269_ vssd1 vssd1 vccd1
+ vccd1 _02186_ sky130_fd_sc_hd__o22a_1
XFILLER_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06973_ _03628_ _03629_ net870 vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__mux2_1
X_08712_ _04566_ net3204 net359 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__mux2_1
X_05924_ top0.CPU.register.registers\[512\] top0.CPU.register.registers\[544\] top0.CPU.register.registers\[576\]
+ top0.CPU.register.registers\[608\] net836 net801 vssd1 vssd1 vccd1 vccd1 _02581_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09504__A top0.MMIO.WBData_i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ top0.CPU.internalMem.pcOut\[3\] net768 top0.CPU.internalMem.pcOut\[4\] vssd1
+ vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09696__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06054__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ net200 net707 net319 net303 net2268 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a32o_1
X_05855_ net579 _02505_ _02511_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__or3_1
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout171_A _04611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05751__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08574_ net2979 net221 net334 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
X_05786_ top0.CPU.register.registers\[407\] top0.CPU.register.registers\[439\] top0.CPU.register.registers\[471\]
+ top0.CPU.register.registers\[503\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02443_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout269_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07525_ _02650_ _03279_ _04124_ _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08656__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
X_07456_ net517 _04111_ _04112_ net450 vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a211o_1
XANTENNA__08408__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _04017_ _04018_ _04031_ _04043_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__o211ai_4
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06407_ top0.CPU.register.registers\[540\] top0.CPU.register.registers\[572\] top0.CPU.register.registers\[604\]
+ top0.CPU.register.registers\[636\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03064_
+ sky130_fd_sc_hd__mux4_1
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09081__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ top0.CPU.register.registers\[75\] net570 net557 vssd1 vssd1 vccd1 vccd1 _04835_
+ sky130_fd_sc_hd__o21a_1
X_06338_ _02993_ _02994_ net732 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_136_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__A2 _05006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06269_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09057_ top0.CPU.register.registers\[121\] net564 vssd1 vssd1 vccd1 vccd1 _04812_
+ sky130_fd_sc_hd__or2_1
X_08008_ top0.CPU.intMem_out\[0\] net629 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__and2_1
XANTENNA__09385__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 top0.CPU.register.registers\[479\] vssd1 vssd1 vccd1 vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold550 top0.CPU.register.registers\[651\] vssd1 vssd1 vccd1 vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 top0.CPU.register.registers\[313\] vssd1 vssd1 vccd1 vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06817__S0 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold594 top0.CPU.register.registers\[916\] vssd1 vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 top0.CPU.register.registers\[430\] vssd1 vssd1 vccd1 vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ _05437_ _05440_ _05439_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06293__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07147__B1 _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921_ net1613 _01560_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[414\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08895__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ net1544 _01491_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[345\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08647__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11452__Q top0.CPU.decoder.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__Q top0.CPU.internalMem.pcOut\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372__1024 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__inv_2
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12775__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
X_11783_ net1475 _01422_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08972__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09072__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ net2096 _02043_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08414__A3 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12335_ net2027 _01974_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12266_ net1958 _01905_ net984 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[759\]
+ sky130_fd_sc_hd__dfrtp_1
X_12197_ net1889 _01836_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[690\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__07386__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__06284__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06036__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06159__S net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__A2 _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_07310_ _03385_ _03407_ _03409_ _03559_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__or4_2
XANTENNA__08638__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08882__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07779__A _02578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ net2939 net224 net414 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
XANTENNA__07498__B net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07241_ _02983_ _03073_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__xnor2_1
X_07172_ _03022_ _03037_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09063__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09602__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06123_ _02778_ _02779_ net786 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XANTENNA__08810__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06054_ top0.CPU.register.registers\[136\] top0.CPU.register.registers\[168\] top0.CPU.register.registers\[200\]
+ top0.CPU.register.registers\[232\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02711_
+ sky130_fd_sc_hd__mux4_1
Xfanout304 _04740_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07377__A0 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 net328 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09813_ _02773_ _04573_ net586 vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__mux2_1
XFILLER_59_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
Xfanout348 _02576_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_2
Xfanout337 _03775_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06275__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ top0.CPU.internalMem.pcOut\[8\] top0.CPU.internalMem.pcOut\[7\] _05228_ vssd1
+ vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_87_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07129__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06956_ top0.CPU.register.registers\[24\] top0.CPU.register.registers\[56\] top0.CPU.register.registers\[88\]
+ top0.CPU.register.registers\[120\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03613_
+ sky130_fd_sc_hd__mux4_1
X_09675_ top0.CPU.internalMem.pcOut\[3\] _05188_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nand2_1
X_06887_ top0.CPU.register.registers\[520\] top0.CPU.register.registers\[552\] top0.CPU.register.registers\[584\]
+ top0.CPU.register.registers\[616\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03544_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05907_ top0.CPU.register.registers\[258\] top0.CPU.register.registers\[290\] top0.CPU.register.registers\[322\]
+ top0.CPU.register.registers\[354\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02564_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08877__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05838_ net867 _02474_ _02472_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a21o_1
XFILLER_55_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08626_ net717 net154 net316 net330 net2902 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a32o_1
XANTENNA__05786__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout720_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ net3048 _04481_ net336 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout818_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
X_05769_ _02424_ _02425_ _02372_ _02374_ _02407_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__o2111a_1
X_08488_ net151 net686 net404 net367 net2295 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__a32o_1
X_07508_ _04021_ _04049_ _04163_ _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_25_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ _02684_ _03404_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09624__A_N _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09054__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09109_ top0.CPU.register.registers\[85\] net569 vssd1 vssd1 vccd1 vccd1 _04828_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08801__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152__804 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__inv_2
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ net1812 _01759_ net1029 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[613\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold380 top0.CPU.register.registers\[100\] vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_12051_ net1743 _01690_ net1065 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[544\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07907__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 top0.CPU.register.registers\[43\] vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08032__B net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__Q top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout871 net873 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
Xfanout893 net895 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_4
Xfanout882 net885 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_51_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08868__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11904_ net1596 _01543_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[397\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1091 top0.CPU.register.registers\[82\] vssd1 vssd1 vccd1 vccd1 net3313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1080 top0.CPU.register.registers\[33\] vssd1 vssd1 vccd1 vccd1 net3302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08332__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11835_ net1527 _01474_ net1010 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[328\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_25_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ net1458 _01405_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[259\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07843__A1 top0.CPU.intMem_out\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760__412 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__inv_2
X_11697_ net1389 _01336_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[190\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08399__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801__453 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__inv_2
XANTENNA__05847__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12318_ net2010 _01957_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[811\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06442__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12249_ net1941 _01888_ net980 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06257__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06582__A1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ _02733_ _02770_ _02750_ net540 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__o211ai_1
X_07790_ net517 _03862_ _03865_ _03850_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_69_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06741_ _03396_ _03397_ net757 vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08859__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09460_ net131 net133 _05048_ net598 net3427 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__o32a_1
XANTENNA__08323__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08411_ net218 net695 net399 net379 net2321 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__a32o_1
XANTENNA__06334__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06672_ net869 _03326_ net862 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_82_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09391_ _02343_ _03709_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_16_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_08342_ net718 net186 net398 net411 net2403 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a32o_1
X_08273_ net512 net194 net675 net419 net2393 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08626__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ _03879_ _03880_ net346 vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__mux2_1
XANTENNA__08832__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09036__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _02579_ _02597_ _03338_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o21ai_1
X_06106_ top0.CPU.register.registers\[268\] top0.CPU.register.registers\[300\] top0.CPU.register.registers\[332\]
+ top0.CPU.register.registers\[364\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05757__A _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ _02428_ _03712_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__or2_4
X_10544__196 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__inv_2
X_06037_ top0.CPU.register.registers\[393\] top0.CPU.register.registers\[425\] top0.CPU.register.registers\[457\]
+ top0.CPU.register.registers\[489\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02694_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07972__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout112 net114 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
X_11371__1023 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__inv_2
Xfanout134 _05040_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_2
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
XFILLER_99_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout156 _04635_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
Xfanout167 _04615_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
X_07988_ top0.CPU.internalMem.pcOut\[4\] net640 net635 _04617_ vssd1 vssd1 vccd1 vccd1
+ _04618_ sky130_fd_sc_hd__o211a_2
Xfanout189 _04592_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout178 _04607_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _05234_ _05235_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06939_ top0.CPU.register.registers\[409\] top0.CPU.register.registers\[441\] top0.CPU.register.registers\[473\]
+ top0.CPU.register.registers\[505\] net910 net876 vssd1 vssd1 vccd1 vccd1 _03596_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _02748_ _05158_ _05166_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__and4_1
XFILLER_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06325__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ top0.display.counter\[3\] top0.display.counter\[2\] _04960_ _05124_ _05130_
+ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a41o_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08609_ net2948 net329 net308 _04562_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ net1312 _01259_ net985 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_11551_ net1243 _01190_ net1095 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06089__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08617__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09027__A0 _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11482_ clknet_leaf_78_clk top0.CPU.addrControl net1114 vssd1 vssd1 vccd1 vccd1 top0.CPU.muxAddr.prev_control
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05931__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1170 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] team_07_1170/LO sky130_fd_sc_hd__conb_1
Xteam_07_1181 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] team_07_1181/LO sky130_fd_sc_hd__conb_1
XANTENNA__07053__A2 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1192 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] team_07_1192/LO sky130_fd_sc_hd__conb_1
XANTENNA__06487__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ net1795 _01742_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[596\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08250__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10295_ net3083 net119 net113 _05667_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a22o_1
X_12034_ net1726 _01673_ net1054 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[527\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09750__A1 top0.CPU.control.funct7\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08553__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06564__A1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05998__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 net692 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11280__932 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__inv_2
XANTENNA__06411__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11321__973 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ net1510 _01457_ net983 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[311\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08069__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487__139 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__inv_2
X_11749_ net1441 _01388_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05827__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09018__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__A1 top0.CPU.decoder.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08792__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__S1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ _04654_ net278 net260 net2814 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__a22o_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
X_07911_ top0.CPU.internalMem.pcOut\[18\] net642 _04553_ _04554_ vssd1 vssd1 vccd1
+ vccd1 _04555_ sky130_fd_sc_hd__a22o_2
X_08891_ _04562_ net552 _04765_ net284 net3267 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__a32o_1
XANTENNA__08544__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07842_ net561 _04494_ _04495_ net625 vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__o211a_1
XANTENNA__10177__A_N net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05989__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ top0.MMIO.WBData_i\[12\] top0.MMIO.WBData_i\[9\] top0.MMIO.WBData_i\[0\]
+ _02357_ net138 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a41o_1
X_07773_ net452 _04239_ _03843_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06650__S1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06724_ _03365_ net530 vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__nand2_1
X_09443_ _02517_ _05002_ _05004_ _05000_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__o211a_1
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout251_A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06655_ _03310_ _03311_ net757 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__mux2_1
X_09374_ net2371 _04546_ net607 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout349_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06586_ _03201_ _03203_ _03221_ _03225_ net533 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__o32a_1
X_08325_ net2877 net409 net392 _04499_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold1199_A top0.CPU.intMem_out\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06166__S0 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07967__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ net2752 net418 _04713_ net501 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08187_ net497 net161 net615 net425 net2587 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a32o_1
X_07207_ net474 _03772_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ _03793_ _03794_ net460 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__mux2_1
XANTENNA__11883__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06469__S1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ _03357_ _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10080_ net3400 net665 net603 _05556_ _05157_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08535__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07338__A3 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264__916 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__inv_2
XANTENNA__06546__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06641__S1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08299__A1 _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__12600__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305__957 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__inv_2
XFILLER_130_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ clknet_leaf_74_clk _02287_ net1125 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ net1295 _01242_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11460__Q top0.CPU.decoder.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158__810 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__inv_2
XANTENNA__06157__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12583_ clknet_leaf_82_clk _02218_ net1108 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05904__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06781__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11534_ net1226 _01173_ net990 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11465_ clknet_leaf_74_clk _01113_ net1123 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.rs2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424__76 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__inv_2
XANTENNA__09420__B1 _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11396_ clknet_leaf_57_clk _01044_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10872__524 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__inv_2
X_10347_ net2252 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06785__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10278_ net144 _05164_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__nand2_1
X_12017_ net1709 _01656_ net1043 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[510\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08526__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913__565 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__inv_2
XFILLER_120_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07117__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__B1 _04033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06632__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05860__A top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__A _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08829__A3 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09051__B net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06440_ top0.CPU.register.registers\[918\] top0.CPU.register.registers\[950\] top0.CPU.register.registers\[982\]
+ top0.CPU.register.registers\[1014\] net922 net888 vssd1 vssd1 vccd1 vccd1 _03097_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06167__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370__1022 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__inv_2
X_06371_ top0.CPU.register.registers\[798\] top0.CPU.register.registers\[830\] top0.CPU.register.registers\[862\]
+ top0.CPU.register.registers\[894\] net935 net901 vssd1 vssd1 vccd1 vccd1 _03028_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06148__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__B net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ net2898 _04487_ net430 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
X_09090_ net157 net614 net268 net255 net2388 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_32_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08041_ net505 net199 net707 net438 net2370 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a32o_1
XANTENNA__07670__C1 _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold913 top0.CPU.register.registers\[823\] vssd1 vssd1 vccd1 vccd1 net3135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold902 top0.CPU.register.registers\[814\] vssd1 vssd1 vccd1 vccd1 net3124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 top0.CPU.register.registers\[819\] vssd1 vssd1 vccd1 vccd1 net3168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 top0.CPU.register.registers\[402\] vssd1 vssd1 vccd1 vccd1 net3146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold935 top0.CPU.register.registers\[283\] vssd1 vssd1 vccd1 vccd1 net3157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 top0.CPU.intMemAddr\[5\] vssd1 vssd1 vccd1 vccd1 net3190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09992_ top0.CPU.internalMem.pcOut\[27\] _05472_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05482_ sky130_fd_sc_hd__o21a_1
Xhold957 top0.CPU.register.registers\[412\] vssd1 vssd1 vccd1 vccd1 net3179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold979 top0.CPU.register.registers\[408\] vssd1 vssd1 vccd1 vccd1 net3201 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08943_ net187 net706 net276 net265 net2503 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__a32o_1
XANTENNA__06871__S1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout299_A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05754__B top0.CPU.control.funct7\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08517__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06528__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ top0.CPU.register.registers\[250\] net564 vssd1 vssd1 vccd1 vccd1 _04758_
+ sky130_fd_sc_hd__or2_1
X_07825_ net634 _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__and2_1
XFILLER_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08557__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _03131_ _03154_ _03914_ _03715_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a31o_1
XFILLER_65_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06707_ _03361_ _03362_ _03302_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ top0.MMIO.WBData_i\[9\] net145 _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout633_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07687_ _03966_ _03989_ _04319_ _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__or4_1
XANTENNA__06585__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06387__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__A1 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06638_ top0.CPU.register.registers\[387\] top0.CPU.register.registers\[419\] top0.CPU.register.registers\[451\]
+ top0.CPU.register.registers\[483\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03295_
+ sky130_fd_sc_hd__mux4_1
X_09357_ net2569 _04623_ net611 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
X_06569_ top0.CPU.register.registers\[656\] top0.CPU.register.registers\[688\] top0.CPU.register.registers\[720\]
+ top0.CPU.register.registers\[752\] net930 net896 vssd1 vssd1 vccd1 vccd1 _03226_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ top0.CPU.internalMem.loadCt\[0\] top0.CPU.internalMem.loadCt\[1\] vssd1 vssd1
+ vccd1 vccd1 _04946_ sky130_fd_sc_hd__nand2_1
XANTENNA__06805__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ net2746 net189 net415 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
XANTENNA__07256__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08239_ net950 net952 net954 vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nor3b_2
XFILLER_121_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07984__X _04615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856__508 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__inv_2
XANTENNA__08205__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10201_ _05011_ net129 net122 net3338 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XANTENNA__09953__A1 top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ top0.display.delayctr\[21\] _05591_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__nand2_1
X_10600__252 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__inv_2
XANTENNA__08321__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08508__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06112__Y _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10063_ _05542_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__nand2_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__Q top0.CPU.control.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09181__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05680__A top0.CPU.Op\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06378__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06495__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12635_ clknet_leaf_74_clk _02270_ net1125 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08444__A1 _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ clknet_leaf_56_clk _02205_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06715__S net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ net1209 _01156_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08995__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ net2189 _02136_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[990\]
+ sky130_fd_sc_hd__dfrtp_1
X_11448_ clknet_leaf_70_clk _01096_ net1117 vssd1 vssd1 vccd1 vccd1 top0.CPU.Op\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06016__A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 top0.CPU.register.registers\[964\] vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08747__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ clknet_leaf_79_clk _01027_ net1111 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07955__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05855__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06450__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06853__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06303__X _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_72_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12593__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09046__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05940_ net584 _02587_ _02595_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__and3_2
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__09172__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05871_ top0.CPU.register.registers\[395\] top0.CPU.register.registers\[427\] top0.CPU.register.registers\[459\]
+ top0.CPU.register.registers\[491\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02528_
+ sky130_fd_sc_hd__mux4_1
X_08590_ net947 net722 _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__nand3_1
XANTENNA__05861__Y _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08380__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07610_ net490 _04010_ _04265_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__o21ai_1
X_07541_ _03022_ _03037_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07472_ _03704_ _03829_ _03883_ _03898_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_17_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ _04524_ _04578_ _04589_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__or4_1
XANTENNA__07891__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06423_ top0.CPU.register.registers\[535\] top0.CPU.register.registers\[567\] top0.CPU.register.registers\[599\]
+ top0.CPU.register.registers\[631\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03080_
+ sky130_fd_sc_hd__mux4_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06354_ top0.CPU.register.registers\[798\] top0.CPU.register.registers\[830\] top0.CPU.register.registers\[862\]
+ top0.CPU.register.registers\[894\] net853 net818 vssd1 vssd1 vccd1 vccd1 _03011_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08435__A1 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ net157 net679 net268 net251 net2701 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a32o_1
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ net196 net622 net278 net257 net2385 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__a32o_1
XANTENNA__12573__D net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08986__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05749__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06285_ net741 _02941_ _02936_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a21oi_4
Xhold710 top0.CPU.register.registers\[542\] vssd1 vssd1 vccd1 vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08840__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold721 top0.CPU.register.registers\[949\] vssd1 vssd1 vccd1 vccd1 net2943 sky130_fd_sc_hd__dlygate4sd3_1
X_08024_ _04516_ net704 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__and2_1
Xhold743 top0.CPU.register.registers\[563\] vssd1 vssd1 vccd1 vccd1 net2965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08738__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold754 top0.CPU.register.registers\[505\] vssd1 vssd1 vccd1 vccd1 net2976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 top0.CPU.register.registers\[898\] vssd1 vssd1 vccd1 vccd1 net2954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 net74 vssd1 vssd1 vccd1 vccd1 net2987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 top0.CPU.register.registers\[1020\] vssd1 vssd1 vccd1 vccd1 net3009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 top0.CPU.register.registers\[536\] vssd1 vssd1 vccd1 vccd1 net2998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ top0.CPU.internalMem.pcOut\[26\] _05455_ vssd1 vssd1 vccd1 vccd1 _05467_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06844__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 top0.CPU.register.registers\[791\] vssd1 vssd1 vccd1 vccd1 net3020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__Y _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ _04644_ net275 net264 net2534 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09671__S net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout750_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ net172 net2937 net353 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__mux2_1
XANTENNA__09163__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ net531 _03317_ _03338_ _03356_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and4_1
XFILLER_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08788_ net217 net683 net318 net291 net2324 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ _03847_ _04029_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__nand2_1
XANTENNA__07021__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09871__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__X _04611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09409_ top0.MMIO.WBData_i\[3\] _04933_ net143 top0.MISOtoMMIO\[3\] _05014_ vssd1
+ vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_101_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12420_ net2112 _02059_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06535__S net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11120__772 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__inv_2
XANTENNA__08977__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ net2043 _01990_ net1094 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[844\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06532__S0 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12282_ net1974 _01921_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[775\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06835__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ top0.display.delayctr\[18\] _05579_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__or2_1
XFILLER_0_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10046_ top0.display.delayctr\[0\] net664 _05132_ _05531_ vssd1 vssd1 vccd1 vccd1
+ _02209_ sky130_fd_sc_hd__a211o_1
Xhold92 top0.CPU.register.registers\[968\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 top0.CPU.register.registers\[587\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06599__S0 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 top0.CPU.register.registers\[162\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__A1 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984__636 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__inv_2
X_11997_ net1689 _01636_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05751__A_N net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12618_ clknet_leaf_74_clk _02253_ net1125 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06445__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12549_ clknet_leaf_60_clk _02188_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_06070_ top0.CPU.register.registers\[10\] top0.CPU.register.registers\[42\] top0.CPU.register.registers\[74\]
+ top0.CPU.register.registers\[106\] net848 net813 vssd1 vssd1 vccd1 vccd1 _02727_
+ sky130_fd_sc_hd__mux4_1
X_10878__530 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__inv_2
XANTENNA_1 _02471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout508 net515 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
Xfanout519 _03685_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06180__S net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919__571 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__inv_2
X_09760_ net241 _05267_ _05268_ _02368_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a31o_1
X_06972_ top0.CPU.register.registers\[923\] top0.CPU.register.registers\[955\] top0.CPU.register.registers\[987\]
+ top0.CPU.register.registers\[1019\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03629_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05735__D net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _05201_ _05203_ net237 vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05923_ top0.CPU.register.registers\[640\] top0.CPU.register.registers\[672\] top0.CPU.register.registers\[704\]
+ top0.CPU.register.registers\[736\] net835 net800 vssd1 vssd1 vccd1 vccd1 _02580_
+ sky130_fd_sc_hd__mux4_1
X_08711_ net222 net3109 net357 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__mux2_1
Xfanout1090 net1092 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07156__A1 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08642_ _04650_ net308 net301 net2819 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a22o_1
X_05854_ net743 _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__and2_2
XANTENNA__09504__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08573_ net3184 _04571_ net335 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
X_11063__715 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__inv_2
XANTENNA__09223__C top0.CPU.internalMem.pcOut\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout164_A _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05785_ top0.CPU.register.registers\[23\] top0.CPU.register.registers\[55\] top0.CPU.register.registers\[87\]
+ top0.CPU.register.registers\[119\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02442_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08105__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ net454 net530 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__nand2_1
XANTENNA__08835__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07864__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ net485 _03865_ _04110_ _03759_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104__756 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__inv_2
XANTENNA__06863__B _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ top0.CPU.register.registers\[668\] top0.CPU.register.registers\[700\] top0.CPU.register.registers\[732\]
+ top0.CPU.register.registers\[764\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout429_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06193__A1_N net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07386_ _04033_ _04042_ net454 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a21o_1
XFILLER_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ net190 net688 _04834_ net254 net3265 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a32o_1
XANTENNA__08959__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__C1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06337_ top0.CPU.register.registers\[29\] top0.CPU.register.registers\[61\] top0.CPU.register.registers\[93\]
+ top0.CPU.register.registers\[125\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02994_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08570__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07092__B1 _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06268_ _02910_ _02924_ net584 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_2
X_09056_ _04677_ net267 net255 net2984 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__a22o_1
XANTENNA__09908__A1 top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ net563 _04631_ _04588_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout798_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold551 top0.CPU.register.registers\[873\] vssd1 vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
X_06199_ top0.CPU.register.registers\[532\] top0.CPU.register.registers\[564\] top0.CPU.register.registers\[596\]
+ top0.CPU.register.registers\[628\] net845 net810 vssd1 vssd1 vccd1 vccd1 _02856_
+ sky130_fd_sc_hd__mux4_1
Xhold562 top0.CPU.register.registers\[294\] vssd1 vssd1 vccd1 vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 top0.CPU.register.registers\[189\] vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06817__S1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 top0.CPU.register.registers\[658\] vssd1 vssd1 vccd1 vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__A3 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold584 top0.CPU.register.registers\[951\] vssd1 vssd1 vccd1 vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold595 top0.CPU.register.registers\[597\] vssd1 vssd1 vccd1 vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
X_09958_ _05449_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__nand2_1
XANTENNA__09136__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ net714 net214 net271 net282 net2555 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__a32o_1
X_10671__323 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__inv_2
X_09889_ top0.CPU.internalMem.pcOut\[20\] _05385_ vssd1 vssd1 vccd1 vccd1 _05387_
+ sky130_fd_sc_hd__xor2_2
XANTENNA__08344__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__10151__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ net1612 _01559_ net1079 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[413\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712__364 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__inv_2
XFILLER_45_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ net1543 _01490_ net1067 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[344\]
+ sky130_fd_sc_hd__dfrtp_1
X_11782_ net1474 _01421_ net1129 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[275\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11397__RESET_B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06265__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ net2095 _02042_ net1060 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__S0 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12334_ net2026 _01973_ net1058 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05957__X _02614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12265_ net1957 _01904_ net1073 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[758\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__08178__A3 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07386__A1 _04033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net1888 _01835_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[689\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__09127__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__A _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08335__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ top0.CPU.internalMem.pcOut\[30\] _05504_ vssd1 vssd1 vccd1 vccd1 _05517_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06992__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09340__A _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08102__A3 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__B _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07240_ _02983_ net538 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__and2_1
XFILLER_20_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07171_ _03022_ net539 vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__nand2b_1
X_06122_ top0.CPU.register.registers\[910\] top0.CPU.register.registers\[942\] top0.CPU.register.registers\[974\]
+ top0.CPU.register.registers\[1006\] net836 net801 vssd1 vssd1 vccd1 vccd1 _02779_
+ sky130_fd_sc_hd__mux4_1
XFILLER_117_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07613__A2 _03317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06053_ _02708_ _02709_ net784 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XFILLER_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08169__A3 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10385__37 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__inv_2
XANTENNA__07377__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_4
X_09812_ top0.CPU.internalMem.pcOut\[14\] net648 vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__nor2_1
XANTENNA__09771__C1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655__307 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__inv_2
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_4
Xfanout338 _03775_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09118__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09743_ _05246_ _05251_ net237 vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_87_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08326__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ top0.CPU.register.registers\[152\] top0.CPU.register.registers\[184\] top0.CPU.register.registers\[216\]
+ top0.CPU.register.registers\[248\] net924 net890 vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__mux4_1
X_09674_ top0.CPU.internalMem.pcOut\[3\] _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__nor2_1
X_06886_ top0.CPU.register.registers\[648\] top0.CPU.register.registers\[680\] top0.CPU.register.registers\[712\]
+ top0.CPU.register.registers\[744\] net928 net894 vssd1 vssd1 vccd1 vccd1 _03543_
+ sky130_fd_sc_hd__mux4_1
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05906_ _02559_ _02560_ _02561_ _02562_ net724 net735 vssd1 vssd1 vccd1 vccd1 _02563_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__08341__A3 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05837_ net581 _02493_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__nand2_1
X_08625_ net713 net158 net306 net329 net2421 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a32o_1
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ _02393_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor2_4
XANTENNA__05786__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05768_ net944 net943 net942 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__and3b_1
X_10549__201 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__inv_2
X_07507_ _03973_ _04004_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__nor2_1
XANTENNA__08565__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05699_ top0.MMIO.WBData_i\[17\] vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__inv_2
X_08487_ net948 net545 _04688_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__or3_4
XANTENNA__06735__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06085__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07438_ net483 _04091_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07369_ net480 net474 _03772_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__or3b_1
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07065__A0 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ _04698_ net273 net252 net2614 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__a22o_1
XFILLER_136_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191__843 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_98_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09039_ net171 net3007 net349 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__mux2_1
X_12050_ net1742 _01689_ net1053 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[543\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold381 top0.CPU.register.registers\[195\] vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 top0.CPU.register.registers\[673\] vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
X_11232__884 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__inv_2
XFILLER_78_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold392 top0.CPU.register.registers\[86\] vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout861 top0.CPU.decoder.instruction\[19\] vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_129_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout850 net853 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_4
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_2
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
Xfanout883 net885 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1092 top0.CPU.register.registers\[396\] vssd1 vssd1 vccd1 vccd1 net3314 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ net1595 _01542_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11463__Q top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12559__Q top0.CPU.internalMem.pcOut\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1070 top0.CPU.register.registers\[68\] vssd1 vssd1 vccd1 vccd1 net3292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 top0.CPU.register.registers\[758\] vssd1 vssd1 vccd1 vccd1 net3303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11834_ net1526 _01473_ net1005 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ net1457 _01404_ net982 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[258\]
+ sky130_fd_sc_hd__dfrtp_1
X_11696_ net1388 _01335_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[189\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10840__492 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__inv_2
XANTENNA__09596__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ net2009 _01956_ net1027 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[810\]
+ sky130_fd_sc_hd__dfrtp_1
X_12248_ net1940 _01887_ net1028 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[741\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08223__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07359__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ net1871 _01818_ net1057 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[672\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355__7 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__inv_2
XFILLER_49_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06740_ top0.CPU.register.registers\[6\] top0.CPU.register.registers\[38\] top0.CPU.register.registers\[70\]
+ top0.CPU.register.registers\[102\] net916 net881 vssd1 vssd1 vccd1 vccd1 _03397_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06671_ net756 _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__or2_1
X_08410_ _04600_ net696 net401 net379 net2285 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a32o_1
XANTENNA__07531__B2 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09390_ _02342_ _02424_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__nand2_1
X_08341_ net722 net192 net407 net412 net2381 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a32o_1
X_08272_ net3124 net418 _04719_ net502 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06717__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07223_ _03722_ _03732_ net460 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__mux2_1
XFILLER_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175__827 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__inv_2
XANTENNA__05877__A1_N _02532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ net455 _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nand2_1
X_06105_ top0.CPU.register.registers\[396\] top0.CPU.register.registers\[428\] top0.CPU.register.registers\[460\]
+ top0.CPU.register.registers\[492\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02762_
+ sky130_fd_sc_hd__mux4_1
X_07085_ _02428_ _03712_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nor2_2
XANTENNA__08795__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06036_ top0.CPU.register.registers\[9\] top0.CPU.register.registers\[41\] top0.CPU.register.registers\[73\]
+ top0.CPU.register.registers\[105\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02693_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1036_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216__868 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_2
XANTENNA__08547__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout135 _05037_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
Xfanout124 _05641_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
X_11069__721 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__inv_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
Xfanout168 _04615_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlymetal6s2s_1
X_07987_ top0.CPU.intMem_out\[4\] net629 _04476_ _04616_ net643 vssd1 vssd1 vccd1
+ vccd1 _04617_ sky130_fd_sc_hd__a221o_1
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_2
X_09726_ _05222_ _05226_ _05220_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06938_ _03593_ _03594_ net756 vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06869_ top0.CPU.register.registers\[777\] top0.CPU.register.registers\[809\] top0.CPU.register.registers\[841\]
+ top0.CPU.register.registers\[873\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03526_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09657_ _02715_ _05151_ _05156_ _02532_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout830_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06325__A2 _02978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06956__S0 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ net719 net202 net319 net331 net2506 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a32o_1
X_09588_ top0.display.state\[0\] _05129_ net666 top0.display.counter\[4\] vssd1 vssd1
+ vccd1 vccd1 _05130_ sky130_fd_sc_hd__o211a_1
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08295__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _04719_ net394 net362 net3104 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a22o_1
X_10783__435 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__inv_2
XANTENNA__06089__A1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ net1242 _01189_ net1007 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05836__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ clknet_leaf_84_clk _01124_ net1107 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824__476 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__inv_2
XANTENNA__05931__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1160 vssd1 vssd1 vccd1 vccd1 team_07_1160/HI gpio_out[26] sky130_fd_sc_hd__conb_1
Xteam_07_1171 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] team_07_1171/LO sky130_fd_sc_hd__conb_1
Xteam_07_1182 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] team_07_1182/LO sky130_fd_sc_hd__conb_1
XANTENNA__08786__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08250__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1193 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] team_07_1193/LO sky130_fd_sc_hd__conb_1
X_12102_ net1794 _01741_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[595\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08043__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _02446_ net551 net144 vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_53_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12033_ net1725 _01672_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[526\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718__370 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__inv_2
XANTENNA__05683__A top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A3 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05998__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_4
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_29_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08710__A0 _04555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06947__S0 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11817_ net1509 _01456_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08069__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05827__A1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11748_ net1440 _01387_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[241\]
+ sky130_fd_sc_hd__dfrtp_1
X_11679_ net1371 _01318_ net1096 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[172\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06961__B net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06453__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ top0.CPU.intMem_out\[18\] net625 _02495_ _02386_ net638 vssd1 vssd1 vccd1
+ vccd1 _04554_ sky130_fd_sc_hd__o221a_1
XFILLER_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08890_ top0.CPU.register.registers\[241\] net567 vssd1 vssd1 vccd1 vccd1 _04765_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08544__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07841_ net591 _02981_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__nand2_1
XANTENNA__05989__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07752__A1 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _03760_ _04428_ _04424_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__o21ai_1
X_09511_ _05089_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__nor2_1
XFILLER_110_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06723_ _03365_ net530 vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__nor2_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470__122 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__inv_2
X_09442_ top0.MMIO.WBData_i\[16\] net145 net135 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__o21a_1
XFILLER_80_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06654_ top0.CPU.register.registers\[2\] top0.CPU.register.registers\[34\] top0.CPU.register.registers\[66\]
+ top0.CPU.register.registers\[98\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03311_
+ sky130_fd_sc_hd__mux4_1
X_10767__419 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ net2866 _04552_ net607 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__mux2_1
X_06585_ _03225_ net533 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout244_A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511__163 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__inv_2
X_08324_ net3130 net410 net397 _04493_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XANTENNA__06166__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05818__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08843__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08255_ _04522_ net671 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__and2_1
XFILLER_137_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06363__S net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ net453 _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nor2_1
X_08186_ net495 net165 net618 net425 net2626 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_95_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08768__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ _03221_ net534 net468 vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ net470 _03338_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06019_ top0.CPU.register.registers\[262\] top0.CPU.register.registers\[294\] top0.CPU.register.registers\[326\]
+ top0.CPU.register.registers\[358\] net833 net797 vssd1 vssd1 vccd1 vccd1 _02676_
+ sky130_fd_sc_hd__mux4_1
XFILLER_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08940__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ top0.CPU.internalMem.pcOut\[6\] _05219_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__or2_1
XANTENNA__06929__S0 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344__996 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__inv_2
X_12651_ clknet_leaf_71_clk _02286_ net1119 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09248__A1 _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ net1294 _01241_ net1052 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06157__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ clknet_leaf_83_clk _02217_ net1110 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08471__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ net1225 _01172_ net956 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11464_ clknet_leaf_70_clk _01112_ net1121 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.rs2\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05904__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238__890 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__inv_2
X_11395_ clknet_leaf_59_clk _01043_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07893__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ net2240 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10277_ net3233 net121 net114 _05660_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XANTENNA__05993__B1 _02649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ net1708 _01655_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[509\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11593__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09184__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10454__106 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__inv_2
XFILLER_66_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07117__B _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06370_ net867 _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__nor2_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06148__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06473__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06183__S net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08040_ net3352 net439 _04650_ net495 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
Xhold903 top0.CPU.register.registers\[268\] vssd1 vssd1 vccd1 vccd1 net3125 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A1 _02355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05875__X _02532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold925 top0.CPU.register.registers\[957\] vssd1 vssd1 vccd1 vccd1 net3147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 top0.CPU.register.registers\[854\] vssd1 vssd1 vccd1 vccd1 net3136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 top0.CPU.register.registers\[855\] vssd1 vssd1 vccd1 vccd1 net3158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ top0.CPU.internalMem.pcOut\[27\] _05472_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05481_ sky130_fd_sc_hd__a21o_1
Xhold958 top0.CPU.register.registers\[770\] vssd1 vssd1 vccd1 vccd1 net3180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 top0.CPU.register.registers\[890\] vssd1 vssd1 vccd1 vccd1 net3191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 top0.CPU.register.registers\[753\] vssd1 vssd1 vccd1 vccd1 net3169 sky130_fd_sc_hd__dlygate4sd3_1
X_08942_ net190 net710 net280 net266 net2474 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__a32o_1
X_11287__939 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09175__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08517__A3 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06084__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08922__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ net3102 net284 net269 _04505_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__a22o_1
X_11031__683 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__inv_2
X_07824_ _04479_ _04480_ top0.CPU.internalMem.pcOut\[31\] net639 vssd1 vssd1 vccd1
+ vccd1 _04481_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__08838__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07755_ _03131_ _03914_ _03154_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout361_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ net343 _04322_ _04330_ _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__a211o_1
XFILLER_65_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06706_ _03302_ _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__and2b_1
X_09425_ net143 net139 _05025_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__and3_2
XANTENNA__08150__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06637_ top0.CPU.register.registers\[259\] top0.CPU.register.registers\[291\] top0.CPU.register.registers\[323\]
+ top0.CPU.register.registers\[355\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03294_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06387__S1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__A2 _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08573__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ net2306 _04627_ net611 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
X_06568_ _02831_ _03199_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__xor2_1
X_09287_ top0.CPU.internalMem.loadCt\[0\] top0.CPU.internalMem.loadCt\[1\] vssd1 vssd1
+ vccd1 vccd1 _04945_ sky130_fd_sc_hd__or2_1
X_08307_ net2913 _04586_ net416 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XANTENNA__08989__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06499_ _02496_ _02833_ _02477_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__RESET_B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08238_ net495 net153 net682 net422 net2396 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_119_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout995_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ _04924_ _05638_ net122 net3335 net115 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a221o_1
X_08169_ net508 net203 net620 net427 net2319 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a32o_1
X_10895__547 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__inv_2
XANTENNA__08205__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08756__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ top0.display.delayctr\[21\] _05591_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__or2_1
X_10936__588 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__inv_2
XANTENNA__09166__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08508__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ top0.display.delayctr\[5\] _05539_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08913__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05822__S0 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05961__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10789__441 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__inv_2
XANTENNA__06268__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06378__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__Q top0.CPU.control.funct7\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08692__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ clknet_leaf_71_clk _02269_ net1122 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_61_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ clknet_leaf_56_clk _02204_ net1038 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_11516_ net1208 _01155_ net1019 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05889__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ net2188 _02135_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[989\]
+ sky130_fd_sc_hd__dfrtp_1
X_11447_ clknet_leaf_70_clk _01095_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.Op\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ clknet_leaf_73_clk top0.CPU.internalMem.loadCt_n\[2\] net1128 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.loadCt\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05855__B _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10329_ net2230 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__clkbuf_1
X_11015__667 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__inv_2
XANTENNA__08904__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09172__A3 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06066__S0 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05870_ top0.CPU.register.registers\[267\] top0.CPU.register.registers\[299\] top0.CPU.register.registers\[331\]
+ top0.CPU.register.registers\[363\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02527_
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05813__S0 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _02945_ _03656_ _04132_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_37_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07471_ _03701_ net519 vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_17_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ _04535_ _04563_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or2_1
X_06422_ top0.CPU.register.registers\[663\] top0.CPU.register.registers\[695\] top0.CPU.register.registers\[727\]
+ top0.CPU.register.registers\[759\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03079_
+ sky130_fd_sc_hd__mux4_1
X_06353_ top0.CPU.register.registers\[926\] top0.CPU.register.registers\[958\] top0.CPU.register.registers\[990\]
+ top0.CPU.register.registers\[1022\] net850 net815 vssd1 vssd1 vccd1 vccd1 _03010_
+ sky130_fd_sc_hd__mux4_1
X_09141_ net3249 net251 _04840_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ net200 net620 _04817_ net257 net3270 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__a32o_1
X_10582__234 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__inv_2
X_06284_ _02937_ _02938_ _02940_ _02939_ net782 net735 vssd1 vssd1 vccd1 vccd1 _02941_
+ sky130_fd_sc_hd__mux4_2
X_08023_ net3212 net437 _04642_ net491 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a22o_1
Xhold700 top0.CPU.register.registers\[392\] vssd1 vssd1 vccd1 vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 top0.CPU.register.registers\[648\] vssd1 vssd1 vccd1 vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 top0.CPU.register.registers\[645\] vssd1 vssd1 vccd1 vccd1 net2977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 top0.CPU.register.registers\[637\] vssd1 vssd1 vccd1 vccd1 net2944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 top0.CPU.register.registers\[668\] vssd1 vssd1 vccd1 vccd1 net2955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 top0.CPU.register.registers\[878\] vssd1 vssd1 vccd1 vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
X_10623__275 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__inv_2
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold766 top0.CPU.register.registers\[258\] vssd1 vssd1 vccd1 vccd1 net2988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 top0.CPU.register.registers\[541\] vssd1 vssd1 vccd1 vccd1 net2999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 top0.CPU.register.registers\[253\] vssd1 vssd1 vccd1 vccd1 net3010 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _05441_ _05463_ _05462_ _05450_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__o211ai_2
Xhold799 top0.CPU.register.registers\[245\] vssd1 vssd1 vccd1 vccd1 net3021 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout576_A _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _04643_ net268 net263 net2635 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold1224_A top0.MMIO.WBData_i\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08856_ net176 net3242 net355 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__mux2_1
XANTENNA__08568__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05804__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ net539 _03053_ net538 net521 vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__and4_1
XANTENNA__08910__A3 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ net180 net685 net322 net291 net2539 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout743_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05999_ top0.CPU.register.registers\[903\] top0.CPU.register.registers\[935\] top0.CPU.register.registers\[967\]
+ top0.CPU.register.registers\[999\] net831 net796 vssd1 vssd1 vccd1 vccd1 _02656_
+ sky130_fd_sc_hd__mux4_1
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07738_ _02925_ _03600_ net341 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a21o_1
XANTENNA__08123__A1 _04561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__Y _03540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ net441 _04156_ net340 vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout910_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ net3386 _04949_ _05017_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_101_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ _02338_ net629 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_134_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ net2042 _01989_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06532__S1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ net1973 _01920_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06296__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _02493_ net550 net141 vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09139__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__Q top0.CPU.control.rs2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10045_ top0.display.delayctr\[0\] net600 vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__nor2_1
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05691__A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 top0.CPU.register.registers\[624\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06599__S1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 top0.CPU.register.registers\[422\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 top0.CPU.register.registers\[354\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 top0.CPU.register.registers\[485\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06912__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ net1688 _01635_ net1021 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[489\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10102__A _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__A1 _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08665__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_14_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10566__218 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__inv_2
X_12617_ clknet_leaf_74_clk _02252_ net1127 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08417__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ clknet_leaf_60_clk _02187_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10224__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607__259 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__inv_2
X_12479_ net2171 _02118_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[972\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_2 _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout509 net511 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
XANTENNA__08050__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06971_ top0.CPU.register.registers\[795\] top0.CPU.register.registers\[827\] top0.CPU.register.registers\[859\]
+ top0.CPU.register.registers\[891\] net920 net886 vssd1 vssd1 vccd1 vccd1 _03628_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06039__S0 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ _05201_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__and2_1
X_08710_ _04555_ net3146 net359 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
X_05922_ net857 _02451_ _02516_ top0.CPU.decoder.instruction\[7\] vssd1 vssd1 vccd1
+ vccd1 _02579_ sky130_fd_sc_hd__a22o_4
XFILLER_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05853_ _02506_ _02507_ _02508_ _02509_ net729 net779 vssd1 vssd1 vccd1 vccd1 _02510_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09550__A0 top0.CPU.control.funct7\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_2
X_08641_ net202 net707 net319 net303 net2531 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a32o_1
XFILLER_67_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1080 net1083 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07156__A2 _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ net2832 _04566_ net335 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__mux2_1
X_05784_ top0.CPU.register.registers\[151\] top0.CPU.register.registers\[183\] top0.CPU.register.registers\[215\]
+ top0.CPU.register.registers\[247\] net825 net790 vssd1 vssd1 vccd1 vccd1 _02441_
+ sky130_fd_sc_hd__mux4_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08105__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07523_ _02684_ _03404_ _04083_ _03261_ _02667_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__o32a_1
XANTENNA__08656__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143__795 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__inv_2
X_07454_ _03861_ _03962_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__a21oi_1
X_06405_ _03060_ _03061_ net758 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XANTENNA__09012__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08408__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07385_ net482 _04040_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1066_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ top0.CPU.register.registers\[76\] net575 _04754_ vssd1 vssd1 vccd1 vccd1
+ _04834_ sky130_fd_sc_hd__o21a_1
XANTENNA__09081__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06336_ top0.CPU.register.registers\[157\] top0.CPU.register.registers\[189\] top0.CPU.register.registers\[221\]
+ top0.CPU.register.registers\[253\] net841 net806 vssd1 vssd1 vccd1 vccd1 _02993_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09055_ _04676_ net269 net255 net2652 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__a22o_1
XANTENNA__11625__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06267_ net772 _02915_ _02919_ _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__o2bb2a_2
X_08006_ _04232_ net233 net228 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__nand3b_1
Xhold530 top0.CPU.register.registers\[824\] vssd1 vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 top0.CPU.register.registers\[467\] vssd1 vssd1 vccd1 vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
X_06198_ top0.CPU.register.registers\[660\] top0.CPU.register.registers\[692\] top0.CPU.register.registers\[724\]
+ top0.CPU.register.registers\[756\] net833 net798 vssd1 vssd1 vccd1 vccd1 _02855_
+ sky130_fd_sc_hd__mux4_1
Xhold563 top0.CPU.register.registers\[348\] vssd1 vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 top0.CPU.register.registers\[346\] vssd1 vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold596 top0.CPU.register.registers\[525\] vssd1 vssd1 vccd1 vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 top0.CPU.register.registers\[663\] vssd1 vssd1 vccd1 vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 top0.CPU.register.registers\[209\] vssd1 vssd1 vccd1 vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ top0.CPU.internalMem.pcOut\[25\] _05448_ vssd1 vssd1 vccd1 vccd1 _05450_
+ sky130_fd_sc_hd__or2_1
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ net720 net167 net278 net283 net2529 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08344__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__A0 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ top0.CPU.internalMem.pcOut\[20\] _05385_ vssd1 vssd1 vccd1 vccd1 _05386_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09670__A2_N net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10151__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__A2 _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ net207 net3017 net354 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__mux2_1
XFILLER_73_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11850_ net1542 _01489_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[343\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08647__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09270__X _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net1473 _01420_ net1035 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout913_X net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ net2094 _02041_ net1051 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[895\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09072__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10206__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ net2025 _01972_ net964 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05686__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12264_ net1956 _01903_ net1076 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[757\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
X_12195_ net1887 _01834_ net1032 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951__603 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__inv_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
X_10028_ _05497_ _05514_ _05512_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08335__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086__738 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__inv_2
XFILLER_64_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127__779 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__inv_2
XANTENNA__09621__A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06992__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07412__Y _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ net1671 _01618_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[472\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07846__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07170_ net446 net539 _03022_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__nor3b_1
XANTENNA__09063__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06121_ top0.CPU.register.registers\[782\] top0.CPU.register.registers\[814\] top0.CPU.register.registers\[846\]
+ top0.CPU.register.registers\[878\] net836 net800 vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08810__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06052_ top0.CPU.register.registers\[392\] top0.CPU.register.registers\[424\] top0.CPU.register.registers\[456\]
+ top0.CPU.register.registers\[488\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02709_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_120_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06191__S net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout328 _04737_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
X_09811_ top0.CPU.internalMem.pcOut\[13\] net648 _05312_ _05315_ vssd1 vssd1 vccd1
+ vccd1 _02190_ sky130_fd_sc_hd__o22a_1
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
X_10694__346 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__inv_2
Xfanout317 _04737_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
Xfanout306 net313 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_4
X_09742_ _05246_ _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkload11_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09007__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06954_ net753 _03606_ net859 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__o21ai_1
X_09673_ _02536_ _04619_ net590 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__mux2_1
X_06885_ _03524_ net525 vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout274_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08877__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05905_ top0.CPU.register.registers\[514\] top0.CPU.register.registers\[546\] top0.CPU.register.registers\[578\]
+ top0.CPU.register.registers\[610\] net824 net789 vssd1 vssd1 vccd1 vccd1 _02562_
+ sky130_fd_sc_hd__mux4_1
X_10735__387 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__inv_2
X_05836_ net743 _02492_ _02485_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__a21oi_4
X_08624_ net714 net162 net309 net330 net2515 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__a32o_1
XANTENNA__06432__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08846__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ _02397_ _02398_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__or2_4
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05767_ net943 net944 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__and2b_2
XFILLER_70_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08629__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _04155_ _04159_ _04161_ _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout539_A _03037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10588__240 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__inv_2
X_05698_ top0.MMIO.WBData_i\[8\] vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__inv_2
XANTENNA__07837__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__A2 _03173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08147__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08486_ net153 net617 net394 net370 net2339 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05848__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout706_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__S1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ net337 _03994_ _04093_ net476 _03841_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__a221o_1
XANTENNA__07986__A _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09054__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10629__281 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__inv_2
X_07368_ net480 _04023_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a21oi_2
XFILLER_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06319_ top0.CPU.register.registers\[284\] top0.CPU.register.registers\[316\] top0.CPU.register.registers\[348\]
+ top0.CPU.register.registers\[380\] net832 net797 vssd1 vssd1 vccd1 vccd1 _02976_
+ sky130_fd_sc_hd__mux4_1
X_09107_ _04697_ net267 net251 net2547 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07299_ _03933_ _03945_ _03946_ _03947_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_111_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ net176 net613 _04806_ net351 net3227 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__a32o_1
XFILLER_123_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold371 top0.CPU.register.registers\[708\] vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 top0.CPU.register.registers\[213\] vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 top0.CPU.register.registers\[351\] vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09706__A top0.CPU.control.funct7\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold393 top0.CPU.register.registers\[722\] vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06114__B _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__A1 _04528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout851 net853 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_4
XFILLER_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
Xfanout873 top0.CPU.decoder.instruction\[17\] vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_4
Xfanout862 net868 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_4
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_51_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08868__A2 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 net904 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
Xhold1060 top0.CPU.register.registers\[205\] vssd1 vssd1 vccd1 vccd1 net3282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1093 top0.CPU.register.registers\[211\] vssd1 vssd1 vccd1 vccd1 net3315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 top0.display.dataforOutput\[13\] vssd1 vssd1 vccd1 vccd1 net3293 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net1594 _01541_ net1007 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[395\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1082 top0.display.dataforOutput\[7\] vssd1 vssd1 vccd1 vccd1 net3304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06423__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ net1525 _01472_ net998 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07540__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08096__A3 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ net1456 _01403_ net961 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[257\]
+ sky130_fd_sc_hd__dfrtp_1
X_11695_ net1387 _01334_ net1001 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[188\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12316_ net2008 _01955_ net1020 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[809\]
+ sky130_fd_sc_hd__dfrtp_1
X_12247_ net1939 _01886_ net972 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[740\]
+ sky130_fd_sc_hd__dfrtp_1
X_12178_ net1870 _01817_ net1053 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[671\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_69_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06414__S0 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06670_ top0.CPU.register.registers\[897\] top0.CPU.register.registers\[929\] top0.CPU.register.registers\[961\]
+ top0.CPU.register.registers\[993\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03327_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_82_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08340_ net721 net194 net401 net411 net2335 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a32o_1
XANTENNA__06717__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08492__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08271_ net221 net671 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and2_1
XANTENNA__06130__A1_N net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ _03729_ _03733_ net456 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux2_1
X_10445__97 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__inv_2
XANTENNA__09036__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07153_ _02579_ _02597_ _03356_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__or3_1
X_06104_ _02759_ _02760_ net734 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XFILLER_106_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ net578 _03718_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__or2_1
X_06035_ top0.CPU.register.registers\[137\] top0.CPU.register.registers\[169\] top0.CPU.register.registers\[201\]
+ top0.CPU.register.registers\[233\] net847 net812 vssd1 vssd1 vccd1 vccd1 _02692_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_93_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
Xfanout147 _04931_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
Xfanout114 _05649_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout169 _04615_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_2
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07986_ _04248_ net232 net228 vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__and3_1
XANTENNA__05766__D1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout158 _04630_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
XANTENNA__06653__S0 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__inv_2
X_06937_ top0.CPU.register.registers\[25\] top0.CPU.register.registers\[57\] top0.CPU.register.registers\[89\]
+ top0.CPU.register.registers\[121\] net909 net875 vssd1 vssd1 vccd1 vccd1 _03594_
+ sky130_fd_sc_hd__mux4_1
X_09656_ top0.MISOtoMMIO\[6\] net3377 _05173_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08607_ net2982 net332 net327 _04551_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a22o_1
XANTENNA__08576__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06868_ top0.CPU.register.registers\[905\] top0.CPU.register.registers\[937\] top0.CPU.register.registers\[969\]
+ top0.CPU.register.registers\[1001\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03525_
+ sky130_fd_sc_hd__mux4_1
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06956__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ top0.CPU.register.registers\[140\] top0.CPU.register.registers\[172\] top0.CPU.register.registers\[204\]
+ top0.CPU.register.registers\[236\] net939 net905 vssd1 vssd1 vccd1 vccd1 _03456_
+ sky130_fd_sc_hd__mux4_1
X_05819_ _02475_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__inv_2
X_09587_ top0.display.state\[0\] _05129_ _05128_ net666 vssd1 vssd1 vccd1 vccd1 _01128_
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout823_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ net198 net675 net404 net363 net2619 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a32o_1
XANTENNA__06096__S net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _04685_ net388 net369 net2884 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22o_1
XANTENNA__08483__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ clknet_leaf_85_clk _01123_ net1107 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_07_1161 vssd1 vssd1 vccd1 vccd1 team_07_1161/HI gpio_out[27] sky130_fd_sc_hd__conb_1
Xteam_07_1150 vssd1 vssd1 vccd1 vccd1 team_07_1150/HI gpio_out[16] sky130_fd_sc_hd__conb_1
Xteam_07_1172 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] team_07_1172/LO sky130_fd_sc_hd__conb_1
XANTENNA__08235__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1194 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] team_07_1194/LO sky130_fd_sc_hd__conb_1
XANTENNA__10042__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1183 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] team_07_1183/LO sky130_fd_sc_hd__conb_1
X_12101_ net1793 _01740_ net1039 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[594\]
+ sky130_fd_sc_hd__dfrtp_1
X_10293_ net3153 net117 net114 _05599_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a22o_1
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ net1724 _01671_ net1042 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold190 top0.CPU.register.registers\[623\] vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11474__Q top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout670 net671 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 net689 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_2
Xfanout692 net700 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06947__S1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11816_ net1508 _01455_ net1075 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[309\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08474__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11747_ net1439 _01386_ net1016 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06485__C1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11678_ net1370 _01317_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[171\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09018__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12587__RESET_B net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__Y _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _03913_ net230 net225 vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and3_1
XANTENNA__09633__X _05162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07771_ net489 _04237_ _04238_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__a21bo_1
X_09510_ _02353_ _02354_ top0.MMIO.WBData_i\[22\] top0.MMIO.WBData_i\[24\] net148
+ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__o41a_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06722_ net745 _03372_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09441_ net143 net139 _05036_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__and3_1
X_06653_ top0.CPU.register.registers\[130\] top0.CPU.register.registers\[162\] top0.CPU.register.registers\[194\]
+ top0.CPU.register.registers\[226\] net914 net880 vssd1 vssd1 vccd1 vccd1 _03310_
+ sky130_fd_sc_hd__mux4_1
X_09372_ net2622 _04557_ net607 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__mux2_1
X_06584_ net860 _03232_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a21oi_4
X_08323_ net3079 net412 net405 _04488_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08465__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10847__499 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__inv_2
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08480__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08254_ net3193 net417 _04712_ net492 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XANTENNA__09020__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05768__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ net498 net215 net615 net425 net2435 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a32o_1
X_07205_ net489 net480 _03860_ _03838_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_95_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07136_ net529 net533 net468 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__mux2_1
XFILLER_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08232__A3 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _03317_ _03301_ net471 vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__mux2_1
XFILLER_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06018_ net778 _02670_ _02673_ _02674_ net773 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__o221a_1
XANTENNA__07328__X _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout773_A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750__402 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__inv_2
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout940_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ top0.CPU.internalMem.pcOut\[6\] _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__nand2_1
X_07969_ top0.CPU.internalMem.pcOut\[8\] net641 net636 _04602_ vssd1 vssd1 vccd1 vccd1
+ _04603_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06819__S net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07063__X _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ _02787_ _05151_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nor2_1
XANTENNA__07504__A _02769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06929__S1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12650_ clknet_leaf_71_clk _02285_ net1122 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07998__X _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11601_ net1293 _01240_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08456__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ clknet_leaf_83_clk _02216_ net1110 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ net1224 _01171_ net966 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06554__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ clknet_leaf_74_clk _01111_ net1125 vssd1 vssd1 vccd1 vccd1 top0.CPU.control.rs2\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08759__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__Q top0.CPU.control.funct7\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11394_ clknet_leaf_57_clk _01042_ net1089 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07431__A1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ net2246 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07893__B net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ _04936_ _05162_ _04930_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__or3b_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05993__A1 top0.CPU.control.funct7\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07238__X _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06617__S0 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ net1707 _01654_ net996 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[508\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09184__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493__145 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__inv_2
XANTENNA__05745__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07042__S0 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05876__A1_N top0.CPU.control.funct7\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10534__186 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__inv_2
XFILLER_34_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__A2 top0.CPU.addrControl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12779_ top0.chipSelectTFT vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08245__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07670__A1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 top0.CPU.register.registers\[904\] vssd1 vssd1 vccd1 vccd1 net3126 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_12_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10415__67 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__inv_2
Xhold926 top0.CPU.register.registers\[783\] vssd1 vssd1 vccd1 vccd1 net3148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold937 top0.display.dataforOutput\[15\] vssd1 vssd1 vccd1 vccd1 net3159 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold915 top0.CPU.register.registers\[244\] vssd1 vssd1 vccd1 vccd1 net3137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06856__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09990_ _05440_ _05449_ _05450_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__and4_1
Xhold959 top0.CPU.register.registers\[1006\] vssd1 vssd1 vccd1 vccd1 net3181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 top0.CPU.register.registers\[273\] vssd1 vssd1 vccd1 vccd1 net3170 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08941_ net193 net711 _04779_ net265 net3282 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_90_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08872_ _04499_ net554 _04757_ net282 net3006 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__a32o_1
X_07823_ top0.CPU.intMem_out\[31\] net628 vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__nand2_1
XFILLER_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06084__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__C1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07754_ _04401_ _04402_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__a21o_1
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06639__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07685_ net344 _03942_ _04332_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o31ai_1
XANTENNA__08686__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ _03285_ net531 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__nand2_1
X_09424_ net3397 net599 net132 _05027_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_91_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout354_A _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06636_ net863 _03288_ _03291_ _03292_ net745 vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__a221o_1
XANTENNA__08854__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ net3128 _04631_ net611 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
X_06567_ _03202_ _03204_ _03222_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__and3_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout521_A _03637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ top0.CPU.internalMem.loadCt\[0\] _04944_ vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.loadCt_n\[0\]
+ sky130_fd_sc_hd__and2b_1
X_08306_ net2907 _04581_ net415 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
XANTENNA__10245__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06498_ _03094_ _03115_ _03132_ _03153_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__or4b_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ net493 net159 net679 net421 net2404 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08168_ net3014 net428 _04684_ net516 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
XFILLER_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11270__922 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__inv_2
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08610__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ net504 net177 net691 net433 net2301 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a32o_1
X_07119_ _02579_ _02597_ net523 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__or3_1
XFILLER_133_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10130_ _04957_ _05594_ net661 vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__o21a_1
X_10477__129 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__inv_2
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10061_ top0.display.delayctr\[5\] _05539_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311__963 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__inv_2
XFILLER_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08913__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05822__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07024__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_82_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_39_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08692__A3 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12633_ clknet_leaf_71_clk _02268_ net1119 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_61_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05689__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12564_ clknet_leaf_55_clk _02203_ net1038 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_11515_ net1207 _01154_ net1008 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07652__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05889__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ net2187 _02134_ net1001 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[988\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12108__RESET_B net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ clknet_leaf_70_clk _01094_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.Op\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_11377_ clknet_leaf_73_clk top0.CPU.internalMem.loadCt_n\[1\] net1127 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.loadCt\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06838__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08601__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07955__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05855__C _02511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10328_ net2251 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08904__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ net3237 net117 net111 _05652_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
XFILLER_22_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06066__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05813__S1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08380__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08668__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08683__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07431__X _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ net342 _04108_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_17_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07891__A1 top0.CPU.intMem_out\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06421_ _02457_ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__xnor2_1
X_06352_ _02454_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__nor2_1
X_09140_ top0.CPU.register.registers\[66\] net565 net160 net680 net553 vssd1 vssd1
+ vccd1 vccd1 _04840_ sky130_fd_sc_hd__o2111a_1
X_09071_ top0.CPU.register.registers\[112\] net570 net557 vssd1 vssd1 vccd1 vccd1
+ _04817_ sky130_fd_sc_hd__o21a_1
X_11254__906 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__inv_2
X_06283_ top0.CPU.register.registers\[26\] top0.CPU.register.registers\[58\] top0.CPU.register.registers\[90\]
+ top0.CPU.register.registers\[122\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02940_
+ sky130_fd_sc_hd__mux4_1
XFILLER_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08022_ net209 net701 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__and2_1
Xhold701 top0.CPU.register.registers\[948\] vssd1 vssd1 vccd1 vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 top0.CPU.register.registers\[603\] vssd1 vssd1 vccd1 vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold723 top0.CPU.intMemAddr\[10\] vssd1 vssd1 vccd1 vccd1 net2945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold745 top0.CPU.register.registers\[314\] vssd1 vssd1 vccd1 vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 top0.CPU.register.registers\[769\] vssd1 vssd1 vccd1 vccd1 net2956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold767 top0.CPU.intMemAddr\[23\] vssd1 vssd1 vccd1 vccd1 net2989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05765__C net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold756 net71 vssd1 vssd1 vccd1 vccd1 net2978 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _05462_ _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__or2_1
Xhold778 top0.CPU.register.registers\[762\] vssd1 vssd1 vccd1 vccd1 net3000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold789 top0.CPU.register.registers\[503\] vssd1 vssd1 vccd1 vccd1 net3011 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ _04642_ net552 _04775_ net263 net3030 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1011_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__X _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148__800 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__inv_2
X_08855_ net220 net3295 net355 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__mux2_1
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08371__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ net183 net685 net323 net291 net2812 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a32o_1
XANTENNA__06369__S net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ net535 _03262_ net532 net529 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout569_A _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05998_ top0.CPU.register.registers\[775\] top0.CPU.register.registers\[807\] top0.CPU.register.registers\[839\]
+ top0.CPU.register.registers\[871\] net842 net807 vssd1 vssd1 vccd1 vccd1 _02655_
+ sky130_fd_sc_hd__mux4_1
X_07737_ _02577_ _03869_ _04393_ net244 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_64_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_111_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout736_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__B1 _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08584__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _03747_ _03759_ _04324_ net452 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06619_ top0.CPU.register.registers\[133\] top0.CPU.register.registers\[165\] top0.CPU.register.registers\[197\]
+ top0.CPU.register.registers\[229\] net934 net900 vssd1 vssd1 vccd1 vccd1 _03276_
+ sky130_fd_sc_hd__mux4_1
X_09407_ top0.MMIO.WBData_i\[2\] net147 net143 top0.MISOtoMMIO\[2\] _05014_ vssd1
+ vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_101_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09627__A_N _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10862__514 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__inv_2
X_07599_ net337 _04077_ _04255_ net476 vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__a22o_1
X_09338_ top0.CPU.internalMem.state\[3\] _04850_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__nor2_1
XANTENNA__09084__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07501__B _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__A1 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903__555 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__inv_2
X_09269_ _04865_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__nand2b_1
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ net1972 _01919_ net1029 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[773\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09387__A1 _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10113_ net3423 net667 _05141_ _05578_ _05581_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a221o_1
XANTENNA__06296__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _05527_ _05530_ top0.CPU.internalMem.pcOut\[31\] net645 vssd1 vssd1 vccd1
+ vccd1 _02208_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06911__A2_N _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 top0.CPU.register.registers\[544\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 top0.CPU.register.registers\[618\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06787__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 top0.CPU.register.registers\[678\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 top0.CPU.register.registers\[35\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 top0.CPU.register.registers\[707\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ net1687 _01634_ net1015 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[488\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_55_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10102__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07899__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ clknet_leaf_80_clk _02251_ net1113 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08417__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ clknet_leaf_60_clk _02186_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_10646__298 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__inv_2
XANTENNA__08822__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ net2170 _02117_ net1014 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[971\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09619__A _02715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _04333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11429_ clknet_leaf_60_clk _01077_ net1094 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10499__151 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__inv_2
XFILLER_112_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06970_ net866 _03626_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
XANTENNA__06039__S1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05921_ net487 net479 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__nand2_2
X_05852_ top0.CPU.register.registers\[271\] top0.CPU.register.registers\[303\] top0.CPU.register.registers\[335\]
+ top0.CPU.register.registers\[367\] net851 net816 vssd1 vssd1 vccd1 vccd1 _02509_
+ sky130_fd_sc_hd__mux4_1
X_08640_ _04649_ net327 net304 net2774 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a22o_1
Xfanout1092 net1106 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_2
Xfanout1081 net1083 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
Xfanout1070 net1088 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_2
XFILLER_27_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05783_ net772 _02439_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__and2_1
X_08571_ net2940 net222 net333 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_35_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09801__B _02734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07522_ _04177_ _04178_ _04167_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__o21bai_1
XFILLER_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07864__A1 top0.CPU.intMem_out\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08656__A3 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ net490 _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__and2_1
X_06404_ top0.CPU.register.registers\[796\] top0.CPU.register.registers\[828\] top0.CPU.register.registers\[860\]
+ top0.CPU.register.registers\[892\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03061_
+ sky130_fd_sc_hd__mux4_1
XFILLER_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09123_ net193 net686 _04833_ net253 net3273 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a32o_1
XANTENNA__08408__A3 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ net488 _04037_ _03743_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21o_1
XANTENNA__08813__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06335_ net781 _02987_ _02990_ _02991_ net771 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__o221ai_4
XANTENNA_fanout317_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07092__A2 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _04675_ net553 _04811_ net256 net3047 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__a32o_1
X_06266_ net735 _02922_ net741 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__o21ai_1
X_08005_ _04232_ _04474_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__nor2_1
Xhold520 top0.CPU.register.registers\[347\] vssd1 vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 top0.CPU.register.registers\[863\] vssd1 vssd1 vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 top0.CPU.register.registers\[958\] vssd1 vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
X_06197_ _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__inv_2
Xhold542 top0.CPU.register.registers\[343\] vssd1 vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 top0.CPU.register.registers\[307\] vssd1 vssd1 vccd1 vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold586 net46 vssd1 vssd1 vccd1 vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 top0.CPU.register.registers\[306\] vssd1 vssd1 vccd1 vccd1 net2797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold597 top0.CPU.register.registers\[465\] vssd1 vssd1 vccd1 vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08579__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__B _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ top0.CPU.internalMem.pcOut\[25\] _05448_ vssd1 vssd1 vccd1 vccd1 _05449_
+ sky130_fd_sc_hd__nand2_1
X_09887_ _02854_ _04541_ net586 vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__mux2_1
XANTENNA__05792__A _02338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ net714 net171 _04770_ net282 net3353 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__a32o_1
Xhold1220 top0.CPU.intMem_out\[25\] vssd1 vssd1 vccd1 vccd1 net3442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ net208 net3253 net353 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__mux2_1
XANTENNA__06099__S net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__B _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _04693_ net307 net289 net2742 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__a22o_1
X_11780_ net1472 _01419_ net987 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[273\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08647__A3 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12401_ net2093 _02040_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08804__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ net2024 _01971_ net986 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06562__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12263_ net1955 _01902_ net1003 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[756\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08062__B net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ net1886 _01833_ net1047 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[687\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
X_10990__642 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__inv_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__B1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _05497_ _05512_ _05514_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_28_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06441__S1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ net1670 _01617_ net963 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05952__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06120_ net780 _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06051_ top0.CPU.register.registers\[264\] top0.CPU.register.registers\[296\] top0.CPU.register.registers\[328\]
+ top0.CPU.register.registers\[360\] net843 net808 vssd1 vssd1 vccd1 vccd1 _02708_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09636__X _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ net235 _05313_ _05314_ net648 vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09771__B2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net321 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_8
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
X_09741_ top0.CPU.internalMem.pcOut\[8\] _05249_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09554__D_N net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06953_ net866 _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__nor2_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05904_ top0.CPU.register.registers\[642\] top0.CPU.register.registers\[674\] top0.CPU.register.registers\[706\]
+ top0.CPU.register.registers\[738\] net829 net794 vssd1 vssd1 vccd1 vccd1 _02561_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08326__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110__762 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _05179_ _05184_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06884_ _03524_ net525 vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__and2_1
XANTENNA__07316__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05835_ _02488_ _02491_ net738 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_08623_ net715 net164 net309 net329 net2481 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06432__S1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _02397_ _02398_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nor2_1
X_05766_ _02338_ _02375_ _02384_ net632 net626 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__o2111a_1
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07603__Y _04260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout267_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _02750_ _03482_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05697_ top0.MMIO.WBData_i\[4\] vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08147__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08485_ net157 net614 net386 net369 net2320 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a32o_1
X_07436_ _04062_ _04092_ net458 vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__mux2_1
XANTENNA__05943__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ net457 _03859_ _03831_ net347 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__o211a_1
X_06318_ net783 _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nand2_1
X_09106_ _04696_ net555 _04827_ net252 net3025 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_98_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ top0.CPU.register.registers\[135\] net570 vssd1 vssd1 vccd1 vccd1 _04806_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08163__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07298_ net485 _03949_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a21o_1
X_10974__626 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__inv_2
X_06249_ net742 _02905_ _02898_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06943__A1_N net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 top0.CPU.register.registers\[842\] vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
X_10376__28 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__inv_2
Xhold361 top0.CPU.register.registers\[378\] vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 top0.CPU.register.registers\[350\] vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 top0.CPU.register.registers\[297\] vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 top0.CPU.register.registers\[429\] vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_2
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
Xfanout841 top0.CPU.control.rs2\[0\] vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ top0.CPU.internalMem.pcOut\[23\] _05421_ _05432_ vssd1 vssd1 vccd1 vccd1
+ _05433_ sky130_fd_sc_hd__o21a_1
Xfanout885 net907 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_51_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout863 net868 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_2
Xfanout874 net876 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_4
Xhold1050 top0.CPU.register.registers\[109\] vssd1 vssd1 vccd1 vccd1 net3272 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout896 net904 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ net1593 _01540_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold1072 _01144_ vssd1 vssd1 vccd1 vccd1 net3294 sky130_fd_sc_hd__dlygate4sd3_1
X_10868__520 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__inv_2
Xhold1083 _01137_ vssd1 vssd1 vccd1 vccd1 net3305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 top0.CPU.register.registers\[131\] vssd1 vssd1 vccd1 vccd1 net3283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 top0.CPU.register.registers\[887\] vssd1 vssd1 vccd1 vccd1 net3316 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06423__S1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ net1524 _01471_ net1026 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[325\]
+ sky130_fd_sc_hd__dfrtp_1
X_10909__561 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11763_ net1455 _01402_ net1064 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[256\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ net1386 _01333_ net991 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ net2007 _01954_ net1017 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11053__705 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__inv_2
XANTENNA__10108__A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ net1938 _01885_ net994 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[739\]
+ sky130_fd_sc_hd__dfrtp_1
X_12177_ net1869 _01816_ net1093 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08520__B _02400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390__42 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__inv_2
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_69_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06414__S1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06178__S0 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08270_ net512 net197 net675 net419 net2395 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a32o_1
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07221_ _03876_ _03877_ net348 vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__mux2_1
X_07152_ _03807_ _03808_ net464 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__mux2_1
X_10661__313 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__inv_2
X_06103_ top0.CPU.register.registers\[12\] top0.CPU.register.registers\[44\] top0.CPU.register.registers\[76\]
+ top0.CPU.register.registers\[108\] net855 net820 vssd1 vssd1 vccd1 vccd1 _02760_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08244__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__A1_N net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ _02430_ _03718_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_8_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
X_10702__354 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__inv_2
XANTENNA__08795__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06034_ _02687_ _02688_ _02689_ _02690_ net728 net737 vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06930__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06102__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 net140 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout126 net128 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
Xfanout115 _05643_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07327__A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07985_ net721 net509 net169 net547 net2682 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a32o_1
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
XFILLER_87_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06653__S1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout159 _04630_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_09724_ top0.CPU.internalMem.pcOut\[7\] _05233_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__or2_1
XANTENNA__08857__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06936_ top0.CPU.register.registers\[153\] top0.CPU.register.registers\[185\] top0.CPU.register.registers\[217\]
+ top0.CPU.register.registers\[249\] net910 net876 vssd1 vssd1 vccd1 vccd1 _03593_
+ sky130_fd_sc_hd__mux4_1
XFILLER_28_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ net3415 top0.MISOtoMMIO\[6\] _05173_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__mux2_1
X_06867_ _02698_ _03523_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_2_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08180__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05818_ net861 _02474_ _02472_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06885__B net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ net3024 net329 net312 _04545_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a22o_1
X_06798_ net754 _03454_ net861 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__o21ai_1
X_09586_ top0.display.counter\[3\] top0.display.counter\[2\] _05124_ vssd1 vssd1 vccd1
+ vccd1 _05129_ sky130_fd_sc_hd__nand3_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08537_ net201 net673 net400 net363 net2540 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a32o_1
X_05749_ net942 net943 net944 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__or3_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ net203 net623 net400 net371 net2275 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a32o_1
XFILLER_51_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ net524 _03262_ net469 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ _04664_ net392 net378 net2846 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a22o_1
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xteam_07_1151 vssd1 vssd1 vccd1 vccd1 team_07_1151/HI gpio_out[17] sky130_fd_sc_hd__conb_1
Xteam_07_1162 vssd1 vssd1 vccd1 vccd1 team_07_1162/HI gpio_out[28] sky130_fd_sc_hd__conb_1
XFILLER_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_07_1140 vssd1 vssd1 vccd1 vccd1 team_07_1140/HI gpio_out[6] sky130_fd_sc_hd__conb_1
XANTENNA__08235__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_07_1173 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] team_07_1173/LO sky130_fd_sc_hd__conb_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_07_1195 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] team_07_1195/LO sky130_fd_sc_hd__conb_1
Xteam_07_1184 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] team_07_1184/LO sky130_fd_sc_hd__conb_1
XANTENNA__08786__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09276__X _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ net3211 net119 net112 _05666_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a22o_1
X_12100_ net1792 _01739_ net989 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[593\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07994__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ net1723 _01670_ net1102 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[524\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 top0.CPU.register.registers\[104\] vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06267__A1_N net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 top0.CPU.register.registers\[875\] vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout660 _04955_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout682 net689 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_4
Xfanout693 net700 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_4
Xfanout671 net678 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ net1507 _01454_ net1031 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[308\]
+ sky130_fd_sc_hd__dfrtp_1
X_11746_ net1438 _01385_ net1045 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05979__X _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05907__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ net1369 _01316_ net1022 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06580__S0 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net1921 _01868_ net1037 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08529__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12556__RESET_B net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07201__A2 _03053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07770_ net442 _04145_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nor2_1
X_06721_ net858 _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__or2_1
X_11181__833 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__inv_2
X_09440_ _05005_ _05006_ _05008_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__10301__A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06652_ net745 _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__or2_1
X_09371_ net2709 _04563_ net607 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__mux2_1
X_06583_ net865 _03235_ _03238_ _03239_ net747 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o221a_1
XANTENNA__05920__C1 _02574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ net721 net151 net404 net411 net2336 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11222__874 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__inv_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ net208 net668 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__and2_1
X_07204_ net481 _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__nand2_1
X_08184_ net509 net169 net621 net428 net2406 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a32o_1
XFILLER_118_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08217__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05768__C net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07135_ _03790_ _03791_ net465 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
XFILLER_134_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1041_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ _03721_ _03722_ net460 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout599_A _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06017_ net729 _02671_ net737 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_7_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_A _02344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08940__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ top0.CPU.intMem_out\[8\] net628 _04476_ _04601_ _02382_ vssd1 vssd1 vccd1
+ vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XFILLER_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08587__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ net590 _04608_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a21o_1
X_06919_ _03562_ _03571_ _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07899_ net715 net223 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ net3328 net605 net659 net3293 _05165_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__a221o_1
XANTENNA__07900__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10830__482 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__inv_2
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ top0.CPU.decoder.instruction\[8\] _02448_ _02535_ net822 net589 vssd1 vssd1
+ vccd1 vccd1 _05116_ sky130_fd_sc_hd__a221o_1
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ clknet_leaf_90_clk _02215_ net1085 vssd1 vssd1 vccd1 vccd1 top0.display.delayctr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11600_ net1292 _01239_ net1078 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_11531_ net1223 _01170_ net1066 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11462_ clknet_leaf_71_clk _01110_ net1119 vssd1 vssd1 vccd1 vccd1 top0.CPU.decoder.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_11393_ clknet_leaf_86_clk _01041_ net1091 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMemAddr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08759__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ net2278 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06314__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10275_ net2869 net121 net114 _05659_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a22o_1
XANTENNA__05993__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__B net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06617__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ net1706 _01653_ net992 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08392__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165__817 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__inv_2
XANTENNA__05745__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout490 _02554_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_2
XANTENNA__08144__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360__12 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__inv_2
XFILLER_0_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07042__S1 top0.CPU.control.rs2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload8_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206__858 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__inv_2
XFILLER_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_12778_ top0.bitDataTFT vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09644__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059__711 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__inv_2
XANTENNA__08998__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11729_ net1421 _01368_ net1048 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08245__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06553__S0 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold927 top0.CPU.register.registers\[671\] vssd1 vssd1 vccd1 vccd1 net3149 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold916 top0.CPU.register.registers\[93\] vssd1 vssd1 vccd1 vccd1 net3138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold905 top0.CPU.register.registers\[859\] vssd1 vssd1 vccd1 vccd1 net3127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05885__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06856__S1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold938 _01145_ vssd1 vssd1 vccd1 vccd1 net3160 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06480__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold949 top0.CPU.register.registers\[1009\] vssd1 vssd1 vccd1 vccd1 net3171 sky130_fd_sc_hd__dlygate4sd3_1
X_08940_ top0.CPU.register.registers\[205\] net572 net558 vssd1 vssd1 vccd1 vccd1
+ _04779_ sky130_fd_sc_hd__o21a_1
X_10773__425 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09175__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ top0.CPU.register.registers\[252\] net566 vssd1 vssd1 vccd1 vccd1 _04757_
+ sky130_fd_sc_hd__or2_1
X_07822_ net591 _03686_ _04478_ net627 vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a211o_1
XFILLER_57_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08922__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814__466 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__inv_2
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ _04407_ _04408_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_121_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07684_ _04338_ _04339_ _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__and3_1
X_06704_ _03320_ _03360_ _03319_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a21o_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09423_ top0.MMIO.WBData_i\[8\] _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__and2_1
X_06635_ net758 _03289_ net750 vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__o21a_1
XANTENNA__06792__S0 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ net34 net36 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.nrst sky130_fd_sc_hd__and2_1
XANTENNA_fanout1089_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout347_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06566_ _03202_ _03204_ _03222_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07340__A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06655__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ net2947 net221 net414 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ top0.CPU.internalMem.state\[1\] top0.CPU.internalMem.state\[0\] _04852_ vssd1
+ vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__and3_1
XANTENNA__10245__B2 top0.MMIO.WBData_i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08989__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06497_ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__inv_2
XANTENNA__08155__B net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708__360 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__inv_2
X_08236_ net497 net161 net680 net421 net2623 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08167_ _04549_ _04671_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ net482 net478 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_132_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08610__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ net506 net219 net694 net434 net2758 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout883_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07049_ _03006_ _03022_ net541 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09166__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10060_ net3402 net663 _05143_ _05541_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a211o_1
XANTENNA__08374__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08110__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07024__S1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_39_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06783__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12632_ clknet_leaf_71_clk _02267_ net1122 vssd1 vssd1 vccd1 vccd1 top0.MMIO.WBData_i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_61_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08429__A1 _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12563_ clknet_leaf_55_clk _02202_ net1038 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_11514_ net1206 _01153_ net975 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12494_ net2186 _02133_ net991 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[987\]
+ sky130_fd_sc_hd__dfrtp_1
X_11445_ clknet_leaf_78_clk _01093_ net1116 vssd1 vssd1 vccd1 vccd1 top0.CPU.Op\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_10460__112 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__inv_2
X_11376_ clknet_leaf_73_clk top0.CPU.internalMem.loadCt_n\[0\] net1127 vssd1 vssd1
+ vccd1 vccd1 top0.CPU.internalMem.loadCt\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06838__S1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757__409 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10327_ net2224 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__05992__X _02649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ _04938_ _05136_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__or2_1
X_10501__153 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08365__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ net129 _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and2_1
XANTENNA__09624__B _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08380__A3 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__09640__A _05141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06420_ _02497_ _02834_ _02870_ _02889_ net541 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__o41a_1
XANTENNA__06774__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06351_ top0.CPU.control.funct7\[5\] _02374_ _02377_ vssd1 vssd1 vccd1 vccd1 _03008_
+ sky130_fd_sc_hd__and3_1
X_11293__945 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__inv_2
X_06282_ top0.CPU.register.registers\[154\] top0.CPU.register.registers\[186\] top0.CPU.register.registers\[218\]
+ top0.CPU.register.registers\[250\] net823 net788 vssd1 vssd1 vccd1 vccd1 _02939_
+ sky130_fd_sc_hd__mux4_1
X_09070_ _04685_ net269 net255 net2493 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__a22o_1
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ net3141 net437 _04641_ net494 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
Xhold702 top0.CPU.register.registers\[514\] vssd1 vssd1 vccd1 vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 top0.CPU.register.registers\[652\] vssd1 vssd1 vccd1 vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 top0.CPU.register.registers\[979\] vssd1 vssd1 vccd1 vccd1 net2968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 top0.CPU.intMemAddr\[7\] vssd1 vssd1 vccd1 vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 top0.CPU.register.registers\[889\] vssd1 vssd1 vccd1 vccd1 net2935 sky130_fd_sc_hd__dlygate4sd3_1
X_11334__986 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__inv_2
Xhold779 top0.CPU.register.registers\[115\] vssd1 vssd1 vccd1 vccd1 net3001 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09972_ _05441_ _05463_ _05450_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__o21a_1
Xhold757 top0.CPU.register.registers\[526\] vssd1 vssd1 vccd1 vccd1 net2979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 top0.CPU.register.registers\[821\] vssd1 vssd1 vccd1 vccd1 net2990 sky130_fd_sc_hd__dlygate4sd3_1
X_08923_ top0.CPU.register.registers\[218\] net564 vssd1 vssd1 vccd1 vccd1 _04775_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08356__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08854_ net180 net3175 net356 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1004_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09026__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ net187 net684 net321 net291 net2462 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a32o_1
X_07805_ net523 net522 net520 _04461_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__and4_1
X_05997_ _02652_ _02653_ net725 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XFILLER_72_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout464_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07736_ net338 _03870_ _04392_ net483 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a22o_1
X_11228__880 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__inv_2
XANTENNA_fanout729_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _04091_ _04101_ net486 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06618_ top0.CPU.register.registers\[389\] top0.CPU.register.registers\[421\] top0.CPU.register.registers\[453\]
+ top0.CPU.register.registers\[485\] net932 net898 vssd1 vssd1 vccd1 vccd1 _03275_
+ sky130_fd_sc_hd__mux4_1
X_09406_ net3394 _04949_ _05016_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_101_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07598_ _04116_ _04254_ net458 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__mux2_1
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09337_ _04851_ _04863_ _04973_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__a22o_1
XFILLER_40_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06549_ top0.CPU.register.registers\[529\] top0.CPU.register.registers\[561\] top0.CPU.register.registers\[593\]
+ top0.CPU.register.registers\[625\] net911 net877 vssd1 vssd1 vccd1 vccd1 _03206_
+ sky130_fd_sc_hd__mux4_1
X_09268_ _04893_ _04897_ _04925_ _04928_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and4b_1
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10942__594 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__inv_2
X_08219_ net222 net679 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__and2_1
X_09199_ _04861_ vssd1 vssd1 vccd1 vccd1 top0.CPU.busy sky130_fd_sc_hd__inv_2
XFILLER_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07398__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05875__A1_N net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10112_ _05579_ _05580_ net600 vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09139__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_112_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _05528_ _05529_ _05110_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a21o_1
Xhold40 top0.CPU.register.registers\[946\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 top0.CPU.register.registers\[607\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 top0.CPU.register.registers\[838\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 top0.CPU.register.registers\[548\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 top0.CPU.register.registers\[300\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold84 top0.CPU.intMemAddr\[1\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11994_ net1686 _01633_ net975 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06756__S0 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11277__929 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__inv_2
X_12615_ clknet_leaf_80_clk _02250_ net1113 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
X_11021__673 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__inv_2
XFILLER_129_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ clknet_leaf_69_clk _02185_ net1099 vssd1 vssd1 vccd1 vccd1 top0.CPU.internalMem.pcOut\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_138_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ net2169 _02116_ net1023 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[970\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09619__B _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ clknet_leaf_61_clk _01076_ net1098 vssd1 vssd1 vccd1 vccd1 top0.CPU.intMem_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05920_ _02552_ _02553_ _02573_ _02574_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__o211a_2
X_05851_ top0.CPU.register.registers\[399\] top0.CPU.register.registers\[431\] top0.CPU.register.registers\[463\]
+ top0.CPU.register.registers\[495\] net851 net816 vssd1 vssd1 vccd1 vccd1 _02508_
+ sky130_fd_sc_hd__mux4_1
XFILLER_94_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout1071 net1074 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08353__A3 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1065 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1093 net1106 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08570_ net2699 _04555_ net335 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XANTENNA__09641__Y _05168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06995__S0 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07521_ net346 _03317_ _04169_ net531 net484 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a32o_1
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10885__537 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__inv_2
X_05782_ _02435_ _02436_ _02437_ _02438_ net726 net736 vssd1 vssd1 vccd1 vccd1 _02439_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08510__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07849__C1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08105__A3 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07452_ _04023_ _04039_ net478 vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__mux2_1
X_06403_ top0.CPU.register.registers\[924\] top0.CPU.register.registers\[956\] top0.CPU.register.registers\[988\]
+ top0.CPU.register.registers\[1020\] net917 net883 vssd1 vssd1 vccd1 vccd1 _03060_
+ sky130_fd_sc_hd__mux4_1
X_10926__578 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__inv_2
X_07383_ _04038_ _04039_ net345 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__mux2_1
X_09122_ top0.CPU.register.registers\[77\] net572 net558 vssd1 vssd1 vccd1 vccd1 _04833_
+ sky130_fd_sc_hd__o21a_1
XFILLER_50_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06334_ net732 _02988_ net739 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a21o_1
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06933__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06824__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ top0.CPU.register.registers\[124\] net565 vssd1 vssd1 vccd1 vccd1 _04811_
+ sky130_fd_sc_hd__or2_1
X_06265_ _02920_ _02921_ net724 vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__mux2_1
X_10779__431 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__inv_2
X_06196_ net857 net644 _02454_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a21oi_2
X_08004_ net713 net493 net159 net546 net2680 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a32o_1
Xhold510 top0.CPU.register.registers\[185\] vssd1 vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 top0.CPU.register.registers\[723\] vssd1 vssd1 vccd1 vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 top0.CPU.register.registers\[905\] vssd1 vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold554 top0.CPU.register.registers\[598\] vssd1 vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 top0.CPU.register.registers\[602\] vssd1 vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 top0.CPU.register.registers\[169\] vssd1 vssd1 vccd1 vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold587 top0.CPU.register.registers\[475\] vssd1 vssd1 vccd1 vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 top0.CPU.register.registers\[57\] vssd1 vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ net585 _04512_ _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a21o_1
Xhold598 top0.CPU.register.registers\[711\] vssd1 vssd1 vccd1 vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
X_09886_ top0.CPU.internalMem.pcOut\[19\] net647 _05384_ vssd1 vssd1 vccd1 vccd1 _02196_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA__05792__B top0.CPU.Op\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ top0.CPU.register.registers\[230\] net565 net553 vssd1 vssd1 vccd1 vccd1
+ _04770_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout679_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1210 top0.CPU.intMem_out\[21\] vssd1 vssd1 vccd1 vccd1 net3432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 top0.CPU.intMem_out\[14\] vssd1 vssd1 vccd1 vccd1 net3443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08344__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08837_ net209 net3121 net353 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout846_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08768_ _04692_ net311 net289 net2785 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07304__A1 _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ net453 _03850_ _03949_ _04372_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__o311a_1
X_08699_ net211 net3179 net357 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__mux2_1
XANTENNA__08501__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07304__B2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06409__A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005__657 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__inv_2
X_12400_ net2092 _02039_ net1080 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ net2023 _01970_ net1072 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[824\]
+ sky130_fd_sc_hd__dfrtp_1
X_12262_ net1954 _01901_ net1126 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[755\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12193_ net1885 _01832_ net1063 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[686\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_1_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07791__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572__224 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__inv_2
X_10026_ _05484_ _05489_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08335__A3 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06977__S0 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10613__265 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__inv_2
X_11977_ net1669 _01616_ net1062 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[470\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07846__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05952__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09599__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12529_ net2221 _02168_ net1049 vssd1 vssd1 vccd1 vccd1 top0.CPU.register.registers\[1022\]
+ sky130_fd_sc_hd__dfrtp_1
X_06050_ net778 _02702_ _02705_ _02706_ net773 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__o221a_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08253__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08023__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_87_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05893__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net313 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
X_09740_ _05248_ top0.CPU.internalMem.pcOut\[8\] _05247_ vssd1 vssd1 vccd1 vccd1 _05250_
+ sky130_fd_sc_hd__nand3b_1
X_06952_ _03607_ _03608_ net764 vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__mux2_1
.ends

