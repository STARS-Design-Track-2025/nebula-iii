`default_nettype none
module t01_ai_MMU_new (
    
); 

  logic [127:0][3:0] d0_w;
  logic [31:0][3:0] d0_b;
  logic [1023:0][3:0] d1_w;
  logic [31:0][3:0] d1_b;
  logic [1023:0][3:0] d2_w;
  logic [31:0][3:0] d2_b;
  logic [31:0][3:0] d3_w;
  logic [3:0] d3_b;
    // --- layer0_w ---
    assign d0_w[0] = 4'h3;
    assign d0_w[1] = 4'h0;
    assign d0_w[2] = 4'hC;
    assign d0_w[3] = 4'h3;
    assign d0_w[4] = 4'hA;
    assign d0_w[5] = 4'h2;
    assign d0_w[6] = 4'h9;
    assign d0_w[7] = 4'hC;
    assign d0_w[8] = 4'hD;
    assign d0_w[9] = 4'hC;
    assign d0_w[10] = 4'hD;
    assign d0_w[11] = 4'hF;
    assign d0_w[12] = 4'hF;
    assign d0_w[13] = 4'hC;
    assign d0_w[14] = 4'h1;
    assign d0_w[15] = 4'hE;
    assign d0_w[16] = 4'h1;
    assign d0_w[17] = 4'hD;
    assign d0_w[18] = 4'h1;
    assign d0_w[19] = 4'h5;
    assign d0_w[20] = 4'h2;
    assign d0_w[21] = 4'hB;
    assign d0_w[22] = 4'h0;
    assign d0_w[23] = 4'h1;
    assign d0_w[24] = 4'hE;
    assign d0_w[25] = 4'hE;
    assign d0_w[26] = 4'h0;
    assign d0_w[27] = 4'h4;
    assign d0_w[28] = 4'hB;
    assign d0_w[29] = 4'h2;
    assign d0_w[30] = 4'hE;
    assign d0_w[31] = 4'hE;
    assign d0_w[32] = 4'hE;
    assign d0_w[33] = 4'hB;
    assign d0_w[34] = 4'h4;
    assign d0_w[35] = 4'h3;
    assign d0_w[36] = 4'h6;
    assign d0_w[37] = 4'hF;
    assign d0_w[38] = 4'h4;
    assign d0_w[39] = 4'hF;
    assign d0_w[40] = 4'h1;
    assign d0_w[41] = 4'hC;
    assign d0_w[42] = 4'hE;
    assign d0_w[43] = 4'hF;
    assign d0_w[44] = 4'h7;
    assign d0_w[45] = 4'hC;
    assign d0_w[46] = 4'hB;
    assign d0_w[47] = 4'h4;
    assign d0_w[48] = 4'hB;
    assign d0_w[49] = 4'h1;
    assign d0_w[50] = 4'h1;
    assign d0_w[51] = 4'hD;
    assign d0_w[52] = 4'h6;
    assign d0_w[53] = 4'h2;
    assign d0_w[54] = 4'h5;
    assign d0_w[55] = 4'hB;
    assign d0_w[56] = 4'h5;
    assign d0_w[57] = 4'hA;
    assign d0_w[58] = 4'h1;
    assign d0_w[59] = 4'hE;
    assign d0_w[60] = 4'h2;
    assign d0_w[61] = 4'h4;
    assign d0_w[62] = 4'hB;
    assign d0_w[63] = 4'hE;
    assign d0_w[64] = 4'h3;
    assign d0_w[65] = 4'hF;
    assign d0_w[66] = 4'hE;
    assign d0_w[67] = 4'hB;
    assign d0_w[68] = 4'hC;
    assign d0_w[69] = 4'h2;
    assign d0_w[70] = 4'h5;
    assign d0_w[71] = 4'hF;
    assign d0_w[72] = 4'h1;
    assign d0_w[73] = 4'hD;
    assign d0_w[74] = 4'h1;
    assign d0_w[75] = 4'h1;
    assign d0_w[76] = 4'h0;
    assign d0_w[77] = 4'hD;
    assign d0_w[78] = 4'hF;
    assign d0_w[79] = 4'hB;
    assign d0_w[80] = 4'h1;
    assign d0_w[81] = 4'hA;
    assign d0_w[82] = 4'hF;
    assign d0_w[83] = 4'hB;
    assign d0_w[84] = 4'hC;
    assign d0_w[85] = 4'h1;
    assign d0_w[86] = 4'hD;
    assign d0_w[87] = 4'hC;
    assign d0_w[88] = 4'hD;
    assign d0_w[89] = 4'hD;
    assign d0_w[90] = 4'h2;
    assign d0_w[91] = 4'h0;
    assign d0_w[92] = 4'h2;
    assign d0_w[93] = 4'hF;
    assign d0_w[94] = 4'hB;
    assign d0_w[95] = 4'h4;
    assign d0_w[96] = 4'h2;
    assign d0_w[97] = 4'h0;
    assign d0_w[98] = 4'hD;
    assign d0_w[99] = 4'hD;
    assign d0_w[100] = 4'h0;
    assign d0_w[101] = 4'hB;
    assign d0_w[102] = 4'hB;
    assign d0_w[103] = 4'h0;
    assign d0_w[104] = 4'h1;
    assign d0_w[105] = 4'h1;
    assign d0_w[106] = 4'h1;
    assign d0_w[107] = 4'hB;
    assign d0_w[108] = 4'h5;
    assign d0_w[109] = 4'h0;
    assign d0_w[110] = 4'h0;
    assign d0_w[111] = 4'hC;
    assign d0_w[112] = 4'h0;
    assign d0_w[113] = 4'h1;
    assign d0_w[114] = 4'h0;
    assign d0_w[115] = 4'hC;
    assign d0_w[116] = 4'h4;
    assign d0_w[117] = 4'hD;
    assign d0_w[118] = 4'hE;
    assign d0_w[119] = 4'h2;
    assign d0_w[120] = 4'hE;
    assign d0_w[121] = 4'h2;
    assign d0_w[122] = 4'hC;
    assign d0_w[123] = 4'hF;
    assign d0_w[124] = 4'h1;
    assign d0_w[125] = 4'h1;
    assign d0_w[126] = 4'h1;
    assign d0_w[127] = 4'hA;

    // --- layer0_b ---
    assign d0_b[0] = 4'h6;
    assign d0_b[1] = 4'h0;
    assign d0_b[2] = 4'h0;
    assign d0_b[3] = 4'h0;
    assign d0_b[4] = 4'hC;
    assign d0_b[5] = 4'h0;
    assign d0_b[6] = 4'hE;
    assign d0_b[7] = 4'h4;
    assign d0_b[8] = 4'h6;
    assign d0_b[9] = 4'h3;
    assign d0_b[10] = 4'hA;
    assign d0_b[11] = 4'h0;
    assign d0_b[12] = 4'hA;
    assign d0_b[13] = 4'h0;
    assign d0_b[14] = 4'h6;
    assign d0_b[15] = 4'h0;
    assign d0_b[16] = 4'h5;
    assign d0_b[17] = 4'hC;
    assign d0_b[18] = 4'h7;
    assign d0_b[19] = 4'h0;
    assign d0_b[20] = 4'hA;
    assign d0_b[21] = 4'h0;
    assign d0_b[22] = 4'h1;
    assign d0_b[23] = 4'h3;
    assign d0_b[24] = 4'h0;
    assign d0_b[25] = 4'h6;
    assign d0_b[26] = 4'h0;
    assign d0_b[27] = 4'h0;
    assign d0_b[28] = 4'h9;
    assign d0_b[29] = 4'hA;
    assign d0_b[30] = 4'hF;
    assign d0_b[31] = 4'h1;

    // --- layer1_w ---
    assign d1_w[0] = 4'h2;
    assign d1_w[1] = 4'h0;
    assign d1_w[2] = 4'h0;
    assign d1_w[3] = 4'hE;
    assign d1_w[4] = 4'h3;
    assign d1_w[5] = 4'h1;
    assign d1_w[6] = 4'h1;
    assign d1_w[7] = 4'h1;
    assign d1_w[8] = 4'h1;
    assign d1_w[9] = 4'hE;
    assign d1_w[10] = 4'h0;
    assign d1_w[11] = 4'h3;
    assign d1_w[12] = 4'h2;
    assign d1_w[13] = 4'hE;
    assign d1_w[14] = 4'hE;
    assign d1_w[15] = 4'h1;
    assign d1_w[16] = 4'h2;
    assign d1_w[17] = 4'hF;
    assign d1_w[18] = 4'h2;
    assign d1_w[19] = 4'hF;
    assign d1_w[20] = 4'h0;
    assign d1_w[21] = 4'hF;
    assign d1_w[22] = 4'hE;
    assign d1_w[23] = 4'hE;
    assign d1_w[24] = 4'hF;
    assign d1_w[25] = 4'h1;
    assign d1_w[26] = 4'hE;
    assign d1_w[27] = 4'h3;
    assign d1_w[28] = 4'hE;
    assign d1_w[29] = 4'hD;
    assign d1_w[30] = 4'hD;
    assign d1_w[31] = 4'h2;
    assign d1_w[32] = 4'hF;
    assign d1_w[33] = 4'h0;
    assign d1_w[34] = 4'h2;
    assign d1_w[35] = 4'hE;
    assign d1_w[36] = 4'hF;
    assign d1_w[37] = 4'hD;
    assign d1_w[38] = 4'hD;
    assign d1_w[39] = 4'hE;
    assign d1_w[40] = 4'h0;
    assign d1_w[41] = 4'h1;
    assign d1_w[42] = 4'hD;
    assign d1_w[43] = 4'h1;
    assign d1_w[44] = 4'hD;
    assign d1_w[45] = 4'h0;
    assign d1_w[46] = 4'h0;
    assign d1_w[47] = 4'hE;
    assign d1_w[48] = 4'hD;
    assign d1_w[49] = 4'hE;
    assign d1_w[50] = 4'hD;
    assign d1_w[51] = 4'hF;
    assign d1_w[52] = 4'hF;
    assign d1_w[53] = 4'h0;
    assign d1_w[54] = 4'h1;
    assign d1_w[55] = 4'hF;
    assign d1_w[56] = 4'h1;
    assign d1_w[57] = 4'hF;
    assign d1_w[58] = 4'h3;
    assign d1_w[59] = 4'h3;
    assign d1_w[60] = 4'h2;
    assign d1_w[61] = 4'hF;
    assign d1_w[62] = 4'hE;
    assign d1_w[63] = 4'h1;
    assign d1_w[64] = 4'h2;
    assign d1_w[65] = 4'h2;
    assign d1_w[66] = 4'hE;
    assign d1_w[67] = 4'h0;
    assign d1_w[68] = 4'h0;
    assign d1_w[69] = 4'h2;
    assign d1_w[70] = 4'hE;
    assign d1_w[71] = 4'hE;
    assign d1_w[72] = 4'hD;
    assign d1_w[73] = 4'h1;
    assign d1_w[74] = 4'h3;
    assign d1_w[75] = 4'hD;
    assign d1_w[76] = 4'hF;
    assign d1_w[77] = 4'hE;
    assign d1_w[78] = 4'h3;
    assign d1_w[79] = 4'hE;
    assign d1_w[80] = 4'hD;
    assign d1_w[81] = 4'h3;
    assign d1_w[82] = 4'hE;
    assign d1_w[83] = 4'h1;
    assign d1_w[84] = 4'hE;
    assign d1_w[85] = 4'hD;
    assign d1_w[86] = 4'hF;
    assign d1_w[87] = 4'h1;
    assign d1_w[88] = 4'h1;
    assign d1_w[89] = 4'h2;
    assign d1_w[90] = 4'hE;
    assign d1_w[91] = 4'h3;
    assign d1_w[92] = 4'h1;
    assign d1_w[93] = 4'h1;
    assign d1_w[94] = 4'h3;
    assign d1_w[95] = 4'h3;
    assign d1_w[96] = 4'hD;
    assign d1_w[97] = 4'h0;
    assign d1_w[98] = 4'hF;
    assign d1_w[99] = 4'h2;
    assign d1_w[100] = 4'h3;
    assign d1_w[101] = 4'h1;
    assign d1_w[102] = 4'h2;
    assign d1_w[103] = 4'hF;
    assign d1_w[104] = 4'hD;
    assign d1_w[105] = 4'hE;
    assign d1_w[106] = 4'h1;
    assign d1_w[107] = 4'h1;
    assign d1_w[108] = 4'h3;
    assign d1_w[109] = 4'h0;
    assign d1_w[110] = 4'hD;
    assign d1_w[111] = 4'hE;
    assign d1_w[112] = 4'h3;
    assign d1_w[113] = 4'hF;
    assign d1_w[114] = 4'h3;
    assign d1_w[115] = 4'h1;
    assign d1_w[116] = 4'h0;
    assign d1_w[117] = 4'h1;
    assign d1_w[118] = 4'h0;
    assign d1_w[119] = 4'h3;
    assign d1_w[120] = 4'hF;
    assign d1_w[121] = 4'hF;
    assign d1_w[122] = 4'h0;
    assign d1_w[123] = 4'h0;
    assign d1_w[124] = 4'hF;
    assign d1_w[125] = 4'h3;
    assign d1_w[126] = 4'hE;
    assign d1_w[127] = 4'h2;
    assign d1_w[128] = 4'h0;
    assign d1_w[129] = 4'h1;
    assign d1_w[130] = 4'hE;
    assign d1_w[131] = 4'h1;
    assign d1_w[132] = 4'h0;
    assign d1_w[133] = 4'hD;
    assign d1_w[134] = 4'h1;
    assign d1_w[135] = 4'h0;
    assign d1_w[136] = 4'hF;
    assign d1_w[137] = 4'h2;
    assign d1_w[138] = 4'h1;
    assign d1_w[139] = 4'h2;
    assign d1_w[140] = 4'hE;
    assign d1_w[141] = 4'h2;
    assign d1_w[142] = 4'h2;
    assign d1_w[143] = 4'h3;
    assign d1_w[144] = 4'h2;
    assign d1_w[145] = 4'hE;
    assign d1_w[146] = 4'hE;
    assign d1_w[147] = 4'hE;
    assign d1_w[148] = 4'h2;
    assign d1_w[149] = 4'h1;
    assign d1_w[150] = 4'h2;
    assign d1_w[151] = 4'h1;
    assign d1_w[152] = 4'h0;
    assign d1_w[153] = 4'h0;
    assign d1_w[154] = 4'h2;
    assign d1_w[155] = 4'h0;
    assign d1_w[156] = 4'hC;
    assign d1_w[157] = 4'hD;
    assign d1_w[158] = 4'hD;
    assign d1_w[159] = 4'hF;
    assign d1_w[160] = 4'hF;
    assign d1_w[161] = 4'h0;
    assign d1_w[162] = 4'hF;
    assign d1_w[163] = 4'h1;
    assign d1_w[164] = 4'h2;
    assign d1_w[165] = 4'hD;
    assign d1_w[166] = 4'h1;
    assign d1_w[167] = 4'h2;
    assign d1_w[168] = 4'h0;
    assign d1_w[169] = 4'h3;
    assign d1_w[170] = 4'h1;
    assign d1_w[171] = 4'hD;
    assign d1_w[172] = 4'h2;
    assign d1_w[173] = 4'h0;
    assign d1_w[174] = 4'h3;
    assign d1_w[175] = 4'h0;
    assign d1_w[176] = 4'hF;
    assign d1_w[177] = 4'h1;
    assign d1_w[178] = 4'hC;
    assign d1_w[179] = 4'h1;
    assign d1_w[180] = 4'h2;
    assign d1_w[181] = 4'hD;
    assign d1_w[182] = 4'h2;
    assign d1_w[183] = 4'hF;
    assign d1_w[184] = 4'h0;
    assign d1_w[185] = 4'h0;
    assign d1_w[186] = 4'hF;
    assign d1_w[187] = 4'h1;
    assign d1_w[188] = 4'h3;
    assign d1_w[189] = 4'hD;
    assign d1_w[190] = 4'h1;
    assign d1_w[191] = 4'h3;
    assign d1_w[192] = 4'h1;
    assign d1_w[193] = 4'hF;
    assign d1_w[194] = 4'hF;
    assign d1_w[195] = 4'hE;
    assign d1_w[196] = 4'h1;
    assign d1_w[197] = 4'h3;
    assign d1_w[198] = 4'h2;
    assign d1_w[199] = 4'hD;
    assign d1_w[200] = 4'h1;
    assign d1_w[201] = 4'hE;
    assign d1_w[202] = 4'h0;
    assign d1_w[203] = 4'h1;
    assign d1_w[204] = 4'h2;
    assign d1_w[205] = 4'h1;
    assign d1_w[206] = 4'hE;
    assign d1_w[207] = 4'h2;
    assign d1_w[208] = 4'hF;
    assign d1_w[209] = 4'h0;
    assign d1_w[210] = 4'hF;
    assign d1_w[211] = 4'h2;
    assign d1_w[212] = 4'h0;
    assign d1_w[213] = 4'h4;
    assign d1_w[214] = 4'h0;
    assign d1_w[215] = 4'hD;
    assign d1_w[216] = 4'hE;
    assign d1_w[217] = 4'hE;
    assign d1_w[218] = 4'hE;
    assign d1_w[219] = 4'h1;
    assign d1_w[220] = 4'h0;
    assign d1_w[221] = 4'h0;
    assign d1_w[222] = 4'hD;
    assign d1_w[223] = 4'h1;
    assign d1_w[224] = 4'h3;
    assign d1_w[225] = 4'h3;
    assign d1_w[226] = 4'hF;
    assign d1_w[227] = 4'h1;
    assign d1_w[228] = 4'h1;
    assign d1_w[229] = 4'h0;
    assign d1_w[230] = 4'h1;
    assign d1_w[231] = 4'hC;
    assign d1_w[232] = 4'hE;
    assign d1_w[233] = 4'h1;
    assign d1_w[234] = 4'hF;
    assign d1_w[235] = 4'h2;
    assign d1_w[236] = 4'h0;
    assign d1_w[237] = 4'hD;
    assign d1_w[238] = 4'h3;
    assign d1_w[239] = 4'hE;
    assign d1_w[240] = 4'h0;
    assign d1_w[241] = 4'h3;
    assign d1_w[242] = 4'h1;
    assign d1_w[243] = 4'h0;
    assign d1_w[244] = 4'hF;
    assign d1_w[245] = 4'h2;
    assign d1_w[246] = 4'hD;
    assign d1_w[247] = 4'h0;
    assign d1_w[248] = 4'h3;
    assign d1_w[249] = 4'hF;
    assign d1_w[250] = 4'h2;
    assign d1_w[251] = 4'h1;
    assign d1_w[252] = 4'hE;
    assign d1_w[253] = 4'h3;
    assign d1_w[254] = 4'hD;
    assign d1_w[255] = 4'hE;
    assign d1_w[256] = 4'h0;
    assign d1_w[257] = 4'h0;
    assign d1_w[258] = 4'h2;
    assign d1_w[259] = 4'h0;
    assign d1_w[260] = 4'hE;
    assign d1_w[261] = 4'h0;
    assign d1_w[262] = 4'h0;
    assign d1_w[263] = 4'hF;
    assign d1_w[264] = 4'hD;
    assign d1_w[265] = 4'h1;
    assign d1_w[266] = 4'h0;
    assign d1_w[267] = 4'hD;
    assign d1_w[268] = 4'h0;
    assign d1_w[269] = 4'h1;
    assign d1_w[270] = 4'hF;
    assign d1_w[271] = 4'hD;
    assign d1_w[272] = 4'h0;
    assign d1_w[273] = 4'h1;
    assign d1_w[274] = 4'hF;
    assign d1_w[275] = 4'h0;
    assign d1_w[276] = 4'hE;
    assign d1_w[277] = 4'hE;
    assign d1_w[278] = 4'h1;
    assign d1_w[279] = 4'hE;
    assign d1_w[280] = 4'hD;
    assign d1_w[281] = 4'hF;
    assign d1_w[282] = 4'h1;
    assign d1_w[283] = 4'h3;
    assign d1_w[284] = 4'h0;
    assign d1_w[285] = 4'h2;
    assign d1_w[286] = 4'hD;
    assign d1_w[287] = 4'hF;
    assign d1_w[288] = 4'h2;
    assign d1_w[289] = 4'h2;
    assign d1_w[290] = 4'h0;
    assign d1_w[291] = 4'h3;
    assign d1_w[292] = 4'hD;
    assign d1_w[293] = 4'hF;
    assign d1_w[294] = 4'h0;
    assign d1_w[295] = 4'hE;
    assign d1_w[296] = 4'h1;
    assign d1_w[297] = 4'hD;
    assign d1_w[298] = 4'h1;
    assign d1_w[299] = 4'h1;
    assign d1_w[300] = 4'hF;
    assign d1_w[301] = 4'hE;
    assign d1_w[302] = 4'h1;
    assign d1_w[303] = 4'hF;
    assign d1_w[304] = 4'h1;
    assign d1_w[305] = 4'h2;
    assign d1_w[306] = 4'h1;
    assign d1_w[307] = 4'hF;
    assign d1_w[308] = 4'h0;
    assign d1_w[309] = 4'hF;
    assign d1_w[310] = 4'hF;
    assign d1_w[311] = 4'hF;
    assign d1_w[312] = 4'h3;
    assign d1_w[313] = 4'h3;
    assign d1_w[314] = 4'h1;
    assign d1_w[315] = 4'hE;
    assign d1_w[316] = 4'hF;
    assign d1_w[317] = 4'h0;
    assign d1_w[318] = 4'hD;
    assign d1_w[319] = 4'hD;
    assign d1_w[320] = 4'h2;
    assign d1_w[321] = 4'hF;
    assign d1_w[322] = 4'h3;
    assign d1_w[323] = 4'hF;
    assign d1_w[324] = 4'h2;
    assign d1_w[325] = 4'hF;
    assign d1_w[326] = 4'hF;
    assign d1_w[327] = 4'hC;
    assign d1_w[328] = 4'h2;
    assign d1_w[329] = 4'h0;
    assign d1_w[330] = 4'hE;
    assign d1_w[331] = 4'hF;
    assign d1_w[332] = 4'hE;
    assign d1_w[333] = 4'h0;
    assign d1_w[334] = 4'h3;
    assign d1_w[335] = 4'h1;
    assign d1_w[336] = 4'h0;
    assign d1_w[337] = 4'h0;
    assign d1_w[338] = 4'hF;
    assign d1_w[339] = 4'h0;
    assign d1_w[340] = 4'h0;
    assign d1_w[341] = 4'hD;
    assign d1_w[342] = 4'hF;
    assign d1_w[343] = 4'hD;
    assign d1_w[344] = 4'h0;
    assign d1_w[345] = 4'hE;
    assign d1_w[346] = 4'h2;
    assign d1_w[347] = 4'hE;
    assign d1_w[348] = 4'hD;
    assign d1_w[349] = 4'h0;
    assign d1_w[350] = 4'h1;
    assign d1_w[351] = 4'hF;
    assign d1_w[352] = 4'h2;
    assign d1_w[353] = 4'h1;
    assign d1_w[354] = 4'hE;
    assign d1_w[355] = 4'h3;
    assign d1_w[356] = 4'h0;
    assign d1_w[357] = 4'h2;
    assign d1_w[358] = 4'hE;
    assign d1_w[359] = 4'hD;
    assign d1_w[360] = 4'h3;
    assign d1_w[361] = 4'hE;
    assign d1_w[362] = 4'h0;
    assign d1_w[363] = 4'hF;
    assign d1_w[364] = 4'h2;
    assign d1_w[365] = 4'hF;
    assign d1_w[366] = 4'hF;
    assign d1_w[367] = 4'h0;
    assign d1_w[368] = 4'h1;
    assign d1_w[369] = 4'hD;
    assign d1_w[370] = 4'hD;
    assign d1_w[371] = 4'h2;
    assign d1_w[372] = 4'hE;
    assign d1_w[373] = 4'hD;
    assign d1_w[374] = 4'h1;
    assign d1_w[375] = 4'hE;
    assign d1_w[376] = 4'h2;
    assign d1_w[377] = 4'hF;
    assign d1_w[378] = 4'h0;
    assign d1_w[379] = 4'hE;
    assign d1_w[380] = 4'h0;
    assign d1_w[381] = 4'h1;
    assign d1_w[382] = 4'hE;
    assign d1_w[383] = 4'hE;
    assign d1_w[384] = 4'hF;
    assign d1_w[385] = 4'h2;
    assign d1_w[386] = 4'h0;
    assign d1_w[387] = 4'hE;
    assign d1_w[388] = 4'hE;
    assign d1_w[389] = 4'h1;
    assign d1_w[390] = 4'h2;
    assign d1_w[391] = 4'h0;
    assign d1_w[392] = 4'hF;
    assign d1_w[393] = 4'h3;
    assign d1_w[394] = 4'hF;
    assign d1_w[395] = 4'hE;
    assign d1_w[396] = 4'hD;
    assign d1_w[397] = 4'hD;
    assign d1_w[398] = 4'h3;
    assign d1_w[399] = 4'hD;
    assign d1_w[400] = 4'hD;
    assign d1_w[401] = 4'hE;
    assign d1_w[402] = 4'hE;
    assign d1_w[403] = 4'h1;
    assign d1_w[404] = 4'hD;
    assign d1_w[405] = 4'h1;
    assign d1_w[406] = 4'hF;
    assign d1_w[407] = 4'hE;
    assign d1_w[408] = 4'hE;
    assign d1_w[409] = 4'h0;
    assign d1_w[410] = 4'h1;
    assign d1_w[411] = 4'hE;
    assign d1_w[412] = 4'h3;
    assign d1_w[413] = 4'hF;
    assign d1_w[414] = 4'h2;
    assign d1_w[415] = 4'hD;
    assign d1_w[416] = 4'h2;
    assign d1_w[417] = 4'hF;
    assign d1_w[418] = 4'h0;
    assign d1_w[419] = 4'h0;
    assign d1_w[420] = 4'hF;
    assign d1_w[421] = 4'hE;
    assign d1_w[422] = 4'h0;
    assign d1_w[423] = 4'hF;
    assign d1_w[424] = 4'hE;
    assign d1_w[425] = 4'h0;
    assign d1_w[426] = 4'hE;
    assign d1_w[427] = 4'h2;
    assign d1_w[428] = 4'h2;
    assign d1_w[429] = 4'h0;
    assign d1_w[430] = 4'hE;
    assign d1_w[431] = 4'h0;
    assign d1_w[432] = 4'hD;
    assign d1_w[433] = 4'h0;
    assign d1_w[434] = 4'hD;
    assign d1_w[435] = 4'hD;
    assign d1_w[436] = 4'h2;
    assign d1_w[437] = 4'hF;
    assign d1_w[438] = 4'h1;
    assign d1_w[439] = 4'h3;
    assign d1_w[440] = 4'h1;
    assign d1_w[441] = 4'hF;
    assign d1_w[442] = 4'hF;
    assign d1_w[443] = 4'hD;
    assign d1_w[444] = 4'h2;
    assign d1_w[445] = 4'h1;
    assign d1_w[446] = 4'hF;
    assign d1_w[447] = 4'h0;
    assign d1_w[448] = 4'h4;
    assign d1_w[449] = 4'hA;
    assign d1_w[450] = 4'h6;
    assign d1_w[451] = 4'h3;
    assign d1_w[452] = 4'h0;
    assign d1_w[453] = 4'hD;
    assign d1_w[454] = 4'hE;
    assign d1_w[455] = 4'hD;
    assign d1_w[456] = 4'hE;
    assign d1_w[457] = 4'hE;
    assign d1_w[458] = 4'h0;
    assign d1_w[459] = 4'hE;
    assign d1_w[460] = 4'h1;
    assign d1_w[461] = 4'hD;
    assign d1_w[462] = 4'hB;
    assign d1_w[463] = 4'hF;
    assign d1_w[464] = 4'hB;
    assign d1_w[465] = 4'h5;
    assign d1_w[466] = 4'h2;
    assign d1_w[467] = 4'hE;
    assign d1_w[468] = 4'hF;
    assign d1_w[469] = 4'h0;
    assign d1_w[470] = 4'hF;
    assign d1_w[471] = 4'hE;
    assign d1_w[472] = 4'hE;
    assign d1_w[473] = 4'h6;
    assign d1_w[474] = 4'hF;
    assign d1_w[475] = 4'h7;
    assign d1_w[476] = 4'h1;
    assign d1_w[477] = 4'hD;
    assign d1_w[478] = 4'h2;
    assign d1_w[479] = 4'h1;
    assign d1_w[480] = 4'h2;
    assign d1_w[481] = 4'h1;
    assign d1_w[482] = 4'hE;
    assign d1_w[483] = 4'hD;
    assign d1_w[484] = 4'h0;
    assign d1_w[485] = 4'h0;
    assign d1_w[486] = 4'h3;
    assign d1_w[487] = 4'h0;
    assign d1_w[488] = 4'h0;
    assign d1_w[489] = 4'h1;
    assign d1_w[490] = 4'h0;
    assign d1_w[491] = 4'h1;
    assign d1_w[492] = 4'h1;
    assign d1_w[493] = 4'hD;
    assign d1_w[494] = 4'hE;
    assign d1_w[495] = 4'hE;
    assign d1_w[496] = 4'h3;
    assign d1_w[497] = 4'hD;
    assign d1_w[498] = 4'h1;
    assign d1_w[499] = 4'hE;
    assign d1_w[500] = 4'h1;
    assign d1_w[501] = 4'hD;
    assign d1_w[502] = 4'hD;
    assign d1_w[503] = 4'hD;
    assign d1_w[504] = 4'h0;
    assign d1_w[505] = 4'hE;
    assign d1_w[506] = 4'h2;
    assign d1_w[507] = 4'h0;
    assign d1_w[508] = 4'hE;
    assign d1_w[509] = 4'h0;
    assign d1_w[510] = 4'hF;
    assign d1_w[511] = 4'h1;
    assign d1_w[512] = 4'h2;
    assign d1_w[513] = 4'h3;
    assign d1_w[514] = 4'hE;
    assign d1_w[515] = 4'h3;
    assign d1_w[516] = 4'h3;
    assign d1_w[517] = 4'h0;
    assign d1_w[518] = 4'hF;
    assign d1_w[519] = 4'h1;
    assign d1_w[520] = 4'hF;
    assign d1_w[521] = 4'h3;
    assign d1_w[522] = 4'h0;
    assign d1_w[523] = 4'h0;
    assign d1_w[524] = 4'hD;
    assign d1_w[525] = 4'h1;
    assign d1_w[526] = 4'h2;
    assign d1_w[527] = 4'hF;
    assign d1_w[528] = 4'h1;
    assign d1_w[529] = 4'h3;
    assign d1_w[530] = 4'h3;
    assign d1_w[531] = 4'hD;
    assign d1_w[532] = 4'hF;
    assign d1_w[533] = 4'hE;
    assign d1_w[534] = 4'h1;
    assign d1_w[535] = 4'h0;
    assign d1_w[536] = 4'hD;
    assign d1_w[537] = 4'hF;
    assign d1_w[538] = 4'hE;
    assign d1_w[539] = 4'h1;
    assign d1_w[540] = 4'h1;
    assign d1_w[541] = 4'hE;
    assign d1_w[542] = 4'hF;
    assign d1_w[543] = 4'hD;
    assign d1_w[544] = 4'hE;
    assign d1_w[545] = 4'h3;
    assign d1_w[546] = 4'hE;
    assign d1_w[547] = 4'h2;
    assign d1_w[548] = 4'h0;
    assign d1_w[549] = 4'h0;
    assign d1_w[550] = 4'h1;
    assign d1_w[551] = 4'h3;
    assign d1_w[552] = 4'h2;
    assign d1_w[553] = 4'h2;
    assign d1_w[554] = 4'hF;
    assign d1_w[555] = 4'h2;
    assign d1_w[556] = 4'h3;
    assign d1_w[557] = 4'h2;
    assign d1_w[558] = 4'h2;
    assign d1_w[559] = 4'h0;
    assign d1_w[560] = 4'h2;
    assign d1_w[561] = 4'hE;
    assign d1_w[562] = 4'h2;
    assign d1_w[563] = 4'h0;
    assign d1_w[564] = 4'h4;
    assign d1_w[565] = 4'hF;
    assign d1_w[566] = 4'hD;
    assign d1_w[567] = 4'hE;
    assign d1_w[568] = 4'h0;
    assign d1_w[569] = 4'h2;
    assign d1_w[570] = 4'hD;
    assign d1_w[571] = 4'hF;
    assign d1_w[572] = 4'h0;
    assign d1_w[573] = 4'h2;
    assign d1_w[574] = 4'h2;
    assign d1_w[575] = 4'h1;
    assign d1_w[576] = 4'hF;
    assign d1_w[577] = 4'hF;
    assign d1_w[578] = 4'h2;
    assign d1_w[579] = 4'h1;
    assign d1_w[580] = 4'hE;
    assign d1_w[581] = 4'h2;
    assign d1_w[582] = 4'hD;
    assign d1_w[583] = 4'h1;
    assign d1_w[584] = 4'h1;
    assign d1_w[585] = 4'h1;
    assign d1_w[586] = 4'h0;
    assign d1_w[587] = 4'h3;
    assign d1_w[588] = 4'hE;
    assign d1_w[589] = 4'h2;
    assign d1_w[590] = 4'h1;
    assign d1_w[591] = 4'h4;
    assign d1_w[592] = 4'hF;
    assign d1_w[593] = 4'h3;
    assign d1_w[594] = 4'h4;
    assign d1_w[595] = 4'h0;
    assign d1_w[596] = 4'h3;
    assign d1_w[597] = 4'h3;
    assign d1_w[598] = 4'hE;
    assign d1_w[599] = 4'hD;
    assign d1_w[600] = 4'hD;
    assign d1_w[601] = 4'hE;
    assign d1_w[602] = 4'hD;
    assign d1_w[603] = 4'h3;
    assign d1_w[604] = 4'hE;
    assign d1_w[605] = 4'hD;
    assign d1_w[606] = 4'h1;
    assign d1_w[607] = 4'h1;
    assign d1_w[608] = 4'h2;
    assign d1_w[609] = 4'h2;
    assign d1_w[610] = 4'hF;
    assign d1_w[611] = 4'h0;
    assign d1_w[612] = 4'h3;
    assign d1_w[613] = 4'hF;
    assign d1_w[614] = 4'h2;
    assign d1_w[615] = 4'h2;
    assign d1_w[616] = 4'h3;
    assign d1_w[617] = 4'h1;
    assign d1_w[618] = 4'hF;
    assign d1_w[619] = 4'h1;
    assign d1_w[620] = 4'h0;
    assign d1_w[621] = 4'hE;
    assign d1_w[622] = 4'h2;
    assign d1_w[623] = 4'hE;
    assign d1_w[624] = 4'h0;
    assign d1_w[625] = 4'h0;
    assign d1_w[626] = 4'hE;
    assign d1_w[627] = 4'h3;
    assign d1_w[628] = 4'h3;
    assign d1_w[629] = 4'h3;
    assign d1_w[630] = 4'h3;
    assign d1_w[631] = 4'hD;
    assign d1_w[632] = 4'h3;
    assign d1_w[633] = 4'hF;
    assign d1_w[634] = 4'hD;
    assign d1_w[635] = 4'h0;
    assign d1_w[636] = 4'h0;
    assign d1_w[637] = 4'h2;
    assign d1_w[638] = 4'h3;
    assign d1_w[639] = 4'h0;
    assign d1_w[640] = 4'hF;
    assign d1_w[641] = 4'hD;
    assign d1_w[642] = 4'h1;
    assign d1_w[643] = 4'h0;
    assign d1_w[644] = 4'h0;
    assign d1_w[645] = 4'h0;
    assign d1_w[646] = 4'h1;
    assign d1_w[647] = 4'hD;
    assign d1_w[648] = 4'h2;
    assign d1_w[649] = 4'hD;
    assign d1_w[650] = 4'hF;
    assign d1_w[651] = 4'h1;
    assign d1_w[652] = 4'hD;
    assign d1_w[653] = 4'h1;
    assign d1_w[654] = 4'h0;
    assign d1_w[655] = 4'hE;
    assign d1_w[656] = 4'h2;
    assign d1_w[657] = 4'hD;
    assign d1_w[658] = 4'hF;
    assign d1_w[659] = 4'hF;
    assign d1_w[660] = 4'hF;
    assign d1_w[661] = 4'h2;
    assign d1_w[662] = 4'h0;
    assign d1_w[663] = 4'hD;
    assign d1_w[664] = 4'hF;
    assign d1_w[665] = 4'hF;
    assign d1_w[666] = 4'h3;
    assign d1_w[667] = 4'hF;
    assign d1_w[668] = 4'hD;
    assign d1_w[669] = 4'h1;
    assign d1_w[670] = 4'h0;
    assign d1_w[671] = 4'hE;
    assign d1_w[672] = 4'hF;
    assign d1_w[673] = 4'h1;
    assign d1_w[674] = 4'hD;
    assign d1_w[675] = 4'hF;
    assign d1_w[676] = 4'hE;
    assign d1_w[677] = 4'h1;
    assign d1_w[678] = 4'h2;
    assign d1_w[679] = 4'h2;
    assign d1_w[680] = 4'h3;
    assign d1_w[681] = 4'h2;
    assign d1_w[682] = 4'h3;
    assign d1_w[683] = 4'hE;
    assign d1_w[684] = 4'h1;
    assign d1_w[685] = 4'hF;
    assign d1_w[686] = 4'hE;
    assign d1_w[687] = 4'h0;
    assign d1_w[688] = 4'hE;
    assign d1_w[689] = 4'h2;
    assign d1_w[690] = 4'h2;
    assign d1_w[691] = 4'hD;
    assign d1_w[692] = 4'hF;
    assign d1_w[693] = 4'hE;
    assign d1_w[694] = 4'h2;
    assign d1_w[695] = 4'hD;
    assign d1_w[696] = 4'hE;
    assign d1_w[697] = 4'h0;
    assign d1_w[698] = 4'h2;
    assign d1_w[699] = 4'hE;
    assign d1_w[700] = 4'h2;
    assign d1_w[701] = 4'h2;
    assign d1_w[702] = 4'hD;
    assign d1_w[703] = 4'hF;
    assign d1_w[704] = 4'h1;
    assign d1_w[705] = 4'h1;
    assign d1_w[706] = 4'hE;
    assign d1_w[707] = 4'h1;
    assign d1_w[708] = 4'h3;
    assign d1_w[709] = 4'h1;
    assign d1_w[710] = 4'hE;
    assign d1_w[711] = 4'h2;
    assign d1_w[712] = 4'h0;
    assign d1_w[713] = 4'hE;
    assign d1_w[714] = 4'h2;
    assign d1_w[715] = 4'hF;
    assign d1_w[716] = 4'hD;
    assign d1_w[717] = 4'h0;
    assign d1_w[718] = 4'hE;
    assign d1_w[719] = 4'h5;
    assign d1_w[720] = 4'h1;
    assign d1_w[721] = 4'h2;
    assign d1_w[722] = 4'hF;
    assign d1_w[723] = 4'h2;
    assign d1_w[724] = 4'h2;
    assign d1_w[725] = 4'hD;
    assign d1_w[726] = 4'h1;
    assign d1_w[727] = 4'h2;
    assign d1_w[728] = 4'h2;
    assign d1_w[729] = 4'h2;
    assign d1_w[730] = 4'h1;
    assign d1_w[731] = 4'hF;
    assign d1_w[732] = 4'h2;
    assign d1_w[733] = 4'hF;
    assign d1_w[734] = 4'hF;
    assign d1_w[735] = 4'h2;
    assign d1_w[736] = 4'hF;
    assign d1_w[737] = 4'h1;
    assign d1_w[738] = 4'h0;
    assign d1_w[739] = 4'hE;
    assign d1_w[740] = 4'hF;
    assign d1_w[741] = 4'hE;
    assign d1_w[742] = 4'hE;
    assign d1_w[743] = 4'hD;
    assign d1_w[744] = 4'h1;
    assign d1_w[745] = 4'hD;
    assign d1_w[746] = 4'h2;
    assign d1_w[747] = 4'h1;
    assign d1_w[748] = 4'h1;
    assign d1_w[749] = 4'hF;
    assign d1_w[750] = 4'h2;
    assign d1_w[751] = 4'h1;
    assign d1_w[752] = 4'h0;
    assign d1_w[753] = 4'h2;
    assign d1_w[754] = 4'h2;
    assign d1_w[755] = 4'hF;
    assign d1_w[756] = 4'h0;
    assign d1_w[757] = 4'h0;
    assign d1_w[758] = 4'h1;
    assign d1_w[759] = 4'h2;
    assign d1_w[760] = 4'h3;
    assign d1_w[761] = 4'hF;
    assign d1_w[762] = 4'h2;
    assign d1_w[763] = 4'h1;
    assign d1_w[764] = 4'hD;
    assign d1_w[765] = 4'h1;
    assign d1_w[766] = 4'h2;
    assign d1_w[767] = 4'hD;
    assign d1_w[768] = 4'hF;
    assign d1_w[769] = 4'h1;
    assign d1_w[770] = 4'h2;
    assign d1_w[771] = 4'h2;
    assign d1_w[772] = 4'h2;
    assign d1_w[773] = 4'h1;
    assign d1_w[774] = 4'h3;
    assign d1_w[775] = 4'h1;
    assign d1_w[776] = 4'hE;
    assign d1_w[777] = 4'hF;
    assign d1_w[778] = 4'hE;
    assign d1_w[779] = 4'hD;
    assign d1_w[780] = 4'h1;
    assign d1_w[781] = 4'h2;
    assign d1_w[782] = 4'hF;
    assign d1_w[783] = 4'h2;
    assign d1_w[784] = 4'h2;
    assign d1_w[785] = 4'hE;
    assign d1_w[786] = 4'hE;
    assign d1_w[787] = 4'h3;
    assign d1_w[788] = 4'h2;
    assign d1_w[789] = 4'hE;
    assign d1_w[790] = 4'h3;
    assign d1_w[791] = 4'h0;
    assign d1_w[792] = 4'hF;
    assign d1_w[793] = 4'hF;
    assign d1_w[794] = 4'h3;
    assign d1_w[795] = 4'hD;
    assign d1_w[796] = 4'hF;
    assign d1_w[797] = 4'hD;
    assign d1_w[798] = 4'hE;
    assign d1_w[799] = 4'h1;
    assign d1_w[800] = 4'h2;
    assign d1_w[801] = 4'h0;
    assign d1_w[802] = 4'h2;
    assign d1_w[803] = 4'h0;
    assign d1_w[804] = 4'h1;
    assign d1_w[805] = 4'hC;
    assign d1_w[806] = 4'hE;
    assign d1_w[807] = 4'h0;
    assign d1_w[808] = 4'hD;
    assign d1_w[809] = 4'h1;
    assign d1_w[810] = 4'h0;
    assign d1_w[811] = 4'hE;
    assign d1_w[812] = 4'h0;
    assign d1_w[813] = 4'hD;
    assign d1_w[814] = 4'hC;
    assign d1_w[815] = 4'h1;
    assign d1_w[816] = 4'h1;
    assign d1_w[817] = 4'h4;
    assign d1_w[818] = 4'h5;
    assign d1_w[819] = 4'h2;
    assign d1_w[820] = 4'h2;
    assign d1_w[821] = 4'hE;
    assign d1_w[822] = 4'hF;
    assign d1_w[823] = 4'h3;
    assign d1_w[824] = 4'hF;
    assign d1_w[825] = 4'h2;
    assign d1_w[826] = 4'hD;
    assign d1_w[827] = 4'h5;
    assign d1_w[828] = 4'h0;
    assign d1_w[829] = 4'h1;
    assign d1_w[830] = 4'hD;
    assign d1_w[831] = 4'h1;
    assign d1_w[832] = 4'h0;
    assign d1_w[833] = 4'h0;
    assign d1_w[834] = 4'hF;
    assign d1_w[835] = 4'h2;
    assign d1_w[836] = 4'h0;
    assign d1_w[837] = 4'h3;
    assign d1_w[838] = 4'hE;
    assign d1_w[839] = 4'h1;
    assign d1_w[840] = 4'h1;
    assign d1_w[841] = 4'h1;
    assign d1_w[842] = 4'hD;
    assign d1_w[843] = 4'h2;
    assign d1_w[844] = 4'h0;
    assign d1_w[845] = 4'hF;
    assign d1_w[846] = 4'h2;
    assign d1_w[847] = 4'hE;
    assign d1_w[848] = 4'hD;
    assign d1_w[849] = 4'hF;
    assign d1_w[850] = 4'h3;
    assign d1_w[851] = 4'hF;
    assign d1_w[852] = 4'h2;
    assign d1_w[853] = 4'hD;
    assign d1_w[854] = 4'h2;
    assign d1_w[855] = 4'hE;
    assign d1_w[856] = 4'hE;
    assign d1_w[857] = 4'hE;
    assign d1_w[858] = 4'hF;
    assign d1_w[859] = 4'h0;
    assign d1_w[860] = 4'hF;
    assign d1_w[861] = 4'h0;
    assign d1_w[862] = 4'h2;
    assign d1_w[863] = 4'hF;
    assign d1_w[864] = 4'hF;
    assign d1_w[865] = 4'hE;
    assign d1_w[866] = 4'hF;
    assign d1_w[867] = 4'hE;
    assign d1_w[868] = 4'hE;
    assign d1_w[869] = 4'hF;
    assign d1_w[870] = 4'h2;
    assign d1_w[871] = 4'hF;
    assign d1_w[872] = 4'h0;
    assign d1_w[873] = 4'h2;
    assign d1_w[874] = 4'hF;
    assign d1_w[875] = 4'hF;
    assign d1_w[876] = 4'h3;
    assign d1_w[877] = 4'h0;
    assign d1_w[878] = 4'hE;
    assign d1_w[879] = 4'h0;
    assign d1_w[880] = 4'hD;
    assign d1_w[881] = 4'hE;
    assign d1_w[882] = 4'hF;
    assign d1_w[883] = 4'hF;
    assign d1_w[884] = 4'hD;
    assign d1_w[885] = 4'h4;
    assign d1_w[886] = 4'h1;
    assign d1_w[887] = 4'hE;
    assign d1_w[888] = 4'h0;
    assign d1_w[889] = 4'h2;
    assign d1_w[890] = 4'hE;
    assign d1_w[891] = 4'h1;
    assign d1_w[892] = 4'h1;
    assign d1_w[893] = 4'h1;
    assign d1_w[894] = 4'h1;
    assign d1_w[895] = 4'hF;
    assign d1_w[896] = 4'hC;
    assign d1_w[897] = 4'h1;
    assign d1_w[898] = 4'h1;
    assign d1_w[899] = 4'hF;
    assign d1_w[900] = 4'h3;
    assign d1_w[901] = 4'h2;
    assign d1_w[902] = 4'h2;
    assign d1_w[903] = 4'h1;
    assign d1_w[904] = 4'hD;
    assign d1_w[905] = 4'h3;
    assign d1_w[906] = 4'h1;
    assign d1_w[907] = 4'hE;
    assign d1_w[908] = 4'hC;
    assign d1_w[909] = 4'hF;
    assign d1_w[910] = 4'h2;
    assign d1_w[911] = 4'hF;
    assign d1_w[912] = 4'h1;
    assign d1_w[913] = 4'h1;
    assign d1_w[914] = 4'hF;
    assign d1_w[915] = 4'h2;
    assign d1_w[916] = 4'h1;
    assign d1_w[917] = 4'h1;
    assign d1_w[918] = 4'h1;
    assign d1_w[919] = 4'h2;
    assign d1_w[920] = 4'hE;
    assign d1_w[921] = 4'hD;
    assign d1_w[922] = 4'h3;
    assign d1_w[923] = 4'hD;
    assign d1_w[924] = 4'h2;
    assign d1_w[925] = 4'hF;
    assign d1_w[926] = 4'hE;
    assign d1_w[927] = 4'hF;
    assign d1_w[928] = 4'h1;
    assign d1_w[929] = 4'hF;
    assign d1_w[930] = 4'hF;
    assign d1_w[931] = 4'h0;
    assign d1_w[932] = 4'hF;
    assign d1_w[933] = 4'h1;
    assign d1_w[934] = 4'h0;
    assign d1_w[935] = 4'hF;
    assign d1_w[936] = 4'h0;
    assign d1_w[937] = 4'h3;
    assign d1_w[938] = 4'hD;
    assign d1_w[939] = 4'h2;
    assign d1_w[940] = 4'hE;
    assign d1_w[941] = 4'h1;
    assign d1_w[942] = 4'hE;
    assign d1_w[943] = 4'h1;
    assign d1_w[944] = 4'h2;
    assign d1_w[945] = 4'hC;
    assign d1_w[946] = 4'hF;
    assign d1_w[947] = 4'hF;
    assign d1_w[948] = 4'h0;
    assign d1_w[949] = 4'hE;
    assign d1_w[950] = 4'h1;
    assign d1_w[951] = 4'h1;
    assign d1_w[952] = 4'hE;
    assign d1_w[953] = 4'hF;
    assign d1_w[954] = 4'h1;
    assign d1_w[955] = 4'hE;
    assign d1_w[956] = 4'h0;
    assign d1_w[957] = 4'h0;
    assign d1_w[958] = 4'h0;
    assign d1_w[959] = 4'hE;
    assign d1_w[960] = 4'hE;
    assign d1_w[961] = 4'h0;
    assign d1_w[962] = 4'h3;
    assign d1_w[963] = 4'hE;
    assign d1_w[964] = 4'hD;
    assign d1_w[965] = 4'h1;
    assign d1_w[966] = 4'hE;
    assign d1_w[967] = 4'hF;
    assign d1_w[968] = 4'h0;
    assign d1_w[969] = 4'h1;
    assign d1_w[970] = 4'hF;
    assign d1_w[971] = 4'hF;
    assign d1_w[972] = 4'h1;
    assign d1_w[973] = 4'h3;
    assign d1_w[974] = 4'h2;
    assign d1_w[975] = 4'hF;
    assign d1_w[976] = 4'hF;
    assign d1_w[977] = 4'hF;
    assign d1_w[978] = 4'hE;
    assign d1_w[979] = 4'hE;
    assign d1_w[980] = 4'h0;
    assign d1_w[981] = 4'hE;
    assign d1_w[982] = 4'h2;
    assign d1_w[983] = 4'hF;
    assign d1_w[984] = 4'hD;
    assign d1_w[985] = 4'h1;
    assign d1_w[986] = 4'h2;
    assign d1_w[987] = 4'h2;
    assign d1_w[988] = 4'h0;
    assign d1_w[989] = 4'h0;
    assign d1_w[990] = 4'h0;
    assign d1_w[991] = 4'h0;
    assign d1_w[992] = 4'h0;
    assign d1_w[993] = 4'h0;
    assign d1_w[994] = 4'h3;
    assign d1_w[995] = 4'h3;
    assign d1_w[996] = 4'hD;
    assign d1_w[997] = 4'h0;
    assign d1_w[998] = 4'h3;
    assign d1_w[999] = 4'h1;
    assign d1_w[1000] = 4'h1;
    assign d1_w[1001] = 4'h2;
    assign d1_w[1002] = 4'h1;
    assign d1_w[1003] = 4'h1;
    assign d1_w[1004] = 4'hD;
    assign d1_w[1005] = 4'hF;
    assign d1_w[1006] = 4'h0;
    assign d1_w[1007] = 4'h0;
    assign d1_w[1008] = 4'h1;
    assign d1_w[1009] = 4'hE;
    assign d1_w[1010] = 4'h2;
    assign d1_w[1011] = 4'h1;
    assign d1_w[1012] = 4'h3;
    assign d1_w[1013] = 4'h1;
    assign d1_w[1014] = 4'hD;
    assign d1_w[1015] = 4'h0;
    assign d1_w[1016] = 4'h1;
    assign d1_w[1017] = 4'h4;
    assign d1_w[1018] = 4'hF;
    assign d1_w[1019] = 4'h1;
    assign d1_w[1020] = 4'h3;
    assign d1_w[1021] = 4'hF;
    assign d1_w[1022] = 4'hE;
    assign d1_w[1023] = 4'hD;

    // --- layer1_b ---
    assign d1_b[0] = 4'h5;
    assign d1_b[1] = 4'hA;
    assign d1_b[2] = 4'h6;
    assign d1_b[3] = 4'h2;
    assign d1_b[4] = 4'hE;
    assign d1_b[5] = 4'h1;
    assign d1_b[6] = 4'hA;
    assign d1_b[7] = 4'h1;
    assign d1_b[8] = 4'hE;
    assign d1_b[9] = 4'hD;
    assign d1_b[10] = 4'h3;
    assign d1_b[11] = 4'h0;
    assign d1_b[12] = 4'h0;
    assign d1_b[13] = 4'h0;
    assign d1_b[14] = 4'hA;
    assign d1_b[15] = 4'h1;
    assign d1_b[16] = 4'hC;
    assign d1_b[17] = 4'h5;
    assign d1_b[18] = 4'h6;
    assign d1_b[19] = 4'h0;
    assign d1_b[20] = 4'h0;
    assign d1_b[21] = 4'h2;
    assign d1_b[22] = 4'h0;
    assign d1_b[23] = 4'h0;
    assign d1_b[24] = 4'h0;
    assign d1_b[25] = 4'h6;
    assign d1_b[26] = 4'hA;
    assign d1_b[27] = 4'h7;
    assign d1_b[28] = 4'h0;
    assign d1_b[29] = 4'hB;
    assign d1_b[30] = 4'h0;
    assign d1_b[31] = 4'h0;

    // --- layer2_w ---
    assign d2_w[0] = 4'h2;
    assign d2_w[1] = 4'hE;
    assign d2_w[2] = 4'h0;
    assign d2_w[3] = 4'h1;
    assign d2_w[4] = 4'hF;
    assign d2_w[5] = 4'h1;
    assign d2_w[6] = 4'h2;
    assign d2_w[7] = 4'hF;
    assign d2_w[8] = 4'hF;
    assign d2_w[9] = 4'h2;
    assign d2_w[10] = 4'hE;
    assign d2_w[11] = 4'h1;
    assign d2_w[12] = 4'h0;
    assign d2_w[13] = 4'h1;
    assign d2_w[14] = 4'hF;
    assign d2_w[15] = 4'h1;
    assign d2_w[16] = 4'h1;
    assign d2_w[17] = 4'hF;
    assign d2_w[18] = 4'h1;
    assign d2_w[19] = 4'h3;
    assign d2_w[20] = 4'h1;
    assign d2_w[21] = 4'hF;
    assign d2_w[22] = 4'h1;
    assign d2_w[23] = 4'hE;
    assign d2_w[24] = 4'hF;
    assign d2_w[25] = 4'hD;
    assign d2_w[26] = 4'h0;
    assign d2_w[27] = 4'h1;
    assign d2_w[28] = 4'hF;
    assign d2_w[29] = 4'h1;
    assign d2_w[30] = 4'h0;
    assign d2_w[31] = 4'h1;
    assign d2_w[32] = 4'h2;
    assign d2_w[33] = 4'hF;
    assign d2_w[34] = 4'hE;
    assign d2_w[35] = 4'hF;
    assign d2_w[36] = 4'h2;
    assign d2_w[37] = 4'h2;
    assign d2_w[38] = 4'h0;
    assign d2_w[39] = 4'hF;
    assign d2_w[40] = 4'h1;
    assign d2_w[41] = 4'h3;
    assign d2_w[42] = 4'hE;
    assign d2_w[43] = 4'h1;
    assign d2_w[44] = 4'h0;
    assign d2_w[45] = 4'h0;
    assign d2_w[46] = 4'h0;
    assign d2_w[47] = 4'hE;
    assign d2_w[48] = 4'hE;
    assign d2_w[49] = 4'hF;
    assign d2_w[50] = 4'h1;
    assign d2_w[51] = 4'hE;
    assign d2_w[52] = 4'hF;
    assign d2_w[53] = 4'hE;
    assign d2_w[54] = 4'hE;
    assign d2_w[55] = 4'h2;
    assign d2_w[56] = 4'h2;
    assign d2_w[57] = 4'h1;
    assign d2_w[58] = 4'h1;
    assign d2_w[59] = 4'h2;
    assign d2_w[60] = 4'hF;
    assign d2_w[61] = 4'h0;
    assign d2_w[62] = 4'h0;
    assign d2_w[63] = 4'h2;
    assign d2_w[64] = 4'hF;
    assign d2_w[65] = 4'h2;
    assign d2_w[66] = 4'h1;
    assign d2_w[67] = 4'h1;
    assign d2_w[68] = 4'hF;
    assign d2_w[69] = 4'h2;
    assign d2_w[70] = 4'h1;
    assign d2_w[71] = 4'hF;
    assign d2_w[72] = 4'h2;
    assign d2_w[73] = 4'h0;
    assign d2_w[74] = 4'hE;
    assign d2_w[75] = 4'h2;
    assign d2_w[76] = 4'hF;
    assign d2_w[77] = 4'h2;
    assign d2_w[78] = 4'h3;
    assign d2_w[79] = 4'h2;
    assign d2_w[80] = 4'hF;
    assign d2_w[81] = 4'h0;
    assign d2_w[82] = 4'h1;
    assign d2_w[83] = 4'h0;
    assign d2_w[84] = 4'h1;
    assign d2_w[85] = 4'h0;
    assign d2_w[86] = 4'h0;
    assign d2_w[87] = 4'hF;
    assign d2_w[88] = 4'h1;
    assign d2_w[89] = 4'hE;
    assign d2_w[90] = 4'hF;
    assign d2_w[91] = 4'h1;
    assign d2_w[92] = 4'hE;
    assign d2_w[93] = 4'h1;
    assign d2_w[94] = 4'hF;
    assign d2_w[95] = 4'h1;
    assign d2_w[96] = 4'h3;
    assign d2_w[97] = 4'h2;
    assign d2_w[98] = 4'h1;
    assign d2_w[99] = 4'h3;
    assign d2_w[100] = 4'h0;
    assign d2_w[101] = 4'hF;
    assign d2_w[102] = 4'h2;
    assign d2_w[103] = 4'h3;
    assign d2_w[104] = 4'hF;
    assign d2_w[105] = 4'h0;
    assign d2_w[106] = 4'hF;
    assign d2_w[107] = 4'h2;
    assign d2_w[108] = 4'hF;
    assign d2_w[109] = 4'h3;
    assign d2_w[110] = 4'h2;
    assign d2_w[111] = 4'h1;
    assign d2_w[112] = 4'hD;
    assign d2_w[113] = 4'hF;
    assign d2_w[114] = 4'hF;
    assign d2_w[115] = 4'hE;
    assign d2_w[116] = 4'h2;
    assign d2_w[117] = 4'h3;
    assign d2_w[118] = 4'h3;
    assign d2_w[119] = 4'h1;
    assign d2_w[120] = 4'h1;
    assign d2_w[121] = 4'h0;
    assign d2_w[122] = 4'h0;
    assign d2_w[123] = 4'hF;
    assign d2_w[124] = 4'hE;
    assign d2_w[125] = 4'hE;
    assign d2_w[126] = 4'h2;
    assign d2_w[127] = 4'hE;
    assign d2_w[128] = 4'h0;
    assign d2_w[129] = 4'h1;
    assign d2_w[130] = 4'hE;
    assign d2_w[131] = 4'h1;
    assign d2_w[132] = 4'h1;
    assign d2_w[133] = 4'h0;
    assign d2_w[134] = 4'h0;
    assign d2_w[135] = 4'hF;
    assign d2_w[136] = 4'h2;
    assign d2_w[137] = 4'hE;
    assign d2_w[138] = 4'hF;
    assign d2_w[139] = 4'h2;
    assign d2_w[140] = 4'hF;
    assign d2_w[141] = 4'hE;
    assign d2_w[142] = 4'h2;
    assign d2_w[143] = 4'hE;
    assign d2_w[144] = 4'hE;
    assign d2_w[145] = 4'h2;
    assign d2_w[146] = 4'h1;
    assign d2_w[147] = 4'h0;
    assign d2_w[148] = 4'hF;
    assign d2_w[149] = 4'h2;
    assign d2_w[150] = 4'h0;
    assign d2_w[151] = 4'h1;
    assign d2_w[152] = 4'hF;
    assign d2_w[153] = 4'hD;
    assign d2_w[154] = 4'h1;
    assign d2_w[155] = 4'hE;
    assign d2_w[156] = 4'hF;
    assign d2_w[157] = 4'hF;
    assign d2_w[158] = 4'hE;
    assign d2_w[159] = 4'hF;
    assign d2_w[160] = 4'h1;
    assign d2_w[161] = 4'h2;
    assign d2_w[162] = 4'h0;
    assign d2_w[163] = 4'h2;
    assign d2_w[164] = 4'h1;
    assign d2_w[165] = 4'h3;
    assign d2_w[166] = 4'hE;
    assign d2_w[167] = 4'h2;
    assign d2_w[168] = 4'h0;
    assign d2_w[169] = 4'h0;
    assign d2_w[170] = 4'h0;
    assign d2_w[171] = 4'h0;
    assign d2_w[172] = 4'h2;
    assign d2_w[173] = 4'hF;
    assign d2_w[174] = 4'hF;
    assign d2_w[175] = 4'hF;
    assign d2_w[176] = 4'hE;
    assign d2_w[177] = 4'h2;
    assign d2_w[178] = 4'h0;
    assign d2_w[179] = 4'h0;
    assign d2_w[180] = 4'h0;
    assign d2_w[181] = 4'hE;
    assign d2_w[182] = 4'hE;
    assign d2_w[183] = 4'hD;
    assign d2_w[184] = 4'h1;
    assign d2_w[185] = 4'hF;
    assign d2_w[186] = 4'hF;
    assign d2_w[187] = 4'h2;
    assign d2_w[188] = 4'h0;
    assign d2_w[189] = 4'h2;
    assign d2_w[190] = 4'h1;
    assign d2_w[191] = 4'hF;
    assign d2_w[192] = 4'h1;
    assign d2_w[193] = 4'hE;
    assign d2_w[194] = 4'hD;
    assign d2_w[195] = 4'h1;
    assign d2_w[196] = 4'h2;
    assign d2_w[197] = 4'h0;
    assign d2_w[198] = 4'hE;
    assign d2_w[199] = 4'h0;
    assign d2_w[200] = 4'hD;
    assign d2_w[201] = 4'h2;
    assign d2_w[202] = 4'hF;
    assign d2_w[203] = 4'hF;
    assign d2_w[204] = 4'h1;
    assign d2_w[205] = 4'hC;
    assign d2_w[206] = 4'hF;
    assign d2_w[207] = 4'hE;
    assign d2_w[208] = 4'h0;
    assign d2_w[209] = 4'hF;
    assign d2_w[210] = 4'h3;
    assign d2_w[211] = 4'h0;
    assign d2_w[212] = 4'hF;
    assign d2_w[213] = 4'h0;
    assign d2_w[214] = 4'hD;
    assign d2_w[215] = 4'h1;
    assign d2_w[216] = 4'h2;
    assign d2_w[217] = 4'h2;
    assign d2_w[218] = 4'hF;
    assign d2_w[219] = 4'h0;
    assign d2_w[220] = 4'h0;
    assign d2_w[221] = 4'h0;
    assign d2_w[222] = 4'h0;
    assign d2_w[223] = 4'hF;
    assign d2_w[224] = 4'h0;
    assign d2_w[225] = 4'h1;
    assign d2_w[226] = 4'h0;
    assign d2_w[227] = 4'hF;
    assign d2_w[228] = 4'h0;
    assign d2_w[229] = 4'h2;
    assign d2_w[230] = 4'hE;
    assign d2_w[231] = 4'h1;
    assign d2_w[232] = 4'hF;
    assign d2_w[233] = 4'hE;
    assign d2_w[234] = 4'h1;
    assign d2_w[235] = 4'h0;
    assign d2_w[236] = 4'h0;
    assign d2_w[237] = 4'h0;
    assign d2_w[238] = 4'h2;
    assign d2_w[239] = 4'h1;
    assign d2_w[240] = 4'hF;
    assign d2_w[241] = 4'h2;
    assign d2_w[242] = 4'hE;
    assign d2_w[243] = 4'hF;
    assign d2_w[244] = 4'hF;
    assign d2_w[245] = 4'hE;
    assign d2_w[246] = 4'h2;
    assign d2_w[247] = 4'h0;
    assign d2_w[248] = 4'h0;
    assign d2_w[249] = 4'h1;
    assign d2_w[250] = 4'h0;
    assign d2_w[251] = 4'h1;
    assign d2_w[252] = 4'hF;
    assign d2_w[253] = 4'h1;
    assign d2_w[254] = 4'h1;
    assign d2_w[255] = 4'hE;
    assign d2_w[256] = 4'h2;
    assign d2_w[257] = 4'hF;
    assign d2_w[258] = 4'h2;
    assign d2_w[259] = 4'hE;
    assign d2_w[260] = 4'hF;
    assign d2_w[261] = 4'h2;
    assign d2_w[262] = 4'hE;
    assign d2_w[263] = 4'h2;
    assign d2_w[264] = 4'h2;
    assign d2_w[265] = 4'hF;
    assign d2_w[266] = 4'hE;
    assign d2_w[267] = 4'h2;
    assign d2_w[268] = 4'h2;
    assign d2_w[269] = 4'h1;
    assign d2_w[270] = 4'h1;
    assign d2_w[271] = 4'hE;
    assign d2_w[272] = 4'hE;
    assign d2_w[273] = 4'h0;
    assign d2_w[274] = 4'h2;
    assign d2_w[275] = 4'h2;
    assign d2_w[276] = 4'hE;
    assign d2_w[277] = 4'h1;
    assign d2_w[278] = 4'h0;
    assign d2_w[279] = 4'h1;
    assign d2_w[280] = 4'h0;
    assign d2_w[281] = 4'hF;
    assign d2_w[282] = 4'h1;
    assign d2_w[283] = 4'hE;
    assign d2_w[284] = 4'hF;
    assign d2_w[285] = 4'hE;
    assign d2_w[286] = 4'h0;
    assign d2_w[287] = 4'hF;
    assign d2_w[288] = 4'hE;
    assign d2_w[289] = 4'h0;
    assign d2_w[290] = 4'h1;
    assign d2_w[291] = 4'hF;
    assign d2_w[292] = 4'h1;
    assign d2_w[293] = 4'h0;
    assign d2_w[294] = 4'h1;
    assign d2_w[295] = 4'h0;
    assign d2_w[296] = 4'h2;
    assign d2_w[297] = 4'hF;
    assign d2_w[298] = 4'h2;
    assign d2_w[299] = 4'hF;
    assign d2_w[300] = 4'h1;
    assign d2_w[301] = 4'h1;
    assign d2_w[302] = 4'h0;
    assign d2_w[303] = 4'hF;
    assign d2_w[304] = 4'hE;
    assign d2_w[305] = 4'hE;
    assign d2_w[306] = 4'h0;
    assign d2_w[307] = 4'h0;
    assign d2_w[308] = 4'hE;
    assign d2_w[309] = 4'hF;
    assign d2_w[310] = 4'h0;
    assign d2_w[311] = 4'h0;
    assign d2_w[312] = 4'h2;
    assign d2_w[313] = 4'h1;
    assign d2_w[314] = 4'h2;
    assign d2_w[315] = 4'hE;
    assign d2_w[316] = 4'h0;
    assign d2_w[317] = 4'h0;
    assign d2_w[318] = 4'h1;
    assign d2_w[319] = 4'hE;
    assign d2_w[320] = 4'h2;
    assign d2_w[321] = 4'h0;
    assign d2_w[322] = 4'hF;
    assign d2_w[323] = 4'hF;
    assign d2_w[324] = 4'h2;
    assign d2_w[325] = 4'h0;
    assign d2_w[326] = 4'h2;
    assign d2_w[327] = 4'h0;
    assign d2_w[328] = 4'hE;
    assign d2_w[329] = 4'h0;
    assign d2_w[330] = 4'h0;
    assign d2_w[331] = 4'hE;
    assign d2_w[332] = 4'hF;
    assign d2_w[333] = 4'hF;
    assign d2_w[334] = 4'h2;
    assign d2_w[335] = 4'hF;
    assign d2_w[336] = 4'h1;
    assign d2_w[337] = 4'h1;
    assign d2_w[338] = 4'h1;
    assign d2_w[339] = 4'h0;
    assign d2_w[340] = 4'hE;
    assign d2_w[341] = 4'h0;
    assign d2_w[342] = 4'h2;
    assign d2_w[343] = 4'hE;
    assign d2_w[344] = 4'hF;
    assign d2_w[345] = 4'hE;
    assign d2_w[346] = 4'h0;
    assign d2_w[347] = 4'h1;
    assign d2_w[348] = 4'h2;
    assign d2_w[349] = 4'h2;
    assign d2_w[350] = 4'h1;
    assign d2_w[351] = 4'h0;
    assign d2_w[352] = 4'hF;
    assign d2_w[353] = 4'hD;
    assign d2_w[354] = 4'h0;
    assign d2_w[355] = 4'h0;
    assign d2_w[356] = 4'h1;
    assign d2_w[357] = 4'h1;
    assign d2_w[358] = 4'hF;
    assign d2_w[359] = 4'hE;
    assign d2_w[360] = 4'h1;
    assign d2_w[361] = 4'h0;
    assign d2_w[362] = 4'h0;
    assign d2_w[363] = 4'hE;
    assign d2_w[364] = 4'hF;
    assign d2_w[365] = 4'h0;
    assign d2_w[366] = 4'h1;
    assign d2_w[367] = 4'hF;
    assign d2_w[368] = 4'h1;
    assign d2_w[369] = 4'hE;
    assign d2_w[370] = 4'h0;
    assign d2_w[371] = 4'h1;
    assign d2_w[372] = 4'h0;
    assign d2_w[373] = 4'hF;
    assign d2_w[374] = 4'hF;
    assign d2_w[375] = 4'hF;
    assign d2_w[376] = 4'h0;
    assign d2_w[377] = 4'hF;
    assign d2_w[378] = 4'h2;
    assign d2_w[379] = 4'hE;
    assign d2_w[380] = 4'hF;
    assign d2_w[381] = 4'h1;
    assign d2_w[382] = 4'hE;
    assign d2_w[383] = 4'hE;
    assign d2_w[384] = 4'h1;
    assign d2_w[385] = 4'h2;
    assign d2_w[386] = 4'hE;
    assign d2_w[387] = 4'h0;
    assign d2_w[388] = 4'h1;
    assign d2_w[389] = 4'hF;
    assign d2_w[390] = 4'h0;
    assign d2_w[391] = 4'h0;
    assign d2_w[392] = 4'h2;
    assign d2_w[393] = 4'hE;
    assign d2_w[394] = 4'h2;
    assign d2_w[395] = 4'hE;
    assign d2_w[396] = 4'h2;
    assign d2_w[397] = 4'h1;
    assign d2_w[398] = 4'hE;
    assign d2_w[399] = 4'hF;
    assign d2_w[400] = 4'h0;
    assign d2_w[401] = 4'hF;
    assign d2_w[402] = 4'hF;
    assign d2_w[403] = 4'h0;
    assign d2_w[404] = 4'h0;
    assign d2_w[405] = 4'h0;
    assign d2_w[406] = 4'h1;
    assign d2_w[407] = 4'hF;
    assign d2_w[408] = 4'hE;
    assign d2_w[409] = 4'h0;
    assign d2_w[410] = 4'h0;
    assign d2_w[411] = 4'hF;
    assign d2_w[412] = 4'hF;
    assign d2_w[413] = 4'hF;
    assign d2_w[414] = 4'h1;
    assign d2_w[415] = 4'hE;
    assign d2_w[416] = 4'hE;
    assign d2_w[417] = 4'h2;
    assign d2_w[418] = 4'h0;
    assign d2_w[419] = 4'h1;
    assign d2_w[420] = 4'h2;
    assign d2_w[421] = 4'h0;
    assign d2_w[422] = 4'h0;
    assign d2_w[423] = 4'hF;
    assign d2_w[424] = 4'h0;
    assign d2_w[425] = 4'hE;
    assign d2_w[426] = 4'hF;
    assign d2_w[427] = 4'hE;
    assign d2_w[428] = 4'hF;
    assign d2_w[429] = 4'hF;
    assign d2_w[430] = 4'hF;
    assign d2_w[431] = 4'h2;
    assign d2_w[432] = 4'hF;
    assign d2_w[433] = 4'hE;
    assign d2_w[434] = 4'hF;
    assign d2_w[435] = 4'h2;
    assign d2_w[436] = 4'h0;
    assign d2_w[437] = 4'h1;
    assign d2_w[438] = 4'h2;
    assign d2_w[439] = 4'h0;
    assign d2_w[440] = 4'h0;
    assign d2_w[441] = 4'hE;
    assign d2_w[442] = 4'h0;
    assign d2_w[443] = 4'h0;
    assign d2_w[444] = 4'h1;
    assign d2_w[445] = 4'h1;
    assign d2_w[446] = 4'hE;
    assign d2_w[447] = 4'h2;
    assign d2_w[448] = 4'hE;
    assign d2_w[449] = 4'h1;
    assign d2_w[450] = 4'hE;
    assign d2_w[451] = 4'h0;
    assign d2_w[452] = 4'hF;
    assign d2_w[453] = 4'hE;
    assign d2_w[454] = 4'h1;
    assign d2_w[455] = 4'hE;
    assign d2_w[456] = 4'h1;
    assign d2_w[457] = 4'hF;
    assign d2_w[458] = 4'hE;
    assign d2_w[459] = 4'hF;
    assign d2_w[460] = 4'h2;
    assign d2_w[461] = 4'hE;
    assign d2_w[462] = 4'h3;
    assign d2_w[463] = 4'hE;
    assign d2_w[464] = 4'hF;
    assign d2_w[465] = 4'h0;
    assign d2_w[466] = 4'hE;
    assign d2_w[467] = 4'h1;
    assign d2_w[468] = 4'h2;
    assign d2_w[469] = 4'h0;
    assign d2_w[470] = 4'hD;
    assign d2_w[471] = 4'h0;
    assign d2_w[472] = 4'h0;
    assign d2_w[473] = 4'h0;
    assign d2_w[474] = 4'hE;
    assign d2_w[475] = 4'h2;
    assign d2_w[476] = 4'h0;
    assign d2_w[477] = 4'h2;
    assign d2_w[478] = 4'hF;
    assign d2_w[479] = 4'hF;
    assign d2_w[480] = 4'hF;
    assign d2_w[481] = 4'h1;
    assign d2_w[482] = 4'h0;
    assign d2_w[483] = 4'h3;
    assign d2_w[484] = 4'h0;
    assign d2_w[485] = 4'h0;
    assign d2_w[486] = 4'h3;
    assign d2_w[487] = 4'hE;
    assign d2_w[488] = 4'h0;
    assign d2_w[489] = 4'h2;
    assign d2_w[490] = 4'hF;
    assign d2_w[491] = 4'hF;
    assign d2_w[492] = 4'h3;
    assign d2_w[493] = 4'h2;
    assign d2_w[494] = 4'h3;
    assign d2_w[495] = 4'h1;
    assign d2_w[496] = 4'h0;
    assign d2_w[497] = 4'h0;
    assign d2_w[498] = 4'hA;
    assign d2_w[499] = 4'hF;
    assign d2_w[500] = 4'h1;
    assign d2_w[501] = 4'h1;
    assign d2_w[502] = 4'h3;
    assign d2_w[503] = 4'hF;
    assign d2_w[504] = 4'h2;
    assign d2_w[505] = 4'h1;
    assign d2_w[506] = 4'h2;
    assign d2_w[507] = 4'h1;
    assign d2_w[508] = 4'h1;
    assign d2_w[509] = 4'h3;
    assign d2_w[510] = 4'h2;
    assign d2_w[511] = 4'hE;
    assign d2_w[512] = 4'hE;
    assign d2_w[513] = 4'h1;
    assign d2_w[514] = 4'hF;
    assign d2_w[515] = 4'h1;
    assign d2_w[516] = 4'h0;
    assign d2_w[517] = 4'hE;
    assign d2_w[518] = 4'h0;
    assign d2_w[519] = 4'h2;
    assign d2_w[520] = 4'h2;
    assign d2_w[521] = 4'h2;
    assign d2_w[522] = 4'h1;
    assign d2_w[523] = 4'h0;
    assign d2_w[524] = 4'h2;
    assign d2_w[525] = 4'hE;
    assign d2_w[526] = 4'h2;
    assign d2_w[527] = 4'h0;
    assign d2_w[528] = 4'hF;
    assign d2_w[529] = 4'h2;
    assign d2_w[530] = 4'h0;
    assign d2_w[531] = 4'h2;
    assign d2_w[532] = 4'h2;
    assign d2_w[533] = 4'hF;
    assign d2_w[534] = 4'h0;
    assign d2_w[535] = 4'hF;
    assign d2_w[536] = 4'h2;
    assign d2_w[537] = 4'hE;
    assign d2_w[538] = 4'h1;
    assign d2_w[539] = 4'hE;
    assign d2_w[540] = 4'hF;
    assign d2_w[541] = 4'hE;
    assign d2_w[542] = 4'h1;
    assign d2_w[543] = 4'hF;
    assign d2_w[544] = 4'h1;
    assign d2_w[545] = 4'h0;
    assign d2_w[546] = 4'h3;
    assign d2_w[547] = 4'hF;
    assign d2_w[548] = 4'h0;
    assign d2_w[549] = 4'hF;
    assign d2_w[550] = 4'h1;
    assign d2_w[551] = 4'h1;
    assign d2_w[552] = 4'h0;
    assign d2_w[553] = 4'h2;
    assign d2_w[554] = 4'hF;
    assign d2_w[555] = 4'h3;
    assign d2_w[556] = 4'hF;
    assign d2_w[557] = 4'h4;
    assign d2_w[558] = 4'h3;
    assign d2_w[559] = 4'h2;
    assign d2_w[560] = 4'h2;
    assign d2_w[561] = 4'h1;
    assign d2_w[562] = 4'h0;
    assign d2_w[563] = 4'hF;
    assign d2_w[564] = 4'h3;
    assign d2_w[565] = 4'h1;
    assign d2_w[566] = 4'h4;
    assign d2_w[567] = 4'h1;
    assign d2_w[568] = 4'h1;
    assign d2_w[569] = 4'h1;
    assign d2_w[570] = 4'hE;
    assign d2_w[571] = 4'hE;
    assign d2_w[572] = 4'hF;
    assign d2_w[573] = 4'h3;
    assign d2_w[574] = 4'h3;
    assign d2_w[575] = 4'hE;
    assign d2_w[576] = 4'h4;
    assign d2_w[577] = 4'h4;
    assign d2_w[578] = 4'h1;
    assign d2_w[579] = 4'h4;
    assign d2_w[580] = 4'h1;
    assign d2_w[581] = 4'hF;
    assign d2_w[582] = 4'h4;
    assign d2_w[583] = 4'h4;
    assign d2_w[584] = 4'h0;
    assign d2_w[585] = 4'h1;
    assign d2_w[586] = 4'hF;
    assign d2_w[587] = 4'h2;
    assign d2_w[588] = 4'hE;
    assign d2_w[589] = 4'h6;
    assign d2_w[590] = 4'h4;
    assign d2_w[591] = 4'h4;
    assign d2_w[592] = 4'h0;
    assign d2_w[593] = 4'hF;
    assign d2_w[594] = 4'h3;
    assign d2_w[595] = 4'hF;
    assign d2_w[596] = 4'h4;
    assign d2_w[597] = 4'h1;
    assign d2_w[598] = 4'h4;
    assign d2_w[599] = 4'h1;
    assign d2_w[600] = 4'hD;
    assign d2_w[601] = 4'h0;
    assign d2_w[602] = 4'hE;
    assign d2_w[603] = 4'hF;
    assign d2_w[604] = 4'hF;
    assign d2_w[605] = 4'h5;
    assign d2_w[606] = 4'h6;
    assign d2_w[607] = 4'hE;
    assign d2_w[608] = 4'h1;
    assign d2_w[609] = 4'h0;
    assign d2_w[610] = 4'h2;
    assign d2_w[611] = 4'hF;
    assign d2_w[612] = 4'h2;
    assign d2_w[613] = 4'h1;
    assign d2_w[614] = 4'hE;
    assign d2_w[615] = 4'hE;
    assign d2_w[616] = 4'hF;
    assign d2_w[617] = 4'h0;
    assign d2_w[618] = 4'h2;
    assign d2_w[619] = 4'h1;
    assign d2_w[620] = 4'h0;
    assign d2_w[621] = 4'hF;
    assign d2_w[622] = 4'hE;
    assign d2_w[623] = 4'h1;
    assign d2_w[624] = 4'h0;
    assign d2_w[625] = 4'h2;
    assign d2_w[626] = 4'hF;
    assign d2_w[627] = 4'h0;
    assign d2_w[628] = 4'hE;
    assign d2_w[629] = 4'h1;
    assign d2_w[630] = 4'hE;
    assign d2_w[631] = 4'hF;
    assign d2_w[632] = 4'hF;
    assign d2_w[633] = 4'h0;
    assign d2_w[634] = 4'hE;
    assign d2_w[635] = 4'h0;
    assign d2_w[636] = 4'h1;
    assign d2_w[637] = 4'h1;
    assign d2_w[638] = 4'hF;
    assign d2_w[639] = 4'hE;
    assign d2_w[640] = 4'h0;
    assign d2_w[641] = 4'h2;
    assign d2_w[642] = 4'h2;
    assign d2_w[643] = 4'h3;
    assign d2_w[644] = 4'h0;
    assign d2_w[645] = 4'hF;
    assign d2_w[646] = 4'h2;
    assign d2_w[647] = 4'h2;
    assign d2_w[648] = 4'h1;
    assign d2_w[649] = 4'hF;
    assign d2_w[650] = 4'h0;
    assign d2_w[651] = 4'h0;
    assign d2_w[652] = 4'h1;
    assign d2_w[653] = 4'h2;
    assign d2_w[654] = 4'h3;
    assign d2_w[655] = 4'h1;
    assign d2_w[656] = 4'hF;
    assign d2_w[657] = 4'h0;
    assign d2_w[658] = 4'h9;
    assign d2_w[659] = 4'h0;
    assign d2_w[660] = 4'h3;
    assign d2_w[661] = 4'h2;
    assign d2_w[662] = 4'h1;
    assign d2_w[663] = 4'h0;
    assign d2_w[664] = 4'hE;
    assign d2_w[665] = 4'h2;
    assign d2_w[666] = 4'hF;
    assign d2_w[667] = 4'hF;
    assign d2_w[668] = 4'hF;
    assign d2_w[669] = 4'h3;
    assign d2_w[670] = 4'hF;
    assign d2_w[671] = 4'h0;
    assign d2_w[672] = 4'hE;
    assign d2_w[673] = 4'h1;
    assign d2_w[674] = 4'h0;
    assign d2_w[675] = 4'hE;
    assign d2_w[676] = 4'hF;
    assign d2_w[677] = 4'hF;
    assign d2_w[678] = 4'h1;
    assign d2_w[679] = 4'h2;
    assign d2_w[680] = 4'hE;
    assign d2_w[681] = 4'hE;
    assign d2_w[682] = 4'h2;
    assign d2_w[683] = 4'h1;
    assign d2_w[684] = 4'hF;
    assign d2_w[685] = 4'h0;
    assign d2_w[686] = 4'hF;
    assign d2_w[687] = 4'h1;
    assign d2_w[688] = 4'h0;
    assign d2_w[689] = 4'h3;
    assign d2_w[690] = 4'h2;
    assign d2_w[691] = 4'h0;
    assign d2_w[692] = 4'h1;
    assign d2_w[693] = 4'hF;
    assign d2_w[694] = 4'h0;
    assign d2_w[695] = 4'h0;
    assign d2_w[696] = 4'hF;
    assign d2_w[697] = 4'h0;
    assign d2_w[698] = 4'h0;
    assign d2_w[699] = 4'h2;
    assign d2_w[700] = 4'h2;
    assign d2_w[701] = 4'h0;
    assign d2_w[702] = 4'h2;
    assign d2_w[703] = 4'hE;
    assign d2_w[704] = 4'h0;
    assign d2_w[705] = 4'h2;
    assign d2_w[706] = 4'hF;
    assign d2_w[707] = 4'hF;
    assign d2_w[708] = 4'h0;
    assign d2_w[709] = 4'hE;
    assign d2_w[710] = 4'h0;
    assign d2_w[711] = 4'hE;
    assign d2_w[712] = 4'hF;
    assign d2_w[713] = 4'h0;
    assign d2_w[714] = 4'h0;
    assign d2_w[715] = 4'h0;
    assign d2_w[716] = 4'h0;
    assign d2_w[717] = 4'h2;
    assign d2_w[718] = 4'hE;
    assign d2_w[719] = 4'hE;
    assign d2_w[720] = 4'hF;
    assign d2_w[721] = 4'hE;
    assign d2_w[722] = 4'hF;
    assign d2_w[723] = 4'h0;
    assign d2_w[724] = 4'h1;
    assign d2_w[725] = 4'h2;
    assign d2_w[726] = 4'h0;
    assign d2_w[727] = 4'hF;
    assign d2_w[728] = 4'hF;
    assign d2_w[729] = 4'h0;
    assign d2_w[730] = 4'h1;
    assign d2_w[731] = 4'h0;
    assign d2_w[732] = 4'h2;
    assign d2_w[733] = 4'h1;
    assign d2_w[734] = 4'hF;
    assign d2_w[735] = 4'h1;
    assign d2_w[736] = 4'h0;
    assign d2_w[737] = 4'hF;
    assign d2_w[738] = 4'h1;
    assign d2_w[739] = 4'hF;
    assign d2_w[740] = 4'hF;
    assign d2_w[741] = 4'h1;
    assign d2_w[742] = 4'h1;
    assign d2_w[743] = 4'hE;
    assign d2_w[744] = 4'hE;
    assign d2_w[745] = 4'hF;
    assign d2_w[746] = 4'hE;
    assign d2_w[747] = 4'h1;
    assign d2_w[748] = 4'hE;
    assign d2_w[749] = 4'h1;
    assign d2_w[750] = 4'h2;
    assign d2_w[751] = 4'h0;
    assign d2_w[752] = 4'hF;
    assign d2_w[753] = 4'h0;
    assign d2_w[754] = 4'h1;
    assign d2_w[755] = 4'hE;
    assign d2_w[756] = 4'h0;
    assign d2_w[757] = 4'hF;
    assign d2_w[758] = 4'h2;
    assign d2_w[759] = 4'h2;
    assign d2_w[760] = 4'h2;
    assign d2_w[761] = 4'h1;
    assign d2_w[762] = 4'h1;
    assign d2_w[763] = 4'hE;
    assign d2_w[764] = 4'hF;
    assign d2_w[765] = 4'h1;
    assign d2_w[766] = 4'hF;
    assign d2_w[767] = 4'h0;
    assign d2_w[768] = 4'h2;
    assign d2_w[769] = 4'h2;
    assign d2_w[770] = 4'h2;
    assign d2_w[771] = 4'h2;
    assign d2_w[772] = 4'h1;
    assign d2_w[773] = 4'hF;
    assign d2_w[774] = 4'hE;
    assign d2_w[775] = 4'h1;
    assign d2_w[776] = 4'h2;
    assign d2_w[777] = 4'h0;
    assign d2_w[778] = 4'h2;
    assign d2_w[779] = 4'h2;
    assign d2_w[780] = 4'hE;
    assign d2_w[781] = 4'hE;
    assign d2_w[782] = 4'hE;
    assign d2_w[783] = 4'h1;
    assign d2_w[784] = 4'hF;
    assign d2_w[785] = 4'hE;
    assign d2_w[786] = 4'h1;
    assign d2_w[787] = 4'h0;
    assign d2_w[788] = 4'hE;
    assign d2_w[789] = 4'hE;
    assign d2_w[790] = 4'h2;
    assign d2_w[791] = 4'hF;
    assign d2_w[792] = 4'hE;
    assign d2_w[793] = 4'h1;
    assign d2_w[794] = 4'hF;
    assign d2_w[795] = 4'h0;
    assign d2_w[796] = 4'h1;
    assign d2_w[797] = 4'hF;
    assign d2_w[798] = 4'hE;
    assign d2_w[799] = 4'h0;
    assign d2_w[800] = 4'h1;
    assign d2_w[801] = 4'h0;
    assign d2_w[802] = 4'h2;
    assign d2_w[803] = 4'h2;
    assign d2_w[804] = 4'h2;
    assign d2_w[805] = 4'h1;
    assign d2_w[806] = 4'hF;
    assign d2_w[807] = 4'h3;
    assign d2_w[808] = 4'hD;
    assign d2_w[809] = 4'h2;
    assign d2_w[810] = 4'h0;
    assign d2_w[811] = 4'h2;
    assign d2_w[812] = 4'h0;
    assign d2_w[813] = 4'h1;
    assign d2_w[814] = 4'hE;
    assign d2_w[815] = 4'h1;
    assign d2_w[816] = 4'h0;
    assign d2_w[817] = 4'hE;
    assign d2_w[818] = 4'h2;
    assign d2_w[819] = 4'h2;
    assign d2_w[820] = 4'h2;
    assign d2_w[821] = 4'hF;
    assign d2_w[822] = 4'h1;
    assign d2_w[823] = 4'h1;
    assign d2_w[824] = 4'h2;
    assign d2_w[825] = 4'h1;
    assign d2_w[826] = 4'h1;
    assign d2_w[827] = 4'h1;
    assign d2_w[828] = 4'hF;
    assign d2_w[829] = 4'h3;
    assign d2_w[830] = 4'h1;
    assign d2_w[831] = 4'h1;
    assign d2_w[832] = 4'hD;
    assign d2_w[833] = 4'h1;
    assign d2_w[834] = 4'hE;
    assign d2_w[835] = 4'h0;
    assign d2_w[836] = 4'hF;
    assign d2_w[837] = 4'hF;
    assign d2_w[838] = 4'h2;
    assign d2_w[839] = 4'hF;
    assign d2_w[840] = 4'hE;
    assign d2_w[841] = 4'h2;
    assign d2_w[842] = 4'hE;
    assign d2_w[843] = 4'hE;
    assign d2_w[844] = 4'h0;
    assign d2_w[845] = 4'hE;
    assign d2_w[846] = 4'hE;
    assign d2_w[847] = 4'h0;
    assign d2_w[848] = 4'h2;
    assign d2_w[849] = 4'h0;
    assign d2_w[850] = 4'hF;
    assign d2_w[851] = 4'hF;
    assign d2_w[852] = 4'h2;
    assign d2_w[853] = 4'hC;
    assign d2_w[854] = 4'h0;
    assign d2_w[855] = 4'hF;
    assign d2_w[856] = 4'h0;
    assign d2_w[857] = 4'h0;
    assign d2_w[858] = 4'h0;
    assign d2_w[859] = 4'h1;
    assign d2_w[860] = 4'h1;
    assign d2_w[861] = 4'h1;
    assign d2_w[862] = 4'hD;
    assign d2_w[863] = 4'hF;
    assign d2_w[864] = 4'h1;
    assign d2_w[865] = 4'h4;
    assign d2_w[866] = 4'h4;
    assign d2_w[867] = 4'h1;
    assign d2_w[868] = 4'h4;
    assign d2_w[869] = 4'h0;
    assign d2_w[870] = 4'h1;
    assign d2_w[871] = 4'h4;
    assign d2_w[872] = 4'h3;
    assign d2_w[873] = 4'h0;
    assign d2_w[874] = 4'h1;
    assign d2_w[875] = 4'h4;
    assign d2_w[876] = 4'hD;
    assign d2_w[877] = 4'h6;
    assign d2_w[878] = 4'h3;
    assign d2_w[879] = 4'h5;
    assign d2_w[880] = 4'hE;
    assign d2_w[881] = 4'hF;
    assign d2_w[882] = 4'h2;
    assign d2_w[883] = 4'hE;
    assign d2_w[884] = 4'h4;
    assign d2_w[885] = 4'h0;
    assign d2_w[886] = 4'h6;
    assign d2_w[887] = 4'h0;
    assign d2_w[888] = 4'h2;
    assign d2_w[889] = 4'hF;
    assign d2_w[890] = 4'h0;
    assign d2_w[891] = 4'h1;
    assign d2_w[892] = 4'h0;
    assign d2_w[893] = 4'h5;
    assign d2_w[894] = 4'h1;
    assign d2_w[895] = 4'hF;
    assign d2_w[896] = 4'hE;
    assign d2_w[897] = 4'h1;
    assign d2_w[898] = 4'h3;
    assign d2_w[899] = 4'hF;
    assign d2_w[900] = 4'h1;
    assign d2_w[901] = 4'hF;
    assign d2_w[902] = 4'h0;
    assign d2_w[903] = 4'h2;
    assign d2_w[904] = 4'hE;
    assign d2_w[905] = 4'h1;
    assign d2_w[906] = 4'hE;
    assign d2_w[907] = 4'h0;
    assign d2_w[908] = 4'h1;
    assign d2_w[909] = 4'hE;
    assign d2_w[910] = 4'h2;
    assign d2_w[911] = 4'h0;
    assign d2_w[912] = 4'h1;
    assign d2_w[913] = 4'h1;
    assign d2_w[914] = 4'h0;
    assign d2_w[915] = 4'h2;
    assign d2_w[916] = 4'h0;
    assign d2_w[917] = 4'h0;
    assign d2_w[918] = 4'h0;
    assign d2_w[919] = 4'hE;
    assign d2_w[920] = 4'hF;
    assign d2_w[921] = 4'h1;
    assign d2_w[922] = 4'h1;
    assign d2_w[923] = 4'h0;
    assign d2_w[924] = 4'h0;
    assign d2_w[925] = 4'h0;
    assign d2_w[926] = 4'hF;
    assign d2_w[927] = 4'hE;
    assign d2_w[928] = 4'h2;
    assign d2_w[929] = 4'h2;
    assign d2_w[930] = 4'h2;
    assign d2_w[931] = 4'h2;
    assign d2_w[932] = 4'h1;
    assign d2_w[933] = 4'h1;
    assign d2_w[934] = 4'h2;
    assign d2_w[935] = 4'hE;
    assign d2_w[936] = 4'hF;
    assign d2_w[937] = 4'hE;
    assign d2_w[938] = 4'hF;
    assign d2_w[939] = 4'hF;
    assign d2_w[940] = 4'h1;
    assign d2_w[941] = 4'hE;
    assign d2_w[942] = 4'h2;
    assign d2_w[943] = 4'hF;
    assign d2_w[944] = 4'hE;
    assign d2_w[945] = 4'hF;
    assign d2_w[946] = 4'hF;
    assign d2_w[947] = 4'h2;
    assign d2_w[948] = 4'hE;
    assign d2_w[949] = 4'h0;
    assign d2_w[950] = 4'h2;
    assign d2_w[951] = 4'h0;
    assign d2_w[952] = 4'hE;
    assign d2_w[953] = 4'hE;
    assign d2_w[954] = 4'hE;
    assign d2_w[955] = 4'h2;
    assign d2_w[956] = 4'hF;
    assign d2_w[957] = 4'hF;
    assign d2_w[958] = 4'hE;
    assign d2_w[959] = 4'h1;
    assign d2_w[960] = 4'h2;
    assign d2_w[961] = 4'h0;
    assign d2_w[962] = 4'hE;
    assign d2_w[963] = 4'hF;
    assign d2_w[964] = 4'h1;
    assign d2_w[965] = 4'h1;
    assign d2_w[966] = 4'h0;
    assign d2_w[967] = 4'h1;
    assign d2_w[968] = 4'h0;
    assign d2_w[969] = 4'hF;
    assign d2_w[970] = 4'h1;
    assign d2_w[971] = 4'hE;
    assign d2_w[972] = 4'h1;
    assign d2_w[973] = 4'h2;
    assign d2_w[974] = 4'h2;
    assign d2_w[975] = 4'h0;
    assign d2_w[976] = 4'h1;
    assign d2_w[977] = 4'hF;
    assign d2_w[978] = 4'h2;
    assign d2_w[979] = 4'hE;
    assign d2_w[980] = 4'hE;
    assign d2_w[981] = 4'hF;
    assign d2_w[982] = 4'h1;
    assign d2_w[983] = 4'hE;
    assign d2_w[984] = 4'hF;
    assign d2_w[985] = 4'h2;
    assign d2_w[986] = 4'h0;
    assign d2_w[987] = 4'hE;
    assign d2_w[988] = 4'hE;
    assign d2_w[989] = 4'hF;
    assign d2_w[990] = 4'hF;
    assign d2_w[991] = 4'h0;
    assign d2_w[992] = 4'h1;
    assign d2_w[993] = 4'h0;
    assign d2_w[994] = 4'hF;
    assign d2_w[995] = 4'hE;
    assign d2_w[996] = 4'hE;
    assign d2_w[997] = 4'h1;
    assign d2_w[998] = 4'hF;
    assign d2_w[999] = 4'hF;
    assign d2_w[1000] = 4'hF;
    assign d2_w[1001] = 4'hE;
    assign d2_w[1002] = 4'hF;
    assign d2_w[1003] = 4'hE;
    assign d2_w[1004] = 4'h2;
    assign d2_w[1005] = 4'hE;
    assign d2_w[1006] = 4'h1;
    assign d2_w[1007] = 4'hF;
    assign d2_w[1008] = 4'h1;
    assign d2_w[1009] = 4'hE;
    assign d2_w[1010] = 4'hE;
    assign d2_w[1011] = 4'hE;
    assign d2_w[1012] = 4'h0;
    assign d2_w[1013] = 4'hF;
    assign d2_w[1014] = 4'h0;
    assign d2_w[1015] = 4'h1;
    assign d2_w[1016] = 4'h2;
    assign d2_w[1017] = 4'h2;
    assign d2_w[1018] = 4'h2;
    assign d2_w[1019] = 4'hF;
    assign d2_w[1020] = 4'hE;
    assign d2_w[1021] = 4'hF;
    assign d2_w[1022] = 4'hE;
    assign d2_w[1023] = 4'h1;

    // --- layer2_b ---
    assign d2_b[0] = 4'h5;
    assign d2_b[1] = 4'h6;
    assign d2_b[2] = 4'h7;
    assign d2_b[3] = 4'h6;
    assign d2_b[4] = 4'h6;
    assign d2_b[5] = 4'hB;
    assign d2_b[6] = 4'h6;
    assign d2_b[7] = 4'h7;
    assign d2_b[8] = 4'h6;
    assign d2_b[9] = 4'h6;
    assign d2_b[10] = 4'h0;
    assign d2_b[11] = 4'h6;
    assign d2_b[12] = 4'hB;
    assign d2_b[13] = 4'h6;
    assign d2_b[14] = 4'h6;
    assign d2_b[15] = 4'h6;
    assign d2_b[16] = 4'h0;
    assign d2_b[17] = 4'hC;
    assign d2_b[18] = 4'h2;
    assign d2_b[19] = 4'hB;
    assign d2_b[20] = 4'h6;
    assign d2_b[21] = 4'h0;
    assign d2_b[22] = 4'h6;
    assign d2_b[23] = 4'h0;
    assign d2_b[24] = 4'hB;
    assign d2_b[25] = 4'h0;
    assign d2_b[26] = 4'h0;
    assign d2_b[27] = 4'hA;
    assign d2_b[28] = 4'h0;
    assign d2_b[29] = 4'h6;
    assign d2_b[30] = 4'h6;
    assign d2_b[31] = 4'h0;

    // --- layer3_w ---
    assign d3_w[0] = 4'h4;
    assign d3_w[1] = 4'h2;
    assign d3_w[2] = 4'h4;
    assign d3_w[3] = 4'h2;
    assign d3_w[4] = 4'h1;
    assign d3_w[5] = 4'hE;
    assign d3_w[6] = 4'h3;
    assign d3_w[7] = 4'h3;
    assign d3_w[8] = 4'h1;
    assign d3_w[9] = 4'h3;
    assign d3_w[10] = 4'hF;
    assign d3_w[11] = 4'h5;
    assign d3_w[12] = 4'hE;
    assign d3_w[13] = 4'h7;
    assign d3_w[14] = 4'h2;
    assign d3_w[15] = 4'h6;
    assign d3_w[16] = 4'hD;
    assign d3_w[17] = 4'hD;
    assign d3_w[18] = 4'h3;
    assign d3_w[19] = 4'hF;
    assign d3_w[20] = 4'h4;
    assign d3_w[21] = 4'hF;
    assign d3_w[22] = 4'h7;
    assign d3_w[23] = 4'hF;
    assign d3_w[24] = 4'hD;
    assign d3_w[25] = 4'hE;
    assign d3_w[26] = 4'h0;
    assign d3_w[27] = 4'hF;
    assign d3_w[28] = 4'hE;
    assign d3_w[29] = 4'h4;
    assign d3_w[30] = 4'h5;
    assign d3_w[31] = 4'hD;

    // --- layer3_b ---
    assign d3_b = 4'h7;


endmodule 